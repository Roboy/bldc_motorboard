// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Aug 25 2019 21:32:08

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    output PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    input PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22317;
    wire N__22316;
    wire N__22315;
    wire N__22308;
    wire N__22307;
    wire N__22306;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22271;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22246;
    wire N__22243;
    wire N__22238;
    wire N__22235;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22213;
    wire N__22210;
    wire N__22205;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22173;
    wire N__22170;
    wire N__22163;
    wire N__22162;
    wire N__22161;
    wire N__22160;
    wire N__22159;
    wire N__22158;
    wire N__22157;
    wire N__22156;
    wire N__22155;
    wire N__22154;
    wire N__22153;
    wire N__22152;
    wire N__22151;
    wire N__22150;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22111;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22096;
    wire N__22093;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22018;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21926;
    wire N__21925;
    wire N__21924;
    wire N__21923;
    wire N__21922;
    wire N__21921;
    wire N__21920;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21916;
    wire N__21915;
    wire N__21914;
    wire N__21913;
    wire N__21912;
    wire N__21911;
    wire N__21910;
    wire N__21909;
    wire N__21908;
    wire N__21907;
    wire N__21906;
    wire N__21905;
    wire N__21904;
    wire N__21903;
    wire N__21902;
    wire N__21901;
    wire N__21900;
    wire N__21899;
    wire N__21898;
    wire N__21897;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21890;
    wire N__21889;
    wire N__21888;
    wire N__21887;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21883;
    wire N__21882;
    wire N__21881;
    wire N__21880;
    wire N__21879;
    wire N__21878;
    wire N__21877;
    wire N__21876;
    wire N__21875;
    wire N__21874;
    wire N__21873;
    wire N__21872;
    wire N__21871;
    wire N__21870;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21866;
    wire N__21865;
    wire N__21864;
    wire N__21863;
    wire N__21862;
    wire N__21861;
    wire N__21860;
    wire N__21859;
    wire N__21858;
    wire N__21857;
    wire N__21856;
    wire N__21855;
    wire N__21854;
    wire N__21853;
    wire N__21852;
    wire N__21851;
    wire N__21850;
    wire N__21849;
    wire N__21848;
    wire N__21847;
    wire N__21846;
    wire N__21845;
    wire N__21844;
    wire N__21843;
    wire N__21842;
    wire N__21841;
    wire N__21840;
    wire N__21839;
    wire N__21838;
    wire N__21837;
    wire N__21836;
    wire N__21835;
    wire N__21834;
    wire N__21833;
    wire N__21832;
    wire N__21831;
    wire N__21830;
    wire N__21829;
    wire N__21828;
    wire N__21827;
    wire N__21826;
    wire N__21825;
    wire N__21824;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21596;
    wire N__21595;
    wire N__21594;
    wire N__21593;
    wire N__21592;
    wire N__21591;
    wire N__21590;
    wire N__21589;
    wire N__21588;
    wire N__21587;
    wire N__21586;
    wire N__21585;
    wire N__21584;
    wire N__21583;
    wire N__21582;
    wire N__21581;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21512;
    wire N__21509;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21497;
    wire N__21496;
    wire N__21495;
    wire N__21494;
    wire N__21491;
    wire N__21486;
    wire N__21485;
    wire N__21482;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21461;
    wire N__21456;
    wire N__21453;
    wire N__21452;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21425;
    wire N__21422;
    wire N__21413;
    wire N__21412;
    wire N__21411;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21396;
    wire N__21395;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21349;
    wire N__21344;
    wire N__21339;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21299;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21282;
    wire N__21279;
    wire N__21278;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21266;
    wire N__21261;
    wire N__21256;
    wire N__21245;
    wire N__21244;
    wire N__21243;
    wire N__21242;
    wire N__21241;
    wire N__21232;
    wire N__21229;
    wire N__21228;
    wire N__21227;
    wire N__21224;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21194;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21179;
    wire N__21174;
    wire N__21171;
    wire N__21164;
    wire N__21159;
    wire N__21156;
    wire N__21149;
    wire N__21146;
    wire N__21145;
    wire N__21144;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21133;
    wire N__21132;
    wire N__21123;
    wire N__21122;
    wire N__21119;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21097;
    wire N__21096;
    wire N__21093;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21071;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21059;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21041;
    wire N__21040;
    wire N__21039;
    wire N__21034;
    wire N__21033;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21011;
    wire N__21010;
    wire N__21009;
    wire N__21006;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20984;
    wire N__20983;
    wire N__20980;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20922;
    wire N__20921;
    wire N__20920;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20908;
    wire N__20903;
    wire N__20902;
    wire N__20901;
    wire N__20896;
    wire N__20891;
    wire N__20884;
    wire N__20879;
    wire N__20878;
    wire N__20875;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20861;
    wire N__20860;
    wire N__20859;
    wire N__20858;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20846;
    wire N__20845;
    wire N__20844;
    wire N__20843;
    wire N__20840;
    wire N__20833;
    wire N__20832;
    wire N__20831;
    wire N__20826;
    wire N__20821;
    wire N__20818;
    wire N__20813;
    wire N__20810;
    wire N__20803;
    wire N__20800;
    wire N__20795;
    wire N__20790;
    wire N__20787;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20749;
    wire N__20746;
    wire N__20745;
    wire N__20742;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20734;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20715;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20666;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20584;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20534;
    wire N__20533;
    wire N__20532;
    wire N__20529;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20515;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20486;
    wire N__20483;
    wire N__20474;
    wire N__20471;
    wire N__20470;
    wire N__20469;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20457;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20443;
    wire N__20442;
    wire N__20439;
    wire N__20434;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20404;
    wire N__20399;
    wire N__20392;
    wire N__20391;
    wire N__20390;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20375;
    wire N__20372;
    wire N__20365;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20355;
    wire N__20354;
    wire N__20349;
    wire N__20346;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20340;
    wire N__20339;
    wire N__20338;
    wire N__20335;
    wire N__20334;
    wire N__20333;
    wire N__20332;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20321;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20290;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20279;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20275;
    wire N__20274;
    wire N__20271;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20255;
    wire N__20252;
    wire N__20245;
    wire N__20242;
    wire N__20237;
    wire N__20234;
    wire N__20229;
    wire N__20216;
    wire N__20211;
    wire N__20204;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20161;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20145;
    wire N__20142;
    wire N__20137;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20090;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20079;
    wire N__20078;
    wire N__20069;
    wire N__20066;
    wire N__20061;
    wire N__20054;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20046;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19967;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19935;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19850;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19804;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19793;
    wire N__19792;
    wire N__19789;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19759;
    wire N__19758;
    wire N__19755;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19739;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19727;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19713;
    wire N__19712;
    wire N__19707;
    wire N__19702;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19648;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19630;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19607;
    wire N__19606;
    wire N__19605;
    wire N__19604;
    wire N__19601;
    wire N__19600;
    wire N__19599;
    wire N__19596;
    wire N__19591;
    wire N__19588;
    wire N__19583;
    wire N__19574;
    wire N__19573;
    wire N__19572;
    wire N__19569;
    wire N__19568;
    wire N__19565;
    wire N__19564;
    wire N__19563;
    wire N__19560;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19542;
    wire N__19541;
    wire N__19540;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19523;
    wire N__19520;
    wire N__19515;
    wire N__19510;
    wire N__19503;
    wire N__19502;
    wire N__19497;
    wire N__19494;
    wire N__19493;
    wire N__19492;
    wire N__19489;
    wire N__19488;
    wire N__19487;
    wire N__19486;
    wire N__19485;
    wire N__19484;
    wire N__19483;
    wire N__19482;
    wire N__19481;
    wire N__19480;
    wire N__19475;
    wire N__19466;
    wire N__19459;
    wire N__19454;
    wire N__19449;
    wire N__19446;
    wire N__19441;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19412;
    wire N__19411;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19403;
    wire N__19402;
    wire N__19401;
    wire N__19400;
    wire N__19399;
    wire N__19398;
    wire N__19397;
    wire N__19396;
    wire N__19393;
    wire N__19388;
    wire N__19381;
    wire N__19376;
    wire N__19375;
    wire N__19374;
    wire N__19373;
    wire N__19372;
    wire N__19371;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19363;
    wire N__19362;
    wire N__19361;
    wire N__19358;
    wire N__19351;
    wire N__19348;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19323;
    wire N__19322;
    wire N__19321;
    wire N__19320;
    wire N__19319;
    wire N__19318;
    wire N__19315;
    wire N__19314;
    wire N__19313;
    wire N__19312;
    wire N__19311;
    wire N__19302;
    wire N__19293;
    wire N__19288;
    wire N__19287;
    wire N__19286;
    wire N__19283;
    wire N__19278;
    wire N__19275;
    wire N__19266;
    wire N__19263;
    wire N__19258;
    wire N__19253;
    wire N__19238;
    wire N__19237;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19222;
    wire N__19219;
    wire N__19218;
    wire N__19215;
    wire N__19214;
    wire N__19213;
    wire N__19210;
    wire N__19209;
    wire N__19206;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19197;
    wire N__19186;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19174;
    wire N__19173;
    wire N__19172;
    wire N__19171;
    wire N__19170;
    wire N__19169;
    wire N__19168;
    wire N__19163;
    wire N__19162;
    wire N__19159;
    wire N__19158;
    wire N__19153;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19129;
    wire N__19120;
    wire N__19115;
    wire N__19114;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19096;
    wire N__19081;
    wire N__19078;
    wire N__19077;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19061;
    wire N__19058;
    wire N__19051;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18971;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18957;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18932;
    wire N__18929;
    wire N__18928;
    wire N__18927;
    wire N__18926;
    wire N__18925;
    wire N__18924;
    wire N__18923;
    wire N__18922;
    wire N__18921;
    wire N__18912;
    wire N__18911;
    wire N__18910;
    wire N__18907;
    wire N__18898;
    wire N__18897;
    wire N__18896;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18881;
    wire N__18874;
    wire N__18873;
    wire N__18868;
    wire N__18861;
    wire N__18858;
    wire N__18853;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18802;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18782;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18746;
    wire N__18743;
    wire N__18742;
    wire N__18739;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18724;
    wire N__18719;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18650;
    wire N__18649;
    wire N__18648;
    wire N__18645;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18627;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18604;
    wire N__18599;
    wire N__18590;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18572;
    wire N__18569;
    wire N__18564;
    wire N__18561;
    wire N__18554;
    wire N__18551;
    wire N__18550;
    wire N__18549;
    wire N__18546;
    wire N__18541;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18500;
    wire N__18497;
    wire N__18496;
    wire N__18495;
    wire N__18494;
    wire N__18493;
    wire N__18492;
    wire N__18487;
    wire N__18486;
    wire N__18483;
    wire N__18482;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18464;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18430;
    wire N__18429;
    wire N__18424;
    wire N__18423;
    wire N__18420;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18412;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18371;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18357;
    wire N__18352;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18323;
    wire N__18322;
    wire N__18321;
    wire N__18318;
    wire N__18313;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18301;
    wire N__18298;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18281;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18273;
    wire N__18272;
    wire N__18269;
    wire N__18262;
    wire N__18257;
    wire N__18254;
    wire N__18253;
    wire N__18252;
    wire N__18249;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18241;
    wire N__18238;
    wire N__18235;
    wire N__18230;
    wire N__18227;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18211;
    wire N__18210;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18178;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18155;
    wire N__18154;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18122;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18080;
    wire N__18073;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18040;
    wire N__18037;
    wire N__18036;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18021;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17999;
    wire N__17996;
    wire N__17995;
    wire N__17992;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17960;
    wire N__17957;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17945;
    wire N__17942;
    wire N__17941;
    wire N__17938;
    wire N__17937;
    wire N__17934;
    wire N__17931;
    wire N__17926;
    wire N__17921;
    wire N__17918;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17906;
    wire N__17905;
    wire N__17904;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17900;
    wire N__17897;
    wire N__17890;
    wire N__17883;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17869;
    wire N__17866;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17858;
    wire N__17857;
    wire N__17856;
    wire N__17851;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17839;
    wire N__17836;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17821;
    wire N__17816;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17795;
    wire N__17790;
    wire N__17787;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17726;
    wire N__17725;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17712;
    wire N__17705;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17693;
    wire N__17692;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17609;
    wire N__17606;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17563;
    wire N__17562;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17554;
    wire N__17553;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17541;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17521;
    wire N__17520;
    wire N__17517;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17505;
    wire N__17504;
    wire N__17503;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17476;
    wire N__17475;
    wire N__17470;
    wire N__17467;
    wire N__17462;
    wire N__17455;
    wire N__17452;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17434;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17419;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17379;
    wire N__17378;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17362;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17345;
    wire N__17344;
    wire N__17343;
    wire N__17342;
    wire N__17341;
    wire N__17340;
    wire N__17339;
    wire N__17338;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17300;
    wire N__17299;
    wire N__17298;
    wire N__17297;
    wire N__17296;
    wire N__17295;
    wire N__17294;
    wire N__17293;
    wire N__17292;
    wire N__17291;
    wire N__17290;
    wire N__17289;
    wire N__17288;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17188;
    wire N__17185;
    wire N__17184;
    wire N__17181;
    wire N__17180;
    wire N__17179;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17171;
    wire N__17168;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17147;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17128;
    wire N__17127;
    wire N__17126;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17111;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17055;
    wire N__17050;
    wire N__17047;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17024;
    wire N__17023;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17004;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16883;
    wire N__16882;
    wire N__16881;
    wire N__16878;
    wire N__16877;
    wire N__16876;
    wire N__16875;
    wire N__16872;
    wire N__16871;
    wire N__16870;
    wire N__16869;
    wire N__16868;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16856;
    wire N__16851;
    wire N__16844;
    wire N__16843;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16809;
    wire N__16808;
    wire N__16807;
    wire N__16800;
    wire N__16795;
    wire N__16788;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16768;
    wire N__16763;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16741;
    wire N__16738;
    wire N__16737;
    wire N__16734;
    wire N__16731;
    wire N__16726;
    wire N__16721;
    wire N__16718;
    wire N__16717;
    wire N__16716;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16708;
    wire N__16703;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16641;
    wire N__16638;
    wire N__16635;
    wire N__16628;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16620;
    wire N__16619;
    wire N__16616;
    wire N__16615;
    wire N__16612;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16588;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16541;
    wire N__16538;
    wire N__16533;
    wire N__16530;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16516;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16462;
    wire N__16461;
    wire N__16458;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16446;
    wire N__16439;
    wire N__16438;
    wire N__16437;
    wire N__16436;
    wire N__16435;
    wire N__16434;
    wire N__16433;
    wire N__16432;
    wire N__16429;
    wire N__16424;
    wire N__16423;
    wire N__16422;
    wire N__16421;
    wire N__16420;
    wire N__16415;
    wire N__16408;
    wire N__16403;
    wire N__16400;
    wire N__16393;
    wire N__16382;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16370;
    wire N__16367;
    wire N__16366;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16352;
    wire N__16351;
    wire N__16350;
    wire N__16349;
    wire N__16348;
    wire N__16347;
    wire N__16346;
    wire N__16341;
    wire N__16338;
    wire N__16331;
    wire N__16326;
    wire N__16321;
    wire N__16318;
    wire N__16307;
    wire N__16306;
    wire N__16305;
    wire N__16304;
    wire N__16303;
    wire N__16302;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16231;
    wire N__16228;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16201;
    wire N__16198;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16186;
    wire N__16181;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16167;
    wire N__16166;
    wire N__16161;
    wire N__16156;
    wire N__16151;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16125;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16103;
    wire N__16100;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16067;
    wire N__16064;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16050;
    wire N__16049;
    wire N__16044;
    wire N__16039;
    wire N__16034;
    wire N__16031;
    wire N__16030;
    wire N__16029;
    wire N__16026;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16007;
    wire N__16004;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15960;
    wire N__15955;
    wire N__15952;
    wire N__15947;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15922;
    wire N__15917;
    wire N__15914;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15902;
    wire N__15899;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15891;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15811;
    wire N__15810;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15791;
    wire N__15782;
    wire N__15781;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15761;
    wire N__15760;
    wire N__15757;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15737;
    wire N__15734;
    wire N__15733;
    wire N__15732;
    wire N__15729;
    wire N__15724;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15698;
    wire N__15695;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15670;
    wire N__15669;
    wire N__15666;
    wire N__15661;
    wire N__15660;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15618;
    wire N__15613;
    wire N__15610;
    wire N__15605;
    wire N__15602;
    wire N__15601;
    wire N__15598;
    wire N__15597;
    wire N__15596;
    wire N__15595;
    wire N__15594;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15526;
    wire N__15525;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15461;
    wire N__15460;
    wire N__15457;
    wire N__15456;
    wire N__15453;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15424;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15407;
    wire N__15406;
    wire N__15403;
    wire N__15402;
    wire N__15401;
    wire N__15398;
    wire N__15391;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15383;
    wire N__15380;
    wire N__15375;
    wire N__15372;
    wire N__15365;
    wire N__15362;
    wire N__15361;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15350;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15332;
    wire N__15331;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15308;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15287;
    wire N__15286;
    wire N__15283;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15265;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15247;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15239;
    wire N__15236;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15217;
    wire N__15214;
    wire N__15209;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15159;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15143;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15135;
    wire N__15130;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15110;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15062;
    wire N__15061;
    wire N__15060;
    wire N__15057;
    wire N__15056;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15023;
    wire N__15022;
    wire N__15021;
    wire N__15018;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14978;
    wire N__14975;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14960;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14940;
    wire N__14939;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14921;
    wire N__14920;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14875;
    wire N__14872;
    wire N__14861;
    wire N__14860;
    wire N__14857;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14843;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14803;
    wire N__14800;
    wire N__14799;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14787;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14719;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14642;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14630;
    wire N__14629;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14618;
    wire N__14615;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14603;
    wire N__14600;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14558;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14550;
    wire N__14547;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14529;
    wire N__14526;
    wire N__14519;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14511;
    wire N__14506;
    wire N__14505;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14474;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14435;
    wire N__14434;
    wire N__14433;
    wire N__14432;
    wire N__14431;
    wire N__14430;
    wire N__14429;
    wire N__14422;
    wire N__14421;
    wire N__14420;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14409;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14391;
    wire N__14384;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14354;
    wire N__14351;
    wire N__14350;
    wire N__14349;
    wire N__14348;
    wire N__14347;
    wire N__14344;
    wire N__14343;
    wire N__14342;
    wire N__14341;
    wire N__14340;
    wire N__14337;
    wire N__14330;
    wire N__14327;
    wire N__14322;
    wire N__14317;
    wire N__14314;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14293;
    wire N__14292;
    wire N__14291;
    wire N__14288;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14233;
    wire N__14232;
    wire N__14229;
    wire N__14226;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14214;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14200;
    wire N__14199;
    wire N__14196;
    wire N__14191;
    wire N__14186;
    wire N__14185;
    wire N__14184;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14151;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14139;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14086;
    wire N__14083;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14066;
    wire N__14065;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14023;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14009;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13982;
    wire N__13979;
    wire N__13970;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13962;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13950;
    wire N__13943;
    wire N__13940;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13928;
    wire N__13927;
    wire N__13924;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13891;
    wire N__13888;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13878;
    wire N__13871;
    wire N__13868;
    wire N__13867;
    wire N__13864;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13847;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13823;
    wire N__13820;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13808;
    wire N__13805;
    wire N__13804;
    wire N__13803;
    wire N__13800;
    wire N__13795;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13783;
    wire N__13782;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13770;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13739;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13731;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13709;
    wire N__13706;
    wire N__13705;
    wire N__13702;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13690;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13660;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13643;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13635;
    wire N__13630;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13613;
    wire N__13610;
    wire N__13609;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13585;
    wire N__13582;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13521;
    wire N__13514;
    wire N__13511;
    wire N__13510;
    wire N__13507;
    wire N__13504;
    wire N__13501;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13418;
    wire N__13415;
    wire N__13410;
    wire N__13405;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13393;
    wire N__13392;
    wire N__13391;
    wire N__13390;
    wire N__13389;
    wire N__13388;
    wire N__13387;
    wire N__13386;
    wire N__13383;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13363;
    wire N__13362;
    wire N__13361;
    wire N__13360;
    wire N__13359;
    wire N__13358;
    wire N__13357;
    wire N__13356;
    wire N__13355;
    wire N__13354;
    wire N__13353;
    wire N__13352;
    wire N__13351;
    wire N__13350;
    wire N__13349;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13331;
    wire N__13330;
    wire N__13327;
    wire N__13320;
    wire N__13315;
    wire N__13304;
    wire N__13303;
    wire N__13302;
    wire N__13301;
    wire N__13300;
    wire N__13299;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13261;
    wire N__13260;
    wire N__13255;
    wire N__13252;
    wire N__13251;
    wire N__13250;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13236;
    wire N__13231;
    wire N__13228;
    wire N__13219;
    wire N__13214;
    wire N__13207;
    wire N__13190;
    wire N__13187;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13163;
    wire N__13160;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13148;
    wire N__13147;
    wire N__13144;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13093;
    wire N__13092;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13060;
    wire N__13059;
    wire N__13056;
    wire N__13051;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13030;
    wire N__13029;
    wire N__13026;
    wire N__13021;
    wire N__13016;
    wire N__13013;
    wire N__13012;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__13000;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12981;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12934;
    wire N__12933;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12896;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12821;
    wire N__12820;
    wire N__12817;
    wire N__12814;
    wire N__12811;
    wire N__12806;
    wire N__12803;
    wire N__12794;
    wire N__12791;
    wire N__12790;
    wire N__12787;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12770;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12587;
    wire N__12584;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12496;
    wire N__12493;
    wire N__12492;
    wire N__12491;
    wire N__12488;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12474;
    wire N__12467;
    wire N__12464;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12362;
    wire N__12361;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12340;
    wire N__12337;
    wire N__12332;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12233;
    wire N__12232;
    wire N__12231;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12148;
    wire N__12145;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12133;
    wire N__12130;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12118;
    wire N__12115;
    wire N__12110;
    wire N__12107;
    wire N__12106;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12098;
    wire N__12097;
    wire N__12094;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12043;
    wire N__12038;
    wire N__12035;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11995;
    wire N__11992;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11960;
    wire N__11957;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11919;
    wire N__11912;
    wire N__11911;
    wire N__11908;
    wire N__11907;
    wire N__11904;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11883;
    wire N__11880;
    wire N__11873;
    wire N__11870;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11837;
    wire N__11834;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11743;
    wire N__11740;
    wire N__11739;
    wire N__11736;
    wire N__11731;
    wire N__11728;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11709;
    wire N__11704;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11653;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11605;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11588;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11498;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11420;
    wire N__11419;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11396;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11372;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11321;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11270;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11249;
    wire N__11246;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11222;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11210;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11150;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11138;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11126;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11114;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11077;
    wire N__11076;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11064;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10787;
    wire N__10784;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10595;
    wire N__10592;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10471;
    wire N__10470;
    wire N__10469;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10454;
    wire N__10453;
    wire N__10450;
    wire N__10445;
    wire N__10442;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10431;
    wire N__10428;
    wire N__10423;
    wire N__10420;
    wire N__10409;
    wire N__10408;
    wire N__10407;
    wire N__10404;
    wire N__10403;
    wire N__10402;
    wire N__10399;
    wire N__10398;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10378;
    wire N__10375;
    wire N__10370;
    wire N__10369;
    wire N__10368;
    wire N__10363;
    wire N__10358;
    wire N__10355;
    wire N__10350;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10328;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10304;
    wire N__10303;
    wire N__10302;
    wire N__10301;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10289;
    wire N__10282;
    wire N__10273;
    wire N__10262;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10256;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10245;
    wire N__10244;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10213;
    wire N__10210;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10190;
    wire N__10187;
    wire N__10182;
    wire N__10175;
    wire N__10172;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10045;
    wire N__10044;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10022;
    wire N__10021;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10017;
    wire N__10012;
    wire N__10007;
    wire N__10002;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9985;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9969;
    wire N__9966;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9924;
    wire N__9919;
    wire N__9916;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9872;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9853;
    wire N__9850;
    wire N__9847;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9800;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9778;
    wire N__9777;
    wire N__9774;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9766;
    wire N__9763;
    wire N__9756;
    wire N__9753;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9653;
    wire N__9650;
    wire N__9649;
    wire N__9644;
    wire N__9641;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9598;
    wire N__9593;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9361;
    wire N__9360;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9348;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9327;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9319;
    wire N__9316;
    wire N__9315;
    wire N__9314;
    wire N__9313;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9297;
    wire N__9292;
    wire N__9289;
    wire N__9278;
    wire N__9277;
    wire N__9276;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9265;
    wire N__9264;
    wire N__9263;
    wire N__9262;
    wire N__9259;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9248;
    wire N__9247;
    wire N__9244;
    wire N__9243;
    wire N__9242;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9225;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9204;
    wire N__9201;
    wire N__9200;
    wire N__9197;
    wire N__9196;
    wire N__9195;
    wire N__9192;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9180;
    wire N__9175;
    wire N__9166;
    wire N__9161;
    wire N__9156;
    wire N__9153;
    wire N__9144;
    wire N__9135;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9109;
    wire N__9108;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9089;
    wire N__9088;
    wire N__9085;
    wire N__9084;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9072;
    wire N__9071;
    wire N__9070;
    wire N__9065;
    wire N__9062;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9031;
    wire N__9022;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8996;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8992;
    wire N__8991;
    wire N__8990;
    wire N__8989;
    wire N__8988;
    wire N__8987;
    wire N__8986;
    wire N__8985;
    wire N__8982;
    wire N__8977;
    wire N__8974;
    wire N__8969;
    wire N__8966;
    wire N__8957;
    wire N__8948;
    wire N__8933;
    wire N__8932;
    wire N__8931;
    wire N__8930;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8905;
    wire N__8902;
    wire N__8901;
    wire N__8900;
    wire N__8899;
    wire N__8896;
    wire N__8895;
    wire N__8894;
    wire N__8893;
    wire N__8890;
    wire N__8883;
    wire N__8880;
    wire N__8879;
    wire N__8878;
    wire N__8877;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8860;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8834;
    wire N__8833;
    wire N__8832;
    wire N__8831;
    wire N__8828;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8813;
    wire N__8808;
    wire N__8807;
    wire N__8806;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8789;
    wire N__8784;
    wire N__8781;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8740;
    wire N__8737;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8720;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8687;
    wire N__8684;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8623;
    wire N__8622;
    wire N__8621;
    wire N__8620;
    wire N__8617;
    wire N__8616;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8612;
    wire N__8611;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8561;
    wire N__8560;
    wire N__8559;
    wire N__8556;
    wire N__8555;
    wire N__8554;
    wire N__8553;
    wire N__8550;
    wire N__8549;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8528;
    wire N__8527;
    wire N__8524;
    wire N__8513;
    wire N__8508;
    wire N__8501;
    wire N__8500;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8419;
    wire N__8418;
    wire N__8415;
    wire N__8410;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8359;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire CLK_ibuf_gb_io_gb_input;
    wire VCCG0;
    wire PIN_2_c;
    wire \c0.rx.r_Rx_Data_RZ0 ;
    wire \c0.rx.rx_data_ready ;
    wire \c0.rx.un1_r_Clock_Count_5_c2_cascade_ ;
    wire \c0.rx.g0_i_o4_0_1_cascade_ ;
    wire \c0.rx.g0_i_o2_2_3_cascade_ ;
    wire \c0.rx.g0_i_a4_1_1 ;
    wire PIN_1_c;
    wire \c0.rx.un1_r_Rx_DV7_0 ;
    wire \c0.rx.g0_i_o2_5 ;
    wire \c0.rx.g0_i_o2_4 ;
    wire \c0.rx.g0_i_o2_6 ;
    wire \c0.rx.g0_i_a4_1_3 ;
    wire \c0.rx.N_7_cascade_ ;
    wire \c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1 ;
    wire \c0.rx.N_10_0 ;
    wire \c0.rx.N_13_0 ;
    wire \c0.rx.N_12_1_cascade_ ;
    wire \c0.rx.un1_r_Clock_Count_5_c2 ;
    wire \c0.rx.N_6_cascade_ ;
    wire \c0.rx.r_Clock_Count_2_sqmuxa_0 ;
    wire \c0.rx.r_Clock_Count_2_sqmuxa_0_cascade_ ;
    wire \c0.rx.g1_4 ;
    wire \c0.rx.g1_5_cascade_ ;
    wire \c0.rx.g1 ;
    wire \c0.rx.g0_0_1_cascade_ ;
    wire \c0.rx.r_Clock_Count14_cascade_ ;
    wire \c0.rx.m6_ns_1 ;
    wire \c0.rx.un1_r_Clock_Count_5_m_0_cascade_ ;
    wire \c0.rx.un1_r_Clock_Count_2_sqmuxa_0 ;
    wire \c0.rx.r_Clock_Count_1_sqmuxa_0 ;
    wire \c0.rx.un1_r_Clock_Count_5_m_1_cascade_ ;
    wire N_12;
    wire N_8_0;
    wire LED_c;
    wire \c0.rx.CO1_cascade_ ;
    wire \c0.rx.g0_i_o3_0_4_cascade_ ;
    wire \c0.rx.N_10 ;
    wire \c0.rx.N_12_0 ;
    wire \c0.rx.N_9_0_cascade_ ;
    wire \c0.rx.N_11_i ;
    wire \c0.rx.r_Clock_CountZ0Z_6 ;
    wire \c0.rx.r_Clock_CountZ0Z_5 ;
    wire \c0.rx.r_Clock_CountZ0Z_7 ;
    wire \c0.rx.r_Clock_CountZ0Z_4 ;
    wire \c0.rx.r_Clock_Count14_3_cascade_ ;
    wire \c0.rx.r_Clock_Count26_cascade_ ;
    wire \c0.rx.r_Clock_CountZ0Z_2 ;
    wire \c0.rx.r_Clock_CountZ0Z_3 ;
    wire \c0.rx.g0_i_a4_0_3_cascade_ ;
    wire \c0.rx.r_Clock_Count14_3 ;
    wire \c0.rx.N_13 ;
    wire \c0.rx.r_Clock_Count26 ;
    wire \c0.rx.r_SM_MainZ0Z_2 ;
    wire \c0.rx.r_Rx_DV_1_sqmuxa_cascade_ ;
    wire \c0.rx.r_SM_MainZ0Z_1 ;
    wire \c0.rx.r_SM_MainZ0Z_0 ;
    wire \c0.rx.r_Clock_Count14 ;
    wire \c0.rx.N_9 ;
    wire \c0.rx.r_Clock_CountZ0Z_0 ;
    wire \c0.rx.r_Clock_CountZ0Z_1 ;
    wire \c0.rx.r_Clock_Count14_1 ;
    wire bfn_5_25_0_;
    wire \c0.tx.un1_r_Clock_Count_cry_0 ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_2 ;
    wire \c0.tx.un1_r_Clock_Count_cry_1 ;
    wire \c0.tx.un1_r_Clock_Count_cry_2 ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_3_cascade_ ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_0 ;
    wire \c0.tx.r_Clock_CountZ0Z_0 ;
    wire \c0.tx.r_Clock_Count_0_sqmuxa ;
    wire \c0.tx.r_Clock_Count_RNO_0Z0Z_1 ;
    wire blink_counterZ0Z_0;
    wire bfn_6_20_0_;
    wire blink_counterZ0Z_1;
    wire blink_counter_cry_0;
    wire blink_counterZ0Z_2;
    wire blink_counter_cry_1;
    wire blink_counterZ0Z_3;
    wire blink_counter_cry_2;
    wire blink_counterZ0Z_4;
    wire blink_counter_cry_3;
    wire blink_counterZ0Z_5;
    wire blink_counter_cry_4;
    wire blink_counterZ0Z_6;
    wire blink_counter_cry_5;
    wire blink_counterZ0Z_7;
    wire blink_counter_cry_6;
    wire blink_counter_cry_7;
    wire blink_counterZ0Z_8;
    wire bfn_6_21_0_;
    wire blink_counterZ0Z_9;
    wire blink_counter_cry_8;
    wire blink_counterZ0Z_10;
    wire blink_counter_cry_9;
    wire blink_counterZ0Z_11;
    wire blink_counter_cry_10;
    wire blink_counterZ0Z_12;
    wire blink_counter_cry_11;
    wire blink_counterZ0Z_13;
    wire blink_counter_cry_12;
    wire blink_counterZ0Z_14;
    wire blink_counter_cry_13;
    wire blink_counterZ0Z_15;
    wire blink_counter_cry_14;
    wire blink_counter_cry_15;
    wire blink_counterZ0Z_16;
    wire bfn_6_22_0_;
    wire blink_counterZ0Z_17;
    wire blink_counter_cry_16;
    wire blink_counterZ0Z_18;
    wire blink_counter_cry_17;
    wire blink_counterZ0Z_19;
    wire blink_counter_cry_18;
    wire blink_counterZ0Z_20;
    wire blink_counter_cry_19;
    wire blink_counterZ0Z_21;
    wire blink_counter_cry_20;
    wire blink_counterZ0Z_22;
    wire blink_counter_cry_21;
    wire blink_counterZ0Z_23;
    wire blink_counter_cry_22;
    wire blink_counter_cry_23;
    wire blink_counterZ0Z_24;
    wire bfn_6_23_0_;
    wire blink_counter_cry_24;
    wire blink_counterZ0Z_25;
    wire \c0.tx.N_287_cascade_ ;
    wire \c0.tx.N_294 ;
    wire \c0.tx.o_Tx_Serial12 ;
    wire \c0.tx.N_294_cascade_ ;
    wire \c0.tx.m5_0_0 ;
    wire \c0.tx.N_287 ;
    wire \c0.tx.N_288_cascade_ ;
    wire \c0.tx.r_Clock_Count_i_0 ;
    wire bfn_6_25_0_;
    wire \c0.tx.r_Clock_CountZ0Z_1 ;
    wire \c0.tx.r_Clock_Count_i_1 ;
    wire \c0.tx.r_Clock_Count12_cry_0 ;
    wire \c0.tx.r_Clock_CountZ0Z_2 ;
    wire \c0.tx.r_Clock_Count_i_2 ;
    wire \c0.tx.r_Clock_Count12_cry_1 ;
    wire \c0.tx.r_Clock_CountZ0Z_3 ;
    wire \c0.tx.r_Clock_Count_i_3 ;
    wire \c0.tx.r_Clock_Count12_cry_2 ;
    wire \c0.tx.r_Clock_Count12 ;
    wire \c0.rx.r_Rx_Bytece_1_1_cascade_ ;
    wire \c0.rx.r_Rx_Bytece_1_5 ;
    wire \c0.rx.r_Rx_DV6 ;
    wire \c0.tx.r_Tx_Active_1_sqmuxa_cascade_ ;
    wire \c0.tx_data_RNO_0Z0Z_1 ;
    wire \c0.tx.r_Tx_DataZ0Z_1 ;
    wire \c0.tx.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_3_cascade_ ;
    wire \c0.tx.r_Tx_DataZ0Z_3 ;
    wire \c0.tx_data_RNO_1Z0Z_5 ;
    wire \c0.tx.r_Tx_DataZ0Z_5 ;
    wire \c0.tx_data_RNO_4Z0Z_3 ;
    wire \c0.tx.r_Bit_IndexZ0Z_2 ;
    wire \c0.tx.r_Bit_IndexZ0Z_1 ;
    wire \c0.tx.r_Tx_Data_pmux_3_i_m2_ns_1_cascade_ ;
    wire \c0.tx.N_354 ;
    wire \c0.tx.r_Bit_IndexZ0Z_0 ;
    wire \c0.tx.N_357_cascade_ ;
    wire \c0.tx.N_320 ;
    wire \c0.tx_data_RNO_3Z0Z_5_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_5 ;
    wire \c0.tx_data_RNO_1Z0Z_0_cascade_ ;
    wire \c0.tx.r_Tx_DataZ0Z_0 ;
    wire \c0.tx.r_Tx_DataZ0Z_4 ;
    wire \c0.data_out_7_Z0Z_5 ;
    wire \c0.rx.r_Rx_Bytece_0_3_cascade_ ;
    wire \c0.rx_data_3 ;
    wire \c0.tx2_data_RNO_3Z0Z_2_cascade_ ;
    wire \c0.tx.r_SM_MainZ0Z_0 ;
    wire \c0.tx.r_SM_MainZ0Z_1 ;
    wire \c0.tx.r_Clock_Count12_THRU_CO ;
    wire \c0.tx.r_SM_MainZ0Z_2 ;
    wire \c0.nextCRC16_3_3_12_cascade_ ;
    wire \c0.nextCRC16_3_4_12 ;
    wire \c0.data_out_6_Z0Z_4 ;
    wire \c0.tx_data_RNO_0Z0Z_4 ;
    wire \c0.tx_data_RNO_4Z0Z_1_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_1 ;
    wire \c0.tx_data_RNO_0Z0Z_3 ;
    wire \c0.nextCRC16_3_0_a2_1_11_cascade_ ;
    wire \c0.data_out_6_Z0Z_3 ;
    wire \c0.d_2_7 ;
    wire \c0.tx_data_RNO_3Z0Z_7_cascade_ ;
    wire \c0.tx_data_RNO_4Z0Z_7 ;
    wire \c0.N_74 ;
    wire \c0.N_74_cascade_ ;
    wire \c0.d_2_19 ;
    wire bfn_9_27_0_;
    wire \c0.dataZ0Z_1 ;
    wire \c0.data_cry_0 ;
    wire \c0.data_cry_1 ;
    wire \c0.data_cry_2 ;
    wire \c0.data_cry_3 ;
    wire \c0.data_cry_4 ;
    wire \c0.data_cry_5 ;
    wire \c0.data_cry_6 ;
    wire \c0.data_cry_7 ;
    wire bfn_9_28_0_;
    wire \c0.data_cry_8 ;
    wire \c0.data_cry_9 ;
    wire \c0.dataZ0Z_11 ;
    wire \c0.data_cry_10 ;
    wire \c0.dataZ0Z_12 ;
    wire \c0.data_cry_11 ;
    wire \c0.data_cry_12 ;
    wire \c0.dataZ0Z_14 ;
    wire \c0.data_cry_13 ;
    wire \c0.data_cry_14 ;
    wire \c0.i12_0_and ;
    wire bfn_10_17_0_;
    wire \c0.i12_0 ;
    wire \c0.i12_2_and ;
    wire \c0.i12_1 ;
    wire \c0.i12_2 ;
    wire \c0.i12_3 ;
    wire \c0.i12_5_and ;
    wire \c0.i12_4 ;
    wire \c0.i12_5 ;
    wire \c0.i12_6 ;
    wire \c0.i12 ;
    wire bfn_10_18_0_;
    wire \c0.i12_1_and ;
    wire \c0.i12_3_and ;
    wire \c0.i12_4_and ;
    wire \c0.i12_6_and ;
    wire \c0.rx_data_5 ;
    wire \c0.tx2_data_RNO_4Z0Z_2 ;
    wire \c0.tx2_data_RNO_1Z0Z_2 ;
    wire \c0.tx2_data_RNO_0Z0Z_2_cascade_ ;
    wire \c0.tx2_data_1_0_i_ns_1_2 ;
    wire \c0.tx2_data_1_iv_4_3 ;
    wire \c0.rx.un1_r_Rx_Byte_7 ;
    wire \c0.tx2.o_Tx_Serial12_cascade_ ;
    wire \c0.tx_data_RNO_3Z0Z_3 ;
    wire \c0.d_2_38 ;
    wire \c0.m115_amcf1 ;
    wire \c0.N_293_cascade_ ;
    wire \c0.tx_data_1_0_i_1_6 ;
    wire \c0.tx_data_RNO_1Z0Z_6_cascade_ ;
    wire \c0.tx.r_Tx_DataZ0Z_6 ;
    wire \c0.tx.r_Tx_DataZ0Z_2 ;
    wire \c0.tx_data_1_0_i_ns_1_7 ;
    wire \c0.tx.r_Tx_DataZ0Z_7 ;
    wire \c0.tx.r_Tx_Data_0_sqmuxa ;
    wire \c0.tx_data_RNO_1Z0Z_4 ;
    wire \c0.data_out_6_Z0Z_1 ;
    wire \c0.tx_data_RNO_0Z0Z_5 ;
    wire \c0.d_2_23 ;
    wire \c0.tx_data_RNO_0Z0Z_7 ;
    wire \c0.tx_data_RNO_1Z0Z_1 ;
    wire \c0.tx_data_RNO_1Z0Z_2 ;
    wire \c0.nextCRC16_3_0_a2_1_15_cascade_ ;
    wire \c0.tx_data_RNO_3Z0Z_4_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_4 ;
    wire \c0.tx_data_RNO_4Z0Z_4 ;
    wire \c0.data_out_7_Z0Z_4 ;
    wire \c0.dataZ0Z_7 ;
    wire \c0.dataZ0Z_3 ;
    wire \c0.dataZ0Z_10 ;
    wire \c0.dataZ0Z_6 ;
    wire \c0.dataZ0Z_2 ;
    wire \c0.data_out_7_Z0Z_2 ;
    wire \c0.dataZ0Z_5 ;
    wire \c0.dataZ0Z_13 ;
    wire \c0.d_2_37 ;
    wire \c0.dataZ0Z_4 ;
    wire \c0.dataZ0Z_9 ;
    wire \c0.i12_7_and ;
    wire \c0.g1_1_cascade_ ;
    wire \c0.N_72_mux ;
    wire \c0.N_249_cascade_ ;
    wire \c0.data_in_4_Z0Z_0 ;
    wire \c0.g1_cascade_ ;
    wire \c0.g0_3 ;
    wire \c0.byte_transmit_counter2_0_sqmuxa_0 ;
    wire \c0.g3_2_0_cascade_ ;
    wire \c0.g0_2 ;
    wire \c0.rx_data_1 ;
    wire \c0.data_in_3_Z0Z_4 ;
    wire \c0.data_in_1_Z0Z_6 ;
    wire \c0.data_in_3_Z0Z_5 ;
    wire \c0.data_in_5_Z0Z_2 ;
    wire bfn_11_22_0_;
    wire \c0.tx2.un1_r_Clock_Count_cry_0 ;
    wire \c0.tx2.r_Clock_Count_RNO_0_0_2 ;
    wire \c0.tx2.un1_r_Clock_Count_cry_1 ;
    wire \c0.tx2.un1_r_Clock_Count_cry_2 ;
    wire \c0.tx2.r_Clock_Count_RNO_0_0_3 ;
    wire \c0.tx2.r_Clock_Count_0_sqmuxa ;
    wire \c0.tx2.r_Clock_Count_RNO_0_0_0 ;
    wire \c0.tx2.r_Clock_CountZ0Z_0 ;
    wire \c0.tx2.r_Clock_Count_RNO_0_0_1 ;
    wire \c0.tx2.r_Clock_Count_i_0 ;
    wire bfn_11_23_0_;
    wire \c0.tx2.r_Clock_CountZ0Z_1 ;
    wire \c0.tx2.r_Clock_Count_i_1 ;
    wire \c0.tx2.r_Clock_Count12_cry_0 ;
    wire \c0.tx2.r_Clock_CountZ0Z_2 ;
    wire \c0.tx2.r_Clock_Count_i_2 ;
    wire \c0.tx2.r_Clock_Count12_cry_1 ;
    wire \c0.tx2.r_Clock_CountZ0Z_3 ;
    wire \c0.tx2.r_Clock_Count_i_3 ;
    wire \c0.tx2.r_Clock_Count12_cry_2 ;
    wire \c0.tx2.r_Clock_Count12 ;
    wire \c0.N_76 ;
    wire \c0.data_out_6_Z0Z_2 ;
    wire \c0.tx_data_RNO_0Z0Z_2 ;
    wire \c0.d_2_21 ;
    wire \c0.tx_data_1_iv_i_m2_0_ns_1_0_cascade_ ;
    wire \c0.N_304_cascade_ ;
    wire \c0.tx_data_1_iv_i_1_0 ;
    wire \c0.nextCRC16_3_0_a2_1_8 ;
    wire \c0.N_77 ;
    wire \c0.data_out_6_Z0Z_0 ;
    wire \c0.dataZ0Z_0 ;
    wire \c0.data_out_7_Z0Z_0 ;
    wire \c0.d_2_8 ;
    wire \c0.tx_data_RNO_0Z0Z_0 ;
    wire \c0.N_93 ;
    wire \c0.nextCRC16_3_0_a2_0_10 ;
    wire \c0.d_2_22 ;
    wire \c0.d_2_6 ;
    wire \c0.nextCRC16_3_9 ;
    wire \c0.nextCRC16_3_0_a2_6_0_15_cascade_ ;
    wire \c0.N_92 ;
    wire \c0.d_2_41 ;
    wire \c0.d_2_12 ;
    wire \c0.d_2_40 ;
    wire \c0.nextCRC16_3_0_a2_2_2 ;
    wire \c0.d_2_3 ;
    wire \c0.N_75 ;
    wire \c0.N_75_cascade_ ;
    wire \c0.d_2_44 ;
    wire \c0.N_95 ;
    wire \c0.d_2_14 ;
    wire \c0.N_95_cascade_ ;
    wire \c0.d_2_25 ;
    wire \c0.d_2_11 ;
    wire \c0.dataZ0Z_8 ;
    wire \c0.dataZ0Z_15 ;
    wire \c0.tx2_active ;
    wire \c0.tx2_data_1_iv_5_1_0_7 ;
    wire \c0.tx2_data_1_iv_5_1_7_cascade_ ;
    wire \c0.data_in_frame_6_Z0Z_7 ;
    wire \c0.tx2_data_1_iv_3_1_3 ;
    wire \c0.tx2_data_1_iv_3_3 ;
    wire \c0.data_in_0_Z0Z_3 ;
    wire \c0.N_247_0 ;
    wire \c0.un1_data_in_6__0_0_a2_5_a2_2_cascade_ ;
    wire \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_ ;
    wire \c0.un1_data_in_7__4_i_cascade_ ;
    wire \c0.un1_data_in_6__0 ;
    wire \c0.d_4_RNIF73E2Z0Z_14_cascade_ ;
    wire \c0.d_4_RNIMKFE3Z0Z_14_cascade_ ;
    wire \c0.un1_data_in_6__7_cascade_ ;
    wire \c0.wait_for_transmission4_12 ;
    wire \c0.data_in_frame_0__0_sqmuxa ;
    wire \c0.wait_for_transmission4_12_cascade_ ;
    wire \c0.un1_data_in_7__4_0_a2_0_a2_4 ;
    wire \c0.data_in_0_Z0Z_2 ;
    wire \c0.d_4_RNID6K21_0Z0Z_15 ;
    wire \c0.d_4_RNID6K21Z0Z_15 ;
    wire \c0.data_in_0_Z0Z_1 ;
    wire \c0.data_in_1_Z0Z_7 ;
    wire \c0.data_in_3_Z0Z_7 ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_2_cascade_ ;
    wire \c0.d_4_2 ;
    wire \c0.N_103 ;
    wire \c0.wait_for_transmission4_13_1_1 ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_6_cascade_ ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_1_cascade_ ;
    wire \c0.un1_data_in_7__1_0_a2_24_a2_5 ;
    wire \c0.d_4_RNITCRCZ0Z_29 ;
    wire \c0.tx2_data_RNO_4Z0Z_0_cascade_ ;
    wire \c0.tx2_data_RNO_0Z0Z_0 ;
    wire \c0.tx2_data_1_0_i_ns_1_0_cascade_ ;
    wire \c0.d_4_1 ;
    wire \c0.tx2_data_RNO_3Z0Z_1_cascade_ ;
    wire \c0.tx2_data_RNO_1Z0Z_1 ;
    wire \c0.tx2_data_1_0_i_ns_1_1_cascade_ ;
    wire \c0.tx2_data_RNO_0Z0Z_1 ;
    wire \c0.tx2_data_RNO_4Z0Z_1 ;
    wire \c0.tx2_data_RNO_1Z0Z_0 ;
    wire \c0.tx2.r_Tx_DataZ0Z_2 ;
    wire \c0.tx2.r_Tx_DataZ0Z_0 ;
    wire \c0.tx2.r_Tx_Data_pmux_3_i_m2_ns_1 ;
    wire \c0.tx2.r_Tx_DataZ0Z_1 ;
    wire \c0.tx2.r_Tx_DataZ0Z_3 ;
    wire \c0.tx2.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_ ;
    wire \c0.tx2.N_349 ;
    wire \c0.tx2.N_346_cascade_ ;
    wire \c0.tx2.N_279_cascade_ ;
    wire PIN_3_c;
    wire \c0.tx2.r_Tx_Active_1_sqmuxa ;
    wire \c0.tx_data_RNO_3Z0Z_1 ;
    wire \c0.tx2.m5_0_0_cascade_ ;
    wire \c0.d_2_9 ;
    wire \c0.N_94 ;
    wire \c0.tx_data_RNO_4Z0Z_5 ;
    wire \c0.d_2_45 ;
    wire \c0.nextCRC16_3_0_a2_0_0 ;
    wire \c0.nextCRC16_3_0_a2_4_0 ;
    wire \c0.d_2_28 ;
    wire \c0.nextCRC16_3_0_a2_1_2 ;
    wire \c0.d_2_0 ;
    wire \c0.nextCRC16_3_4_0 ;
    wire \c0.d_2_13 ;
    wire \c0.d_2_26 ;
    wire \c0.nextCRC16_3_4_0_cascade_ ;
    wire \c0.N_99 ;
    wire \c0.nextCRC16_3_0_a2_3_0 ;
    wire \c0.d_2_39 ;
    wire \c0.data_out_6_Z0Z_5 ;
    wire \c0.nextCRC16_3_0_a2_4_15 ;
    wire \c0.nextCRC16_3_0_a2_3_15 ;
    wire \c0.data_out_6_Z0Z_7 ;
    wire \c0.d_2_16 ;
    wire \c0.d_2_24 ;
    wire CONSTANT_ONE_NET;
    wire \c0.N_105 ;
    wire \c0.nextCRC16_3_2_1 ;
    wire \c0.N_106 ;
    wire \c0.data_out_7_Z0Z_1 ;
    wire \c0.data_in_frame_7_Z0Z_5 ;
    wire \c0.data_in_frame_7_Z0Z_7 ;
    wire \c0.wait_for_transmission_RNOZ0Z_10_cascade_ ;
    wire \c0.g0_5_4 ;
    wire \c0.d_4_3 ;
    wire \c0.d_4_45 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_2 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_3_cascade_ ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_5 ;
    wire \c0.g3_2_1 ;
    wire \c0.g0_3_0 ;
    wire \c0.un1_data_in_7__0_0_a2_1_a2_3_cascade_ ;
    wire \c0.un1_data_in_7__0_0_a2_1_a2_5_0_cascade_ ;
    wire \c0.tx2_transmit_0_sqmuxa_1 ;
    wire \c0.un1_data_in_7__3_0_a2_0_a2_3_cascade_ ;
    wire \c0.N_129 ;
    wire \c0.data_in_2_Z0Z_1 ;
    wire \c0.d_4_17 ;
    wire \c0.data_in_3_Z0Z_6 ;
    wire \c0.data_in_0_Z0Z_0 ;
    wire \c0.data_in_2_Z0Z_0 ;
    wire \c0.d_4_16 ;
    wire \c0.d_4_0 ;
    wire \c0.tx2_data_RNO_3Z0Z_0 ;
    wire \c0.data_in_0_Z0Z_4 ;
    wire \c0.data_in_4_Z0Z_2 ;
    wire \c0.data_in_1_Z0Z_3 ;
    wire \c0.data_in_1_Z0Z_5 ;
    wire \c0.data_in_2_Z0Z_5 ;
    wire \c0.data_in_3_Z0Z_1 ;
    wire \c0.data_in_5_Z0Z_1 ;
    wire \c0.data_in_3_Z0Z_3 ;
    wire \c0.tx2_data_1_iv_3_1_6_cascade_ ;
    wire \c0.d_4_34 ;
    wire \c0.un1_data_in_7__7_i ;
    wire \c0.tx2_data_1_0_i_1_3 ;
    wire \c0.tx2_data_1_iv_4_1_0_3 ;
    wire \c0.data_in_1_Z0Z_4 ;
    wire \c0.data_in_7_Z0Z_3 ;
    wire \c0.data_in_frame_7_Z0Z_3 ;
    wire \c0.d_4_14 ;
    wire \c0.d_4_30 ;
    wire \c0.tx2_data_1_iv_4_1_6_cascade_ ;
    wire \c0.data_in_5_Z0Z_3 ;
    wire \c0.tx2.r_SM_MainZ0Z_2 ;
    wire \c0.tx2.r_SM_MainZ0Z_0 ;
    wire \c0.tx2.N_257_cascade_ ;
    wire \c0.tx2.N_261 ;
    wire \c0.tx2.o_Tx_Serial12 ;
    wire \c0.tx2.N_261_cascade_ ;
    wire \c0.tx2.r_Bit_IndexZ0Z_2 ;
    wire \c0.tx_transmitZ0 ;
    wire \c0.tx_active ;
    wire \c0.tx2_data_1_iv_4_6 ;
    wire \c0.tx2_data_1_iv_3_6 ;
    wire \c0.tx2.r_Tx_DataZ0Z_6 ;
    wire \c0.d_2_27 ;
    wire \c0.tx_data_RNO_1Z0Z_3 ;
    wire \c0.data_out_7_Z0Z_7 ;
    wire \c0.tx_data_RNO_1Z0Z_7 ;
    wire \c0.tx_data_RNO_3Z0Z_2_cascade_ ;
    wire \c0.tx_data_1_0_i_ns_1_2 ;
    wire \c0.d_2_10 ;
    wire \c0.d_2_42 ;
    wire \c0.tx_data_RNO_4Z0Z_2 ;
    wire \c0.N_81 ;
    wire \c0.d_2_29 ;
    wire \c0.d_2_30 ;
    wire \c0.data_out_7_Z0Z_3 ;
    wire \c0.d_2_31 ;
    wire \c0.d_2_43 ;
    wire \c0.d_2_15 ;
    wire \c0.d_2_2 ;
    wire \c0.d_2_47 ;
    wire \c0.un105_newcrc_0_a2_3_cascade_ ;
    wire \c0.un105_newcrc_0_a2_4 ;
    wire \c0.d_2_5 ;
    wire \c0.d_2_32 ;
    wire \c0.d_2_18 ;
    wire \c0.d_2_46 ;
    wire \c0.d_2_20 ;
    wire \c0.nextCRC16_3_3_1 ;
    wire \c0.d_2_17 ;
    wire \c0.d_2_1 ;
    wire \c0.d_2_4 ;
    wire \c0.nextCRC16_3_0_a2_1_1 ;
    wire \c0.un1_data_in_6__4_0_a2_5_a2_1 ;
    wire \c0.N_133 ;
    wire \c0.un1_data_in_7__2_0_a2_0_a2_5 ;
    wire \c0.un1_data_in_6__4 ;
    wire \c0.wait_for_transmission4_12_5_1_cascade_ ;
    wire \c0.N_108 ;
    wire \c0.d_4_32 ;
    wire \c0.un1_data_in_7__6_0_a2_5_a2_2 ;
    wire \c0.wait_for_transmission_RNOZ0Z_11 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_4_1 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_4_1_cascade_ ;
    wire \c0.d_4_47 ;
    wire \c0.N_125 ;
    wire \c0.data_in_0_Z0Z_6 ;
    wire \c0.d_4_6 ;
    wire \c0.data_in_2_Z0Z_3 ;
    wire \c0.d_4_19 ;
    wire \c0.un1_data_in_6__7_0_a2_17_a2_4_1_0 ;
    wire \c0.data_in_4_Z0Z_3 ;
    wire \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_ ;
    wire \c0.g3_2 ;
    wire \c0.un1_data_in_6__6_0_a2_0_a2_3_cascade_ ;
    wire \c0.N_128 ;
    wire \c0.d_4_41 ;
    wire \c0.un1_data_in_6__5_0_a2_5_a2_2_cascade_ ;
    wire \c0.N_132 ;
    wire \c0.un1_data_in_6__6_0_a2_0_a2_3 ;
    wire \c0.un1_data_in_6__5_cascade_ ;
    wire \c0.g0_2_0 ;
    wire \c0.d_4_43 ;
    wire \c0.un1_data_in_7__0_0_a2_1_a2_2 ;
    wire \c0.un1_data_in_6__3_0_a2_5_a2_2_cascade_ ;
    wire \c0.d_4_25 ;
    wire \c0.un1_data_in_6__3 ;
    wire \c0.un1_data_in_6__3_0_a2_5_a2_1 ;
    wire \c0.data_in_1_Z0Z_1 ;
    wire \c0.data_in_2_Z0Z_7 ;
    wire \c0.data_in_5_Z0Z_0 ;
    wire \c0.d_4_40 ;
    wire \c0.un1_data_in_7__7_0_a2_0_a2_2 ;
    wire \c0.data_in_0_Z0Z_5 ;
    wire \c0.wait_for_transmission_RNOZ0Z_9 ;
    wire \c0.data_in_2_Z0Z_2 ;
    wire \c0.data_in_2_Z0Z_4 ;
    wire \c0.d_4_18 ;
    wire \c0.N_124 ;
    wire \c0.N_124_cascade_ ;
    wire \c0.d_4_RNI21N6Z0Z_11 ;
    wire \c0.d_4_RNIPF9J2Z0Z_37 ;
    wire \c0.data_in_4_Z0Z_1 ;
    wire \c0.d_4_33 ;
    wire \c0.data_in_frame_6_Z0Z_0 ;
    wire \c0.data_in_3_Z0Z_2 ;
    wire \c0.d_4_26 ;
    wire \c0.data_in_frame_6_Z0Z_1 ;
    wire \c0.data_in_1_Z0Z_2 ;
    wire \c0.d_4_10 ;
    wire \c0.data_in_frame_7_Z0Z_0 ;
    wire \c0.d_2_36 ;
    wire \c0.d_2_35 ;
    wire \c0.N_71 ;
    wire \c0.tx2.r_Bit_IndexZ0Z_0 ;
    wire \c0.tx2.r_Clock_Count12_THRU_CO ;
    wire \c0.tx2.N_257 ;
    wire \c0.tx2.N_258_cascade_ ;
    wire \c0.tx2.r_SM_MainZ0Z_1 ;
    wire \c0.tx2.r_Bit_IndexZ0Z_1 ;
    wire \c0.data_out_6_Z0Z_6 ;
    wire \c0.N_4_0_cascade_ ;
    wire \c0.N_197 ;
    wire \c0.data_out_0__1_sqmuxa ;
    wire \c0.byte_transmit_counterZ0Z_6 ;
    wire \c0.byte_transmit_counterZ0Z_3 ;
    wire \c0.m2_e_1_cascade_ ;
    wire \c0.N_129_mux_cascade_ ;
    wire \c0.N_86 ;
    wire \c0.byte_transmit_counterZ0Z_1 ;
    wire \c0.byte_transmit_counterZ0Z_4 ;
    wire \c0.byte_transmit_counterZ0Z_0 ;
    wire \c0.un144_newcrc_3 ;
    wire \c0.d_2_34 ;
    wire \c0.un144_newcrc_4 ;
    wire \c0.d_2_33 ;
    wire \c0.data_out_7_Z0Z_6 ;
    wire \c0.data_out_0__1_sqmuxa_g ;
    wire \c0.d_4_12 ;
    wire \c0.d_4_44 ;
    wire \c0.tx2_data_1_iv_5_7 ;
    wire \c0.tx2_data_1_0_i_1_7 ;
    wire \c0.tx2.r_Tx_DataZ0Z_7 ;
    wire \c0.d_4_13 ;
    wire \c0.d_4_29 ;
    wire \c0.data_in_frame_1__m_5_cascade_ ;
    wire \c0.tx2_data_1_0_i_1_5 ;
    wire \c0.tx2_data_1_iv_1_5_cascade_ ;
    wire \c0.tx2.r_Tx_DataZ0Z_5 ;
    wire \c0.d_4_15 ;
    wire \c0.data_in_frame_1__m_7_cascade_ ;
    wire \c0.d_4_31 ;
    wire \c0.tx2_data_1_iv_1_7 ;
    wire \c0.N_205 ;
    wire \c0.d_4_27 ;
    wire \c0.N_205_cascade_ ;
    wire \c0.d_4_11 ;
    wire \c0.tx2_data_1_iv_4_1_3 ;
    wire \c0.un1_data_in_6__5 ;
    wire \c0.i12_THRU_CO ;
    wire \c0.N_136 ;
    wire \c0.wait_for_transmission4_13_1 ;
    wire \c0.g1_3_cascade_ ;
    wire \c0.un1_data_in_7__0_0_a2_1_a2_5_0 ;
    wire \c0.i12_7_c_RNIP740G_cascade_ ;
    wire \c0.g1_2 ;
    wire \c0.wait_for_transmission4_12_5 ;
    wire \c0.un1_data_in_7__3_i ;
    wire \c0.g1_5_cascade_ ;
    wire \c0.wait_for_transmission4_12_4 ;
    wire \c0.d_4_RNI9LFUVZ0Z_43_cascade_ ;
    wire \c0.wait_for_transmission_RNI9PP5BZ0Z1_cascade_ ;
    wire \c0.un1_data_in_6__1_1 ;
    wire \c0.g0_2_3 ;
    wire \c0.d_4_23 ;
    wire \c0.N_126_cascade_ ;
    wire \c0.un1_data_in_6__1 ;
    wire \c0.d_4_35 ;
    wire \c0.data_in_0_Z0Z_7 ;
    wire \c0.d_4_7 ;
    wire \c0.data_in_1_Z0Z_0 ;
    wire \c0.d_4_8 ;
    wire \c0.d_4_9 ;
    wire \c0.d_4_39 ;
    wire \c0.un1_data_in_6__2_0 ;
    wire \c0.N_107 ;
    wire \c0.un1_data_in_6__2_0_a2_6_a2_2 ;
    wire \c0.N_107_cascade_ ;
    wire \c0.un1_data_in_6__2 ;
    wire \c0.data_in_2_Z0Z_6 ;
    wire \c0.d_4_22 ;
    wire \c0.d_4_RNIU6U8Z0Z_22 ;
    wire \c0.d_4_RNIU6U8_0Z0Z_22_cascade_ ;
    wire \c0.d_4_RNIMI4KZ0Z_37 ;
    wire \c0.data_in_3_Z0Z_0 ;
    wire \c0.d_4_24 ;
    wire \c0.N_126 ;
    wire \c0.un1_data_in_6__1_0_a2_4_a2_1 ;
    wire \c0.un1_data_in_6__1_0 ;
    wire \c0.data_in_4_Z0Z_4 ;
    wire \c0.d_4_36 ;
    wire \c0.data_in_frame_6_Z0Z_4 ;
    wire \c0.tx2_data_1_iv_4_1_0_6 ;
    wire \c0.data_in_frame_7_Z0Z_6 ;
    wire \c0.d_4_42 ;
    wire \c0.d_4_46 ;
    wire \c0.un1_data_in_7__2_0_a2_0_a2_4 ;
    wire \c0.data_in_4_Z0Z_7 ;
    wire \c0.rx_data_7 ;
    wire \c0.data_in_6_Z0Z_1 ;
    wire \c0.data_in_6_Z0Z_0 ;
    wire \c0.data_in_7_Z0Z_0 ;
    wire \c0.data_in_5_Z0Z_4 ;
    wire \c0.byte_transmit_counterZ0Z_5 ;
    wire \c0.N_201 ;
    wire \c0.N_129_mux ;
    wire \c0.byte_transmit_counterZ0Z_2 ;
    wire GNDG0;
    wire \c0.byte_transmit_counterZ0Z_7 ;
    wire \c0.byte_transmit_counter15 ;
    wire \c0.tx2_data_1_iv_5_1_0_4 ;
    wire \c0.N_207 ;
    wire \c0.N_207_cascade_ ;
    wire \c0.d_4_28 ;
    wire \c0.m2_e_0_2_cascade_ ;
    wire \c0.N_71_mux ;
    wire \c0.d_4_RNII9QU3Z0Z_14 ;
    wire \c0.wait_for_transmission_RNI94LSZ0Z6 ;
    wire \c0.wait_for_transmissionZ0 ;
    wire \c0.d_4_RNI9LFUVZ0Z_43 ;
    wire \c0.tx2_transmitZ0 ;
    wire \c0.m2_e_0_2 ;
    wire \c0.d_4_20 ;
    wire \c0.N_203_cascade_ ;
    wire \c0.d_4_4 ;
    wire \c0.tx2_data_1_iv_5_1_4 ;
    wire \c0.un1_m4_0_a2_2_cascade_ ;
    wire \c0.byte_transmit_counter2Z0Z_7 ;
    wire \c0.un1_m4_0_a2_1_0 ;
    wire \c0.byte_transmit_counter2Z0Z_6 ;
    wire \c0.byte_transmit_counter2Z0Z_5 ;
    wire \c0.byte_transmit_counter2Z0Z_0 ;
    wire \c0.un1_byte_transmit_counter2_1_ac0_3_out_cascade_ ;
    wire \c0.wait_for_transmission_RNI9PP5BZ0Z1 ;
    wire \c0.tx2_transmit_0_sqmuxa ;
    wire \c0.data_in_4_Z0Z_5 ;
    wire \c0.data_in_5_Z0Z_5 ;
    wire \c0.data_in_7_Z0Z_5 ;
    wire \c0.data_in_6_Z0Z_5 ;
    wire \c0.data_in_5_Z0Z_6 ;
    wire \c0.data_in_7_Z0Z_6 ;
    wire \c0.data_in_6_Z0Z_3 ;
    wire \c0.data_in_frame_6_Z0Z_3 ;
    wire \c0.tx2_data_1_0_i_1_6 ;
    wire \c0.data_in_6_Z0Z_6 ;
    wire \c0.data_in_frame_6_Z0Z_6 ;
    wire \c0.data_in_4_Z0Z_6 ;
    wire \c0.d_4_38 ;
    wire \c0.d_4_5 ;
    wire \c0.d_4_21 ;
    wire \c0.N_203 ;
    wire \c0.tx2_data_1_iv_5_1_5_cascade_ ;
    wire \c0.byte_transmit_counter2Z0Z_2 ;
    wire \c0.tx2_data_1_iv_5_5 ;
    wire \c0.data_in_frame_6_Z0Z_5 ;
    wire \c0.d_4_37 ;
    wire \c0.tx2_data_1_iv_5_1_0_5 ;
    wire \c0.rx.r_Rx_Bytece_1_6 ;
    wire \c0.rx_data_6 ;
    wire \c0.rx.r_Rx_Bytece_1_2 ;
    wire \c0.rx_data_2 ;
    wire \c0.rx.r_Rx_Bytece_1_4_cascade_ ;
    wire \c0.rx_data_4 ;
    wire \c0.rx.r_Bit_IndexZ0Z_2 ;
    wire \c0.rx.r_Bit_IndexZ0Z_1 ;
    wire \c0.rx.r_Bit_IndexZ0Z_0 ;
    wire \c0.rx.r_Rx_DataZ0 ;
    wire \c0.rx.r_Rx_Bytece_1_0_cascade_ ;
    wire \c0.rx.r_Rx_Byte_1_sqmuxa ;
    wire \c0.rx_data_0 ;
    wire \c0.un1_byte_transmit_counter2_1_ac0_3_out ;
    wire \c0.byte_transmit_counter2Z0Z_3 ;
    wire \c0.byte_transmit_counter2Z0Z_4 ;
    wire \c0.un1_byte_transmit_counter2_1_ac0_7_out_0 ;
    wire \c0.tx2_data_1_iv_5_4 ;
    wire \c0.tx2_data_1_0_i_1_4 ;
    wire \c0.tx2_data_1_0_i_1_0_4 ;
    wire \c0.byte_transmit_counter2Z0Z_1 ;
    wire \c0.tx2.r_Tx_DataZ0Z_4 ;
    wire \c0.tx2.r_Tx_Data_0_sqmuxa ;
    wire \c0.data_in_5_Z0Z_7 ;
    wire \c0.data_in_6_Z0Z_4 ;
    wire \c0.data_in_7_Z0Z_7 ;
    wire \c0.data_in_6_Z0Z_7 ;
    wire \c0.rx_data_ready_g ;
    wire \c0.data_in_6_Z0Z_2 ;
    wire \c0.data_in_frame_6_Z0Z_2 ;
    wire \c0.data_in_7_Z0Z_1 ;
    wire \c0.data_in_frame_7_Z0Z_1 ;
    wire \c0.data_in_7_Z0Z_2 ;
    wire \c0.data_in_frame_7_Z0Z_2 ;
    wire \c0.data_in_7_Z0Z_4 ;
    wire \c0.data_in_frame_7_Z0Z_4 ;
    wire CLK_c_g;
    wire \c0.data_in_frame_0__0_sqmuxa_g ;
    wire _gnd_net_;

    IO_PAD LED_obuf_iopad (
            .OE(N__22335),
            .DIN(N__22334),
            .DOUT(N__22333),
            .PACKAGEPIN(LED));
    defparam LED_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_preio (
            .PADOEN(N__22335),
            .PADOUT(N__22334),
            .PADIN(N__22333),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8477),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PIN_1_obuf_iopad (
            .OE(N__22326),
            .DIN(N__22325),
            .DOUT(N__22324),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIN_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIN_1_obuf_preio (
            .PADOEN(N__22326),
            .PADOUT(N__22325),
            .PADIN(N__22324),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8336),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PIN_2_ibuf_iopad (
            .OE(N__22317),
            .DIN(N__22316),
            .DOUT(N__22315),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PIN_2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PIN_2_ibuf_preio (
            .PADOEN(N__22317),
            .PADOUT(N__22316),
            .PADIN(N__22315),
            .CLOCKENABLE(),
            .DIN0(PIN_2_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD PIN_3_obuf_iopad (
            .OE(N__22308),
            .DIN(N__22307),
            .DOUT(N__22306),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIN_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIN_3_obuf_preio (
            .PADOEN(N__22308),
            .PADOUT(N__22307),
            .PADIN(N__22306),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12668),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD USBPU_obuf_iopad (
            .OE(N__22299),
            .DIN(N__22298),
            .DOUT(N__22297),
            .PACKAGEPIN(USBPU));
    defparam USBPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam USBPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO USBPU_obuf_preio (
            .PADOEN(N__22299),
            .PADOUT(N__22298),
            .PADIN(N__22297),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__22290),
            .DIN(N__22289),
            .DOUT(N__22288),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__22290),
            .PADOUT(N__22289),
            .PADIN(N__22288),
            .CLOCKENABLE(),
            .DIN0(CLK_ibuf_gb_io_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__5372 (
            .O(N__22271),
            .I(N__22267));
    InMux I__5371 (
            .O(N__22270),
            .I(N__22264));
    InMux I__5370 (
            .O(N__22267),
            .I(N__22260));
    LocalMux I__5369 (
            .O(N__22264),
            .I(N__22257));
    InMux I__5368 (
            .O(N__22263),
            .I(N__22254));
    LocalMux I__5367 (
            .O(N__22260),
            .I(N__22251));
    Span4Mux_v I__5366 (
            .O(N__22257),
            .I(N__22246));
    LocalMux I__5365 (
            .O(N__22254),
            .I(N__22246));
    Span4Mux_h I__5364 (
            .O(N__22251),
            .I(N__22243));
    Odrv4 I__5363 (
            .O(N__22246),
            .I(\c0.data_in_6_Z0Z_4 ));
    Odrv4 I__5362 (
            .O(N__22243),
            .I(\c0.data_in_6_Z0Z_4 ));
    InMux I__5361 (
            .O(N__22238),
            .I(N__22235));
    LocalMux I__5360 (
            .O(N__22235),
            .I(N__22231));
    InMux I__5359 (
            .O(N__22234),
            .I(N__22228));
    Span4Mux_h I__5358 (
            .O(N__22231),
            .I(N__22224));
    LocalMux I__5357 (
            .O(N__22228),
            .I(N__22221));
    CascadeMux I__5356 (
            .O(N__22227),
            .I(N__22218));
    Span4Mux_v I__5355 (
            .O(N__22224),
            .I(N__22213));
    Span4Mux_h I__5354 (
            .O(N__22221),
            .I(N__22213));
    InMux I__5353 (
            .O(N__22218),
            .I(N__22210));
    Odrv4 I__5352 (
            .O(N__22213),
            .I(\c0.data_in_7_Z0Z_7 ));
    LocalMux I__5351 (
            .O(N__22210),
            .I(\c0.data_in_7_Z0Z_7 ));
    InMux I__5350 (
            .O(N__22205),
            .I(N__22202));
    LocalMux I__5349 (
            .O(N__22202),
            .I(N__22197));
    InMux I__5348 (
            .O(N__22201),
            .I(N__22194));
    InMux I__5347 (
            .O(N__22200),
            .I(N__22191));
    Span4Mux_h I__5346 (
            .O(N__22197),
            .I(N__22187));
    LocalMux I__5345 (
            .O(N__22194),
            .I(N__22184));
    LocalMux I__5344 (
            .O(N__22191),
            .I(N__22181));
    InMux I__5343 (
            .O(N__22190),
            .I(N__22178));
    Span4Mux_v I__5342 (
            .O(N__22187),
            .I(N__22173));
    Span4Mux_h I__5341 (
            .O(N__22184),
            .I(N__22173));
    Span4Mux_h I__5340 (
            .O(N__22181),
            .I(N__22170));
    LocalMux I__5339 (
            .O(N__22178),
            .I(\c0.data_in_6_Z0Z_7 ));
    Odrv4 I__5338 (
            .O(N__22173),
            .I(\c0.data_in_6_Z0Z_7 ));
    Odrv4 I__5337 (
            .O(N__22170),
            .I(\c0.data_in_6_Z0Z_7 ));
    CEMux I__5336 (
            .O(N__22163),
            .I(N__22121));
    CEMux I__5335 (
            .O(N__22162),
            .I(N__22121));
    CEMux I__5334 (
            .O(N__22161),
            .I(N__22121));
    CEMux I__5333 (
            .O(N__22160),
            .I(N__22121));
    CEMux I__5332 (
            .O(N__22159),
            .I(N__22121));
    CEMux I__5331 (
            .O(N__22158),
            .I(N__22121));
    CEMux I__5330 (
            .O(N__22157),
            .I(N__22121));
    CEMux I__5329 (
            .O(N__22156),
            .I(N__22121));
    CEMux I__5328 (
            .O(N__22155),
            .I(N__22121));
    CEMux I__5327 (
            .O(N__22154),
            .I(N__22121));
    CEMux I__5326 (
            .O(N__22153),
            .I(N__22121));
    CEMux I__5325 (
            .O(N__22152),
            .I(N__22121));
    CEMux I__5324 (
            .O(N__22151),
            .I(N__22121));
    CEMux I__5323 (
            .O(N__22150),
            .I(N__22121));
    GlobalMux I__5322 (
            .O(N__22121),
            .I(N__22118));
    gio2CtrlBuf I__5321 (
            .O(N__22118),
            .I(\c0.rx_data_ready_g ));
    InMux I__5320 (
            .O(N__22115),
            .I(N__22112));
    LocalMux I__5319 (
            .O(N__22112),
            .I(N__22107));
    InMux I__5318 (
            .O(N__22111),
            .I(N__22104));
    CascadeMux I__5317 (
            .O(N__22110),
            .I(N__22101));
    Span4Mux_h I__5316 (
            .O(N__22107),
            .I(N__22096));
    LocalMux I__5315 (
            .O(N__22104),
            .I(N__22096));
    InMux I__5314 (
            .O(N__22101),
            .I(N__22093));
    Odrv4 I__5313 (
            .O(N__22096),
            .I(\c0.data_in_6_Z0Z_2 ));
    LocalMux I__5312 (
            .O(N__22093),
            .I(\c0.data_in_6_Z0Z_2 ));
    InMux I__5311 (
            .O(N__22088),
            .I(N__22085));
    LocalMux I__5310 (
            .O(N__22085),
            .I(N__22082));
    Span4Mux_h I__5309 (
            .O(N__22082),
            .I(N__22079));
    Span4Mux_h I__5308 (
            .O(N__22079),
            .I(N__22076));
    Odrv4 I__5307 (
            .O(N__22076),
            .I(\c0.data_in_frame_6_Z0Z_2 ));
    InMux I__5306 (
            .O(N__22073),
            .I(N__22070));
    LocalMux I__5305 (
            .O(N__22070),
            .I(N__22066));
    InMux I__5304 (
            .O(N__22069),
            .I(N__22063));
    Span4Mux_v I__5303 (
            .O(N__22066),
            .I(N__22060));
    LocalMux I__5302 (
            .O(N__22063),
            .I(N__22057));
    Span4Mux_h I__5301 (
            .O(N__22060),
            .I(N__22053));
    Span4Mux_h I__5300 (
            .O(N__22057),
            .I(N__22050));
    InMux I__5299 (
            .O(N__22056),
            .I(N__22047));
    Odrv4 I__5298 (
            .O(N__22053),
            .I(\c0.data_in_7_Z0Z_1 ));
    Odrv4 I__5297 (
            .O(N__22050),
            .I(\c0.data_in_7_Z0Z_1 ));
    LocalMux I__5296 (
            .O(N__22047),
            .I(\c0.data_in_7_Z0Z_1 ));
    CascadeMux I__5295 (
            .O(N__22040),
            .I(N__22037));
    InMux I__5294 (
            .O(N__22037),
            .I(N__22034));
    LocalMux I__5293 (
            .O(N__22034),
            .I(N__22031));
    Span4Mux_h I__5292 (
            .O(N__22031),
            .I(N__22028));
    Span4Mux_h I__5291 (
            .O(N__22028),
            .I(N__22025));
    Odrv4 I__5290 (
            .O(N__22025),
            .I(\c0.data_in_frame_7_Z0Z_1 ));
    InMux I__5289 (
            .O(N__22022),
            .I(N__22019));
    LocalMux I__5288 (
            .O(N__22019),
            .I(N__22014));
    InMux I__5287 (
            .O(N__22018),
            .I(N__22011));
    InMux I__5286 (
            .O(N__22017),
            .I(N__22008));
    Span4Mux_v I__5285 (
            .O(N__22014),
            .I(N__22005));
    LocalMux I__5284 (
            .O(N__22011),
            .I(N__22002));
    LocalMux I__5283 (
            .O(N__22008),
            .I(N__21999));
    Odrv4 I__5282 (
            .O(N__22005),
            .I(\c0.data_in_7_Z0Z_2 ));
    Odrv4 I__5281 (
            .O(N__22002),
            .I(\c0.data_in_7_Z0Z_2 ));
    Odrv4 I__5280 (
            .O(N__21999),
            .I(\c0.data_in_7_Z0Z_2 ));
    InMux I__5279 (
            .O(N__21992),
            .I(N__21989));
    LocalMux I__5278 (
            .O(N__21989),
            .I(N__21986));
    Span12Mux_h I__5277 (
            .O(N__21986),
            .I(N__21983));
    Odrv12 I__5276 (
            .O(N__21983),
            .I(\c0.data_in_frame_7_Z0Z_2 ));
    CascadeMux I__5275 (
            .O(N__21980),
            .I(N__21977));
    InMux I__5274 (
            .O(N__21977),
            .I(N__21972));
    InMux I__5273 (
            .O(N__21976),
            .I(N__21969));
    InMux I__5272 (
            .O(N__21975),
            .I(N__21966));
    LocalMux I__5271 (
            .O(N__21972),
            .I(N__21963));
    LocalMux I__5270 (
            .O(N__21969),
            .I(N__21958));
    LocalMux I__5269 (
            .O(N__21966),
            .I(N__21958));
    Span4Mux_h I__5268 (
            .O(N__21963),
            .I(N__21955));
    Span4Mux_v I__5267 (
            .O(N__21958),
            .I(N__21952));
    Span4Mux_h I__5266 (
            .O(N__21955),
            .I(N__21949));
    Odrv4 I__5265 (
            .O(N__21952),
            .I(\c0.data_in_7_Z0Z_4 ));
    Odrv4 I__5264 (
            .O(N__21949),
            .I(\c0.data_in_7_Z0Z_4 ));
    InMux I__5263 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__5262 (
            .O(N__21941),
            .I(N__21938));
    Span4Mux_h I__5261 (
            .O(N__21938),
            .I(N__21935));
    Odrv4 I__5260 (
            .O(N__21935),
            .I(\c0.data_in_frame_7_Z0Z_4 ));
    ClkMux I__5259 (
            .O(N__21932),
            .I(N__21605));
    ClkMux I__5258 (
            .O(N__21931),
            .I(N__21605));
    ClkMux I__5257 (
            .O(N__21930),
            .I(N__21605));
    ClkMux I__5256 (
            .O(N__21929),
            .I(N__21605));
    ClkMux I__5255 (
            .O(N__21928),
            .I(N__21605));
    ClkMux I__5254 (
            .O(N__21927),
            .I(N__21605));
    ClkMux I__5253 (
            .O(N__21926),
            .I(N__21605));
    ClkMux I__5252 (
            .O(N__21925),
            .I(N__21605));
    ClkMux I__5251 (
            .O(N__21924),
            .I(N__21605));
    ClkMux I__5250 (
            .O(N__21923),
            .I(N__21605));
    ClkMux I__5249 (
            .O(N__21922),
            .I(N__21605));
    ClkMux I__5248 (
            .O(N__21921),
            .I(N__21605));
    ClkMux I__5247 (
            .O(N__21920),
            .I(N__21605));
    ClkMux I__5246 (
            .O(N__21919),
            .I(N__21605));
    ClkMux I__5245 (
            .O(N__21918),
            .I(N__21605));
    ClkMux I__5244 (
            .O(N__21917),
            .I(N__21605));
    ClkMux I__5243 (
            .O(N__21916),
            .I(N__21605));
    ClkMux I__5242 (
            .O(N__21915),
            .I(N__21605));
    ClkMux I__5241 (
            .O(N__21914),
            .I(N__21605));
    ClkMux I__5240 (
            .O(N__21913),
            .I(N__21605));
    ClkMux I__5239 (
            .O(N__21912),
            .I(N__21605));
    ClkMux I__5238 (
            .O(N__21911),
            .I(N__21605));
    ClkMux I__5237 (
            .O(N__21910),
            .I(N__21605));
    ClkMux I__5236 (
            .O(N__21909),
            .I(N__21605));
    ClkMux I__5235 (
            .O(N__21908),
            .I(N__21605));
    ClkMux I__5234 (
            .O(N__21907),
            .I(N__21605));
    ClkMux I__5233 (
            .O(N__21906),
            .I(N__21605));
    ClkMux I__5232 (
            .O(N__21905),
            .I(N__21605));
    ClkMux I__5231 (
            .O(N__21904),
            .I(N__21605));
    ClkMux I__5230 (
            .O(N__21903),
            .I(N__21605));
    ClkMux I__5229 (
            .O(N__21902),
            .I(N__21605));
    ClkMux I__5228 (
            .O(N__21901),
            .I(N__21605));
    ClkMux I__5227 (
            .O(N__21900),
            .I(N__21605));
    ClkMux I__5226 (
            .O(N__21899),
            .I(N__21605));
    ClkMux I__5225 (
            .O(N__21898),
            .I(N__21605));
    ClkMux I__5224 (
            .O(N__21897),
            .I(N__21605));
    ClkMux I__5223 (
            .O(N__21896),
            .I(N__21605));
    ClkMux I__5222 (
            .O(N__21895),
            .I(N__21605));
    ClkMux I__5221 (
            .O(N__21894),
            .I(N__21605));
    ClkMux I__5220 (
            .O(N__21893),
            .I(N__21605));
    ClkMux I__5219 (
            .O(N__21892),
            .I(N__21605));
    ClkMux I__5218 (
            .O(N__21891),
            .I(N__21605));
    ClkMux I__5217 (
            .O(N__21890),
            .I(N__21605));
    ClkMux I__5216 (
            .O(N__21889),
            .I(N__21605));
    ClkMux I__5215 (
            .O(N__21888),
            .I(N__21605));
    ClkMux I__5214 (
            .O(N__21887),
            .I(N__21605));
    ClkMux I__5213 (
            .O(N__21886),
            .I(N__21605));
    ClkMux I__5212 (
            .O(N__21885),
            .I(N__21605));
    ClkMux I__5211 (
            .O(N__21884),
            .I(N__21605));
    ClkMux I__5210 (
            .O(N__21883),
            .I(N__21605));
    ClkMux I__5209 (
            .O(N__21882),
            .I(N__21605));
    ClkMux I__5208 (
            .O(N__21881),
            .I(N__21605));
    ClkMux I__5207 (
            .O(N__21880),
            .I(N__21605));
    ClkMux I__5206 (
            .O(N__21879),
            .I(N__21605));
    ClkMux I__5205 (
            .O(N__21878),
            .I(N__21605));
    ClkMux I__5204 (
            .O(N__21877),
            .I(N__21605));
    ClkMux I__5203 (
            .O(N__21876),
            .I(N__21605));
    ClkMux I__5202 (
            .O(N__21875),
            .I(N__21605));
    ClkMux I__5201 (
            .O(N__21874),
            .I(N__21605));
    ClkMux I__5200 (
            .O(N__21873),
            .I(N__21605));
    ClkMux I__5199 (
            .O(N__21872),
            .I(N__21605));
    ClkMux I__5198 (
            .O(N__21871),
            .I(N__21605));
    ClkMux I__5197 (
            .O(N__21870),
            .I(N__21605));
    ClkMux I__5196 (
            .O(N__21869),
            .I(N__21605));
    ClkMux I__5195 (
            .O(N__21868),
            .I(N__21605));
    ClkMux I__5194 (
            .O(N__21867),
            .I(N__21605));
    ClkMux I__5193 (
            .O(N__21866),
            .I(N__21605));
    ClkMux I__5192 (
            .O(N__21865),
            .I(N__21605));
    ClkMux I__5191 (
            .O(N__21864),
            .I(N__21605));
    ClkMux I__5190 (
            .O(N__21863),
            .I(N__21605));
    ClkMux I__5189 (
            .O(N__21862),
            .I(N__21605));
    ClkMux I__5188 (
            .O(N__21861),
            .I(N__21605));
    ClkMux I__5187 (
            .O(N__21860),
            .I(N__21605));
    ClkMux I__5186 (
            .O(N__21859),
            .I(N__21605));
    ClkMux I__5185 (
            .O(N__21858),
            .I(N__21605));
    ClkMux I__5184 (
            .O(N__21857),
            .I(N__21605));
    ClkMux I__5183 (
            .O(N__21856),
            .I(N__21605));
    ClkMux I__5182 (
            .O(N__21855),
            .I(N__21605));
    ClkMux I__5181 (
            .O(N__21854),
            .I(N__21605));
    ClkMux I__5180 (
            .O(N__21853),
            .I(N__21605));
    ClkMux I__5179 (
            .O(N__21852),
            .I(N__21605));
    ClkMux I__5178 (
            .O(N__21851),
            .I(N__21605));
    ClkMux I__5177 (
            .O(N__21850),
            .I(N__21605));
    ClkMux I__5176 (
            .O(N__21849),
            .I(N__21605));
    ClkMux I__5175 (
            .O(N__21848),
            .I(N__21605));
    ClkMux I__5174 (
            .O(N__21847),
            .I(N__21605));
    ClkMux I__5173 (
            .O(N__21846),
            .I(N__21605));
    ClkMux I__5172 (
            .O(N__21845),
            .I(N__21605));
    ClkMux I__5171 (
            .O(N__21844),
            .I(N__21605));
    ClkMux I__5170 (
            .O(N__21843),
            .I(N__21605));
    ClkMux I__5169 (
            .O(N__21842),
            .I(N__21605));
    ClkMux I__5168 (
            .O(N__21841),
            .I(N__21605));
    ClkMux I__5167 (
            .O(N__21840),
            .I(N__21605));
    ClkMux I__5166 (
            .O(N__21839),
            .I(N__21605));
    ClkMux I__5165 (
            .O(N__21838),
            .I(N__21605));
    ClkMux I__5164 (
            .O(N__21837),
            .I(N__21605));
    ClkMux I__5163 (
            .O(N__21836),
            .I(N__21605));
    ClkMux I__5162 (
            .O(N__21835),
            .I(N__21605));
    ClkMux I__5161 (
            .O(N__21834),
            .I(N__21605));
    ClkMux I__5160 (
            .O(N__21833),
            .I(N__21605));
    ClkMux I__5159 (
            .O(N__21832),
            .I(N__21605));
    ClkMux I__5158 (
            .O(N__21831),
            .I(N__21605));
    ClkMux I__5157 (
            .O(N__21830),
            .I(N__21605));
    ClkMux I__5156 (
            .O(N__21829),
            .I(N__21605));
    ClkMux I__5155 (
            .O(N__21828),
            .I(N__21605));
    ClkMux I__5154 (
            .O(N__21827),
            .I(N__21605));
    ClkMux I__5153 (
            .O(N__21826),
            .I(N__21605));
    ClkMux I__5152 (
            .O(N__21825),
            .I(N__21605));
    ClkMux I__5151 (
            .O(N__21824),
            .I(N__21605));
    GlobalMux I__5150 (
            .O(N__21605),
            .I(N__21602));
    gio2CtrlBuf I__5149 (
            .O(N__21602),
            .I(CLK_c_g));
    CEMux I__5148 (
            .O(N__21599),
            .I(N__21542));
    CEMux I__5147 (
            .O(N__21598),
            .I(N__21542));
    CEMux I__5146 (
            .O(N__21597),
            .I(N__21542));
    CEMux I__5145 (
            .O(N__21596),
            .I(N__21542));
    CEMux I__5144 (
            .O(N__21595),
            .I(N__21542));
    CEMux I__5143 (
            .O(N__21594),
            .I(N__21542));
    CEMux I__5142 (
            .O(N__21593),
            .I(N__21542));
    CEMux I__5141 (
            .O(N__21592),
            .I(N__21542));
    CEMux I__5140 (
            .O(N__21591),
            .I(N__21542));
    CEMux I__5139 (
            .O(N__21590),
            .I(N__21542));
    CEMux I__5138 (
            .O(N__21589),
            .I(N__21542));
    CEMux I__5137 (
            .O(N__21588),
            .I(N__21542));
    CEMux I__5136 (
            .O(N__21587),
            .I(N__21542));
    CEMux I__5135 (
            .O(N__21586),
            .I(N__21542));
    CEMux I__5134 (
            .O(N__21585),
            .I(N__21542));
    CEMux I__5133 (
            .O(N__21584),
            .I(N__21542));
    CEMux I__5132 (
            .O(N__21583),
            .I(N__21542));
    CEMux I__5131 (
            .O(N__21582),
            .I(N__21542));
    CEMux I__5130 (
            .O(N__21581),
            .I(N__21542));
    GlobalMux I__5129 (
            .O(N__21542),
            .I(N__21539));
    gio2CtrlBuf I__5128 (
            .O(N__21539),
            .I(\c0.data_in_frame_0__0_sqmuxa_g ));
    InMux I__5127 (
            .O(N__21536),
            .I(N__21533));
    LocalMux I__5126 (
            .O(N__21533),
            .I(N__21530));
    Odrv12 I__5125 (
            .O(N__21530),
            .I(\c0.rx.r_Rx_Bytece_1_2 ));
    CascadeMux I__5124 (
            .O(N__21527),
            .I(N__21523));
    InMux I__5123 (
            .O(N__21526),
            .I(N__21520));
    InMux I__5122 (
            .O(N__21523),
            .I(N__21517));
    LocalMux I__5121 (
            .O(N__21520),
            .I(\c0.rx_data_2 ));
    LocalMux I__5120 (
            .O(N__21517),
            .I(\c0.rx_data_2 ));
    CascadeMux I__5119 (
            .O(N__21512),
            .I(\c0.rx.r_Rx_Bytece_1_4_cascade_ ));
    InMux I__5118 (
            .O(N__21509),
            .I(N__21505));
    InMux I__5117 (
            .O(N__21508),
            .I(N__21502));
    LocalMux I__5116 (
            .O(N__21505),
            .I(\c0.rx_data_4 ));
    LocalMux I__5115 (
            .O(N__21502),
            .I(\c0.rx_data_4 ));
    InMux I__5114 (
            .O(N__21497),
            .I(N__21491));
    InMux I__5113 (
            .O(N__21496),
            .I(N__21486));
    InMux I__5112 (
            .O(N__21495),
            .I(N__21486));
    InMux I__5111 (
            .O(N__21494),
            .I(N__21482));
    LocalMux I__5110 (
            .O(N__21491),
            .I(N__21478));
    LocalMux I__5109 (
            .O(N__21486),
            .I(N__21475));
    InMux I__5108 (
            .O(N__21485),
            .I(N__21472));
    LocalMux I__5107 (
            .O(N__21482),
            .I(N__21468));
    InMux I__5106 (
            .O(N__21481),
            .I(N__21465));
    Span4Mux_v I__5105 (
            .O(N__21478),
            .I(N__21462));
    Span4Mux_h I__5104 (
            .O(N__21475),
            .I(N__21456));
    LocalMux I__5103 (
            .O(N__21472),
            .I(N__21456));
    InMux I__5102 (
            .O(N__21471),
            .I(N__21453));
    Span4Mux_h I__5101 (
            .O(N__21468),
            .I(N__21447));
    LocalMux I__5100 (
            .O(N__21465),
            .I(N__21447));
    Span4Mux_h I__5099 (
            .O(N__21462),
            .I(N__21444));
    InMux I__5098 (
            .O(N__21461),
            .I(N__21441));
    Span4Mux_h I__5097 (
            .O(N__21456),
            .I(N__21436));
    LocalMux I__5096 (
            .O(N__21453),
            .I(N__21436));
    InMux I__5095 (
            .O(N__21452),
            .I(N__21433));
    Span4Mux_h I__5094 (
            .O(N__21447),
            .I(N__21430));
    Span4Mux_h I__5093 (
            .O(N__21444),
            .I(N__21425));
    LocalMux I__5092 (
            .O(N__21441),
            .I(N__21425));
    Span4Mux_h I__5091 (
            .O(N__21436),
            .I(N__21422));
    LocalMux I__5090 (
            .O(N__21433),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__5089 (
            .O(N__21430),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__5088 (
            .O(N__21425),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__5087 (
            .O(N__21422),
            .I(\c0.rx.r_Bit_IndexZ0Z_2 ));
    InMux I__5086 (
            .O(N__21413),
            .I(N__21407));
    CascadeMux I__5085 (
            .O(N__21412),
            .I(N__21404));
    InMux I__5084 (
            .O(N__21411),
            .I(N__21400));
    InMux I__5083 (
            .O(N__21410),
            .I(N__21397));
    LocalMux I__5082 (
            .O(N__21407),
            .I(N__21392));
    InMux I__5081 (
            .O(N__21404),
            .I(N__21385));
    InMux I__5080 (
            .O(N__21403),
            .I(N__21385));
    LocalMux I__5079 (
            .O(N__21400),
            .I(N__21382));
    LocalMux I__5078 (
            .O(N__21397),
            .I(N__21379));
    InMux I__5077 (
            .O(N__21396),
            .I(N__21376));
    InMux I__5076 (
            .O(N__21395),
            .I(N__21373));
    Span4Mux_v I__5075 (
            .O(N__21392),
            .I(N__21370));
    InMux I__5074 (
            .O(N__21391),
            .I(N__21367));
    CascadeMux I__5073 (
            .O(N__21390),
            .I(N__21364));
    LocalMux I__5072 (
            .O(N__21385),
            .I(N__21360));
    Span4Mux_h I__5071 (
            .O(N__21382),
            .I(N__21357));
    Span4Mux_h I__5070 (
            .O(N__21379),
            .I(N__21354));
    LocalMux I__5069 (
            .O(N__21376),
            .I(N__21349));
    LocalMux I__5068 (
            .O(N__21373),
            .I(N__21349));
    Span4Mux_h I__5067 (
            .O(N__21370),
            .I(N__21344));
    LocalMux I__5066 (
            .O(N__21367),
            .I(N__21344));
    InMux I__5065 (
            .O(N__21364),
            .I(N__21339));
    InMux I__5064 (
            .O(N__21363),
            .I(N__21339));
    Odrv12 I__5063 (
            .O(N__21360),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__5062 (
            .O(N__21357),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__5061 (
            .O(N__21354),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__5060 (
            .O(N__21349),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__5059 (
            .O(N__21344),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__5058 (
            .O(N__21339),
            .I(\c0.rx.r_Bit_IndexZ0Z_1 ));
    InMux I__5057 (
            .O(N__21326),
            .I(N__21319));
    InMux I__5056 (
            .O(N__21325),
            .I(N__21319));
    InMux I__5055 (
            .O(N__21324),
            .I(N__21316));
    LocalMux I__5054 (
            .O(N__21319),
            .I(N__21312));
    LocalMux I__5053 (
            .O(N__21316),
            .I(N__21309));
    InMux I__5052 (
            .O(N__21315),
            .I(N__21305));
    Span4Mux_h I__5051 (
            .O(N__21312),
            .I(N__21299));
    Span4Mux_v I__5050 (
            .O(N__21309),
            .I(N__21299));
    InMux I__5049 (
            .O(N__21308),
            .I(N__21296));
    LocalMux I__5048 (
            .O(N__21305),
            .I(N__21290));
    InMux I__5047 (
            .O(N__21304),
            .I(N__21287));
    Span4Mux_h I__5046 (
            .O(N__21299),
            .I(N__21282));
    LocalMux I__5045 (
            .O(N__21296),
            .I(N__21282));
    InMux I__5044 (
            .O(N__21295),
            .I(N__21279));
    InMux I__5043 (
            .O(N__21294),
            .I(N__21274));
    InMux I__5042 (
            .O(N__21293),
            .I(N__21271));
    Span4Mux_v I__5041 (
            .O(N__21290),
            .I(N__21266));
    LocalMux I__5040 (
            .O(N__21287),
            .I(N__21266));
    Span4Mux_h I__5039 (
            .O(N__21282),
            .I(N__21261));
    LocalMux I__5038 (
            .O(N__21279),
            .I(N__21261));
    InMux I__5037 (
            .O(N__21278),
            .I(N__21256));
    InMux I__5036 (
            .O(N__21277),
            .I(N__21256));
    LocalMux I__5035 (
            .O(N__21274),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__5034 (
            .O(N__21271),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__5033 (
            .O(N__21266),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__5032 (
            .O(N__21261),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__5031 (
            .O(N__21256),
            .I(\c0.rx.r_Bit_IndexZ0Z_0 ));
    InMux I__5030 (
            .O(N__21245),
            .I(N__21232));
    InMux I__5029 (
            .O(N__21244),
            .I(N__21232));
    InMux I__5028 (
            .O(N__21243),
            .I(N__21232));
    InMux I__5027 (
            .O(N__21242),
            .I(N__21232));
    CascadeMux I__5026 (
            .O(N__21241),
            .I(N__21229));
    LocalMux I__5025 (
            .O(N__21232),
            .I(N__21224));
    InMux I__5024 (
            .O(N__21229),
            .I(N__21219));
    InMux I__5023 (
            .O(N__21228),
            .I(N__21219));
    InMux I__5022 (
            .O(N__21227),
            .I(N__21215));
    Span4Mux_v I__5021 (
            .O(N__21224),
            .I(N__21210));
    LocalMux I__5020 (
            .O(N__21219),
            .I(N__21207));
    InMux I__5019 (
            .O(N__21218),
            .I(N__21204));
    LocalMux I__5018 (
            .O(N__21215),
            .I(N__21201));
    InMux I__5017 (
            .O(N__21214),
            .I(N__21198));
    CascadeMux I__5016 (
            .O(N__21213),
            .I(N__21195));
    Sp12to4 I__5015 (
            .O(N__21210),
            .I(N__21190));
    Span4Mux_v I__5014 (
            .O(N__21207),
            .I(N__21187));
    LocalMux I__5013 (
            .O(N__21204),
            .I(N__21184));
    Span4Mux_v I__5012 (
            .O(N__21201),
            .I(N__21179));
    LocalMux I__5011 (
            .O(N__21198),
            .I(N__21179));
    InMux I__5010 (
            .O(N__21195),
            .I(N__21174));
    InMux I__5009 (
            .O(N__21194),
            .I(N__21174));
    CascadeMux I__5008 (
            .O(N__21193),
            .I(N__21171));
    Span12Mux_h I__5007 (
            .O(N__21190),
            .I(N__21164));
    Sp12to4 I__5006 (
            .O(N__21187),
            .I(N__21164));
    Span12Mux_v I__5005 (
            .O(N__21184),
            .I(N__21164));
    Span4Mux_h I__5004 (
            .O(N__21179),
            .I(N__21159));
    LocalMux I__5003 (
            .O(N__21174),
            .I(N__21159));
    InMux I__5002 (
            .O(N__21171),
            .I(N__21156));
    Odrv12 I__5001 (
            .O(N__21164),
            .I(\c0.rx.r_Rx_DataZ0 ));
    Odrv4 I__5000 (
            .O(N__21159),
            .I(\c0.rx.r_Rx_DataZ0 ));
    LocalMux I__4999 (
            .O(N__21156),
            .I(\c0.rx.r_Rx_DataZ0 ));
    CascadeMux I__4998 (
            .O(N__21149),
            .I(\c0.rx.r_Rx_Bytece_1_0_cascade_ ));
    InMux I__4997 (
            .O(N__21146),
            .I(N__21138));
    InMux I__4996 (
            .O(N__21145),
            .I(N__21133));
    InMux I__4995 (
            .O(N__21144),
            .I(N__21123));
    InMux I__4994 (
            .O(N__21143),
            .I(N__21123));
    InMux I__4993 (
            .O(N__21142),
            .I(N__21123));
    InMux I__4992 (
            .O(N__21141),
            .I(N__21123));
    LocalMux I__4991 (
            .O(N__21138),
            .I(N__21119));
    InMux I__4990 (
            .O(N__21137),
            .I(N__21114));
    InMux I__4989 (
            .O(N__21136),
            .I(N__21114));
    LocalMux I__4988 (
            .O(N__21133),
            .I(N__21111));
    InMux I__4987 (
            .O(N__21132),
            .I(N__21108));
    LocalMux I__4986 (
            .O(N__21123),
            .I(N__21105));
    InMux I__4985 (
            .O(N__21122),
            .I(N__21102));
    Span4Mux_h I__4984 (
            .O(N__21119),
            .I(N__21097));
    LocalMux I__4983 (
            .O(N__21114),
            .I(N__21097));
    Span4Mux_h I__4982 (
            .O(N__21111),
            .I(N__21093));
    LocalMux I__4981 (
            .O(N__21108),
            .I(N__21086));
    Span12Mux_h I__4980 (
            .O(N__21105),
            .I(N__21086));
    LocalMux I__4979 (
            .O(N__21102),
            .I(N__21086));
    Span4Mux_h I__4978 (
            .O(N__21097),
            .I(N__21083));
    InMux I__4977 (
            .O(N__21096),
            .I(N__21080));
    Odrv4 I__4976 (
            .O(N__21093),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    Odrv12 I__4975 (
            .O(N__21086),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    Odrv4 I__4974 (
            .O(N__21083),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    LocalMux I__4973 (
            .O(N__21080),
            .I(\c0.rx.r_Rx_Byte_1_sqmuxa ));
    InMux I__4972 (
            .O(N__21071),
            .I(N__21067));
    InMux I__4971 (
            .O(N__21070),
            .I(N__21064));
    LocalMux I__4970 (
            .O(N__21067),
            .I(\c0.rx_data_0 ));
    LocalMux I__4969 (
            .O(N__21064),
            .I(\c0.rx_data_0 ));
    InMux I__4968 (
            .O(N__21059),
            .I(N__21055));
    InMux I__4967 (
            .O(N__21058),
            .I(N__21052));
    LocalMux I__4966 (
            .O(N__21055),
            .I(N__21049));
    LocalMux I__4965 (
            .O(N__21052),
            .I(N__21046));
    Odrv12 I__4964 (
            .O(N__21049),
            .I(\c0.un1_byte_transmit_counter2_1_ac0_3_out ));
    Odrv4 I__4963 (
            .O(N__21046),
            .I(\c0.un1_byte_transmit_counter2_1_ac0_3_out ));
    InMux I__4962 (
            .O(N__21041),
            .I(N__21034));
    InMux I__4961 (
            .O(N__21040),
            .I(N__21034));
    InMux I__4960 (
            .O(N__21039),
            .I(N__21029));
    LocalMux I__4959 (
            .O(N__21034),
            .I(N__21026));
    InMux I__4958 (
            .O(N__21033),
            .I(N__21023));
    InMux I__4957 (
            .O(N__21032),
            .I(N__21020));
    LocalMux I__4956 (
            .O(N__21029),
            .I(\c0.byte_transmit_counter2Z0Z_3 ));
    Odrv4 I__4955 (
            .O(N__21026),
            .I(\c0.byte_transmit_counter2Z0Z_3 ));
    LocalMux I__4954 (
            .O(N__21023),
            .I(\c0.byte_transmit_counter2Z0Z_3 ));
    LocalMux I__4953 (
            .O(N__21020),
            .I(\c0.byte_transmit_counter2Z0Z_3 ));
    InMux I__4952 (
            .O(N__21011),
            .I(N__21006));
    InMux I__4951 (
            .O(N__21010),
            .I(N__21002));
    InMux I__4950 (
            .O(N__21009),
            .I(N__20999));
    LocalMux I__4949 (
            .O(N__21006),
            .I(N__20996));
    InMux I__4948 (
            .O(N__21005),
            .I(N__20993));
    LocalMux I__4947 (
            .O(N__21002),
            .I(\c0.byte_transmit_counter2Z0Z_4 ));
    LocalMux I__4946 (
            .O(N__20999),
            .I(\c0.byte_transmit_counter2Z0Z_4 ));
    Odrv4 I__4945 (
            .O(N__20996),
            .I(\c0.byte_transmit_counter2Z0Z_4 ));
    LocalMux I__4944 (
            .O(N__20993),
            .I(\c0.byte_transmit_counter2Z0Z_4 ));
    CascadeMux I__4943 (
            .O(N__20984),
            .I(N__20980));
    InMux I__4942 (
            .O(N__20983),
            .I(N__20975));
    InMux I__4941 (
            .O(N__20980),
            .I(N__20975));
    LocalMux I__4940 (
            .O(N__20975),
            .I(N__20972));
    Odrv4 I__4939 (
            .O(N__20972),
            .I(\c0.un1_byte_transmit_counter2_1_ac0_7_out_0 ));
    InMux I__4938 (
            .O(N__20969),
            .I(N__20966));
    LocalMux I__4937 (
            .O(N__20966),
            .I(\c0.tx2_data_1_iv_5_4 ));
    InMux I__4936 (
            .O(N__20963),
            .I(N__20960));
    LocalMux I__4935 (
            .O(N__20960),
            .I(\c0.tx2_data_1_0_i_1_4 ));
    CascadeMux I__4934 (
            .O(N__20957),
            .I(N__20954));
    InMux I__4933 (
            .O(N__20954),
            .I(N__20951));
    LocalMux I__4932 (
            .O(N__20951),
            .I(N__20948));
    Span4Mux_h I__4931 (
            .O(N__20948),
            .I(N__20945));
    Odrv4 I__4930 (
            .O(N__20945),
            .I(\c0.tx2_data_1_0_i_1_0_4 ));
    InMux I__4929 (
            .O(N__20942),
            .I(N__20934));
    InMux I__4928 (
            .O(N__20941),
            .I(N__20934));
    CascadeMux I__4927 (
            .O(N__20940),
            .I(N__20929));
    InMux I__4926 (
            .O(N__20939),
            .I(N__20916));
    LocalMux I__4925 (
            .O(N__20934),
            .I(N__20913));
    InMux I__4924 (
            .O(N__20933),
            .I(N__20908));
    InMux I__4923 (
            .O(N__20932),
            .I(N__20908));
    InMux I__4922 (
            .O(N__20929),
            .I(N__20903));
    InMux I__4921 (
            .O(N__20928),
            .I(N__20903));
    InMux I__4920 (
            .O(N__20927),
            .I(N__20896));
    InMux I__4919 (
            .O(N__20926),
            .I(N__20896));
    InMux I__4918 (
            .O(N__20925),
            .I(N__20891));
    InMux I__4917 (
            .O(N__20924),
            .I(N__20891));
    InMux I__4916 (
            .O(N__20923),
            .I(N__20884));
    InMux I__4915 (
            .O(N__20922),
            .I(N__20884));
    InMux I__4914 (
            .O(N__20921),
            .I(N__20884));
    InMux I__4913 (
            .O(N__20920),
            .I(N__20879));
    InMux I__4912 (
            .O(N__20919),
            .I(N__20879));
    LocalMux I__4911 (
            .O(N__20916),
            .I(N__20875));
    Span4Mux_h I__4910 (
            .O(N__20913),
            .I(N__20868));
    LocalMux I__4909 (
            .O(N__20908),
            .I(N__20868));
    LocalMux I__4908 (
            .O(N__20903),
            .I(N__20868));
    InMux I__4907 (
            .O(N__20902),
            .I(N__20865));
    CascadeMux I__4906 (
            .O(N__20901),
            .I(N__20862));
    LocalMux I__4905 (
            .O(N__20896),
            .I(N__20853));
    LocalMux I__4904 (
            .O(N__20891),
            .I(N__20853));
    LocalMux I__4903 (
            .O(N__20884),
            .I(N__20850));
    LocalMux I__4902 (
            .O(N__20879),
            .I(N__20847));
    InMux I__4901 (
            .O(N__20878),
            .I(N__20840));
    Span4Mux_v I__4900 (
            .O(N__20875),
            .I(N__20833));
    Span4Mux_v I__4899 (
            .O(N__20868),
            .I(N__20833));
    LocalMux I__4898 (
            .O(N__20865),
            .I(N__20833));
    InMux I__4897 (
            .O(N__20862),
            .I(N__20826));
    InMux I__4896 (
            .O(N__20861),
            .I(N__20826));
    InMux I__4895 (
            .O(N__20860),
            .I(N__20821));
    InMux I__4894 (
            .O(N__20859),
            .I(N__20821));
    InMux I__4893 (
            .O(N__20858),
            .I(N__20818));
    Span4Mux_v I__4892 (
            .O(N__20853),
            .I(N__20813));
    Span4Mux_v I__4891 (
            .O(N__20850),
            .I(N__20813));
    Span4Mux_v I__4890 (
            .O(N__20847),
            .I(N__20810));
    InMux I__4889 (
            .O(N__20846),
            .I(N__20803));
    InMux I__4888 (
            .O(N__20845),
            .I(N__20803));
    InMux I__4887 (
            .O(N__20844),
            .I(N__20803));
    InMux I__4886 (
            .O(N__20843),
            .I(N__20800));
    LocalMux I__4885 (
            .O(N__20840),
            .I(N__20795));
    Span4Mux_h I__4884 (
            .O(N__20833),
            .I(N__20795));
    InMux I__4883 (
            .O(N__20832),
            .I(N__20790));
    InMux I__4882 (
            .O(N__20831),
            .I(N__20790));
    LocalMux I__4881 (
            .O(N__20826),
            .I(N__20787));
    LocalMux I__4880 (
            .O(N__20821),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    LocalMux I__4879 (
            .O(N__20818),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    Odrv4 I__4878 (
            .O(N__20813),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    Odrv4 I__4877 (
            .O(N__20810),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    LocalMux I__4876 (
            .O(N__20803),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    LocalMux I__4875 (
            .O(N__20800),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    Odrv4 I__4874 (
            .O(N__20795),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    LocalMux I__4873 (
            .O(N__20790),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    Odrv12 I__4872 (
            .O(N__20787),
            .I(\c0.byte_transmit_counter2Z0Z_1 ));
    CascadeMux I__4871 (
            .O(N__20768),
            .I(N__20765));
    InMux I__4870 (
            .O(N__20765),
            .I(N__20762));
    LocalMux I__4869 (
            .O(N__20762),
            .I(N__20759));
    Span4Mux_v I__4868 (
            .O(N__20759),
            .I(N__20756));
    Span4Mux_h I__4867 (
            .O(N__20756),
            .I(N__20753));
    Odrv4 I__4866 (
            .O(N__20753),
            .I(\c0.tx2.r_Tx_DataZ0Z_4 ));
    CEMux I__4865 (
            .O(N__20750),
            .I(N__20746));
    InMux I__4864 (
            .O(N__20749),
            .I(N__20742));
    LocalMux I__4863 (
            .O(N__20746),
            .I(N__20738));
    CEMux I__4862 (
            .O(N__20745),
            .I(N__20735));
    LocalMux I__4861 (
            .O(N__20742),
            .I(N__20730));
    CEMux I__4860 (
            .O(N__20741),
            .I(N__20727));
    Span4Mux_v I__4859 (
            .O(N__20738),
            .I(N__20722));
    LocalMux I__4858 (
            .O(N__20735),
            .I(N__20722));
    CEMux I__4857 (
            .O(N__20734),
            .I(N__20719));
    CEMux I__4856 (
            .O(N__20733),
            .I(N__20716));
    Span4Mux_v I__4855 (
            .O(N__20730),
            .I(N__20710));
    LocalMux I__4854 (
            .O(N__20727),
            .I(N__20710));
    Span4Mux_h I__4853 (
            .O(N__20722),
            .I(N__20707));
    LocalMux I__4852 (
            .O(N__20719),
            .I(N__20704));
    LocalMux I__4851 (
            .O(N__20716),
            .I(N__20701));
    CascadeMux I__4850 (
            .O(N__20715),
            .I(N__20698));
    Span4Mux_v I__4849 (
            .O(N__20710),
            .I(N__20695));
    Span4Mux_h I__4848 (
            .O(N__20707),
            .I(N__20690));
    Span4Mux_h I__4847 (
            .O(N__20704),
            .I(N__20690));
    Span4Mux_v I__4846 (
            .O(N__20701),
            .I(N__20687));
    InMux I__4845 (
            .O(N__20698),
            .I(N__20684));
    Span4Mux_h I__4844 (
            .O(N__20695),
            .I(N__20681));
    Sp12to4 I__4843 (
            .O(N__20690),
            .I(N__20678));
    Span4Mux_h I__4842 (
            .O(N__20687),
            .I(N__20675));
    LocalMux I__4841 (
            .O(N__20684),
            .I(\c0.tx2.r_Tx_Data_0_sqmuxa ));
    Odrv4 I__4840 (
            .O(N__20681),
            .I(\c0.tx2.r_Tx_Data_0_sqmuxa ));
    Odrv12 I__4839 (
            .O(N__20678),
            .I(\c0.tx2.r_Tx_Data_0_sqmuxa ));
    Odrv4 I__4838 (
            .O(N__20675),
            .I(\c0.tx2.r_Tx_Data_0_sqmuxa ));
    InMux I__4837 (
            .O(N__20666),
            .I(N__20662));
    InMux I__4836 (
            .O(N__20665),
            .I(N__20659));
    LocalMux I__4835 (
            .O(N__20662),
            .I(N__20656));
    LocalMux I__4834 (
            .O(N__20659),
            .I(N__20653));
    Span12Mux_v I__4833 (
            .O(N__20656),
            .I(N__20650));
    Span4Mux_h I__4832 (
            .O(N__20653),
            .I(N__20647));
    Odrv12 I__4831 (
            .O(N__20650),
            .I(\c0.data_in_5_Z0Z_7 ));
    Odrv4 I__4830 (
            .O(N__20647),
            .I(\c0.data_in_5_Z0Z_7 ));
    InMux I__4829 (
            .O(N__20642),
            .I(N__20638));
    CascadeMux I__4828 (
            .O(N__20641),
            .I(N__20635));
    LocalMux I__4827 (
            .O(N__20638),
            .I(N__20632));
    InMux I__4826 (
            .O(N__20635),
            .I(N__20628));
    Span12Mux_h I__4825 (
            .O(N__20632),
            .I(N__20625));
    InMux I__4824 (
            .O(N__20631),
            .I(N__20622));
    LocalMux I__4823 (
            .O(N__20628),
            .I(N__20619));
    Odrv12 I__4822 (
            .O(N__20625),
            .I(\c0.data_in_6_Z0Z_3 ));
    LocalMux I__4821 (
            .O(N__20622),
            .I(\c0.data_in_6_Z0Z_3 ));
    Odrv12 I__4820 (
            .O(N__20619),
            .I(\c0.data_in_6_Z0Z_3 ));
    InMux I__4819 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__4818 (
            .O(N__20609),
            .I(N__20606));
    Span4Mux_h I__4817 (
            .O(N__20606),
            .I(N__20603));
    Odrv4 I__4816 (
            .O(N__20603),
            .I(\c0.data_in_frame_6_Z0Z_3 ));
    InMux I__4815 (
            .O(N__20600),
            .I(N__20597));
    LocalMux I__4814 (
            .O(N__20597),
            .I(N__20594));
    Span4Mux_h I__4813 (
            .O(N__20594),
            .I(N__20591));
    Odrv4 I__4812 (
            .O(N__20591),
            .I(\c0.tx2_data_1_0_i_1_6 ));
    InMux I__4811 (
            .O(N__20588),
            .I(N__20585));
    LocalMux I__4810 (
            .O(N__20585),
            .I(N__20580));
    InMux I__4809 (
            .O(N__20584),
            .I(N__20577));
    InMux I__4808 (
            .O(N__20583),
            .I(N__20574));
    Span4Mux_h I__4807 (
            .O(N__20580),
            .I(N__20571));
    LocalMux I__4806 (
            .O(N__20577),
            .I(\c0.data_in_6_Z0Z_6 ));
    LocalMux I__4805 (
            .O(N__20574),
            .I(\c0.data_in_6_Z0Z_6 ));
    Odrv4 I__4804 (
            .O(N__20571),
            .I(\c0.data_in_6_Z0Z_6 ));
    CascadeMux I__4803 (
            .O(N__20564),
            .I(N__20561));
    InMux I__4802 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__4801 (
            .O(N__20558),
            .I(\c0.data_in_frame_6_Z0Z_6 ));
    InMux I__4800 (
            .O(N__20555),
            .I(N__20552));
    LocalMux I__4799 (
            .O(N__20552),
            .I(N__20549));
    Span4Mux_v I__4798 (
            .O(N__20549),
            .I(N__20546));
    Span4Mux_h I__4797 (
            .O(N__20546),
            .I(N__20542));
    InMux I__4796 (
            .O(N__20545),
            .I(N__20539));
    Odrv4 I__4795 (
            .O(N__20542),
            .I(\c0.data_in_4_Z0Z_6 ));
    LocalMux I__4794 (
            .O(N__20539),
            .I(\c0.data_in_4_Z0Z_6 ));
    InMux I__4793 (
            .O(N__20534),
            .I(N__20529));
    InMux I__4792 (
            .O(N__20533),
            .I(N__20525));
    InMux I__4791 (
            .O(N__20532),
            .I(N__20522));
    LocalMux I__4790 (
            .O(N__20529),
            .I(N__20519));
    InMux I__4789 (
            .O(N__20528),
            .I(N__20516));
    LocalMux I__4788 (
            .O(N__20525),
            .I(N__20508));
    LocalMux I__4787 (
            .O(N__20522),
            .I(N__20508));
    Span4Mux_h I__4786 (
            .O(N__20519),
            .I(N__20508));
    LocalMux I__4785 (
            .O(N__20516),
            .I(N__20501));
    InMux I__4784 (
            .O(N__20515),
            .I(N__20498));
    Span4Mux_v I__4783 (
            .O(N__20508),
            .I(N__20495));
    InMux I__4782 (
            .O(N__20507),
            .I(N__20486));
    InMux I__4781 (
            .O(N__20506),
            .I(N__20486));
    InMux I__4780 (
            .O(N__20505),
            .I(N__20486));
    InMux I__4779 (
            .O(N__20504),
            .I(N__20486));
    Span4Mux_v I__4778 (
            .O(N__20501),
            .I(N__20483));
    LocalMux I__4777 (
            .O(N__20498),
            .I(\c0.d_4_38 ));
    Odrv4 I__4776 (
            .O(N__20495),
            .I(\c0.d_4_38 ));
    LocalMux I__4775 (
            .O(N__20486),
            .I(\c0.d_4_38 ));
    Odrv4 I__4774 (
            .O(N__20483),
            .I(\c0.d_4_38 ));
    InMux I__4773 (
            .O(N__20474),
            .I(N__20471));
    LocalMux I__4772 (
            .O(N__20471),
            .I(N__20465));
    InMux I__4771 (
            .O(N__20470),
            .I(N__20462));
    InMux I__4770 (
            .O(N__20469),
            .I(N__20457));
    InMux I__4769 (
            .O(N__20468),
            .I(N__20457));
    Odrv4 I__4768 (
            .O(N__20465),
            .I(\c0.d_4_5 ));
    LocalMux I__4767 (
            .O(N__20462),
            .I(\c0.d_4_5 ));
    LocalMux I__4766 (
            .O(N__20457),
            .I(\c0.d_4_5 ));
    CascadeMux I__4765 (
            .O(N__20450),
            .I(N__20447));
    InMux I__4764 (
            .O(N__20447),
            .I(N__20444));
    LocalMux I__4763 (
            .O(N__20444),
            .I(N__20439));
    InMux I__4762 (
            .O(N__20443),
            .I(N__20434));
    InMux I__4761 (
            .O(N__20442),
            .I(N__20434));
    Span4Mux_v I__4760 (
            .O(N__20439),
            .I(N__20431));
    LocalMux I__4759 (
            .O(N__20434),
            .I(N__20427));
    Span4Mux_h I__4758 (
            .O(N__20431),
            .I(N__20424));
    InMux I__4757 (
            .O(N__20430),
            .I(N__20421));
    Span4Mux_h I__4756 (
            .O(N__20427),
            .I(N__20418));
    Odrv4 I__4755 (
            .O(N__20424),
            .I(\c0.d_4_21 ));
    LocalMux I__4754 (
            .O(N__20421),
            .I(\c0.d_4_21 ));
    Odrv4 I__4753 (
            .O(N__20418),
            .I(\c0.d_4_21 ));
    CascadeMux I__4752 (
            .O(N__20411),
            .I(N__20404));
    InMux I__4751 (
            .O(N__20410),
            .I(N__20399));
    InMux I__4750 (
            .O(N__20409),
            .I(N__20399));
    InMux I__4749 (
            .O(N__20408),
            .I(N__20392));
    InMux I__4748 (
            .O(N__20407),
            .I(N__20392));
    InMux I__4747 (
            .O(N__20404),
            .I(N__20392));
    LocalMux I__4746 (
            .O(N__20399),
            .I(N__20385));
    LocalMux I__4745 (
            .O(N__20392),
            .I(N__20382));
    InMux I__4744 (
            .O(N__20391),
            .I(N__20375));
    InMux I__4743 (
            .O(N__20390),
            .I(N__20375));
    InMux I__4742 (
            .O(N__20389),
            .I(N__20375));
    InMux I__4741 (
            .O(N__20388),
            .I(N__20372));
    Span4Mux_h I__4740 (
            .O(N__20385),
            .I(N__20365));
    Span4Mux_h I__4739 (
            .O(N__20382),
            .I(N__20365));
    LocalMux I__4738 (
            .O(N__20375),
            .I(N__20365));
    LocalMux I__4737 (
            .O(N__20372),
            .I(\c0.N_203 ));
    Odrv4 I__4736 (
            .O(N__20365),
            .I(\c0.N_203 ));
    CascadeMux I__4735 (
            .O(N__20360),
            .I(\c0.tx2_data_1_iv_5_1_5_cascade_ ));
    InMux I__4734 (
            .O(N__20357),
            .I(N__20349));
    InMux I__4733 (
            .O(N__20356),
            .I(N__20349));
    InMux I__4732 (
            .O(N__20355),
            .I(N__20346));
    InMux I__4731 (
            .O(N__20354),
            .I(N__20335));
    LocalMux I__4730 (
            .O(N__20349),
            .I(N__20329));
    LocalMux I__4729 (
            .O(N__20346),
            .I(N__20321));
    InMux I__4728 (
            .O(N__20345),
            .I(N__20312));
    InMux I__4727 (
            .O(N__20344),
            .I(N__20312));
    InMux I__4726 (
            .O(N__20343),
            .I(N__20312));
    InMux I__4725 (
            .O(N__20342),
            .I(N__20312));
    InMux I__4724 (
            .O(N__20341),
            .I(N__20309));
    InMux I__4723 (
            .O(N__20340),
            .I(N__20306));
    InMux I__4722 (
            .O(N__20339),
            .I(N__20301));
    InMux I__4721 (
            .O(N__20338),
            .I(N__20301));
    LocalMux I__4720 (
            .O(N__20335),
            .I(N__20298));
    InMux I__4719 (
            .O(N__20334),
            .I(N__20295));
    InMux I__4718 (
            .O(N__20333),
            .I(N__20290));
    InMux I__4717 (
            .O(N__20332),
            .I(N__20290));
    Span4Mux_h I__4716 (
            .O(N__20329),
            .I(N__20286));
    InMux I__4715 (
            .O(N__20328),
            .I(N__20283));
    InMux I__4714 (
            .O(N__20327),
            .I(N__20280));
    CascadeMux I__4713 (
            .O(N__20326),
            .I(N__20271));
    CascadeMux I__4712 (
            .O(N__20325),
            .I(N__20267));
    CascadeMux I__4711 (
            .O(N__20324),
            .I(N__20264));
    Span4Mux_v I__4710 (
            .O(N__20321),
            .I(N__20255));
    LocalMux I__4709 (
            .O(N__20312),
            .I(N__20255));
    LocalMux I__4708 (
            .O(N__20309),
            .I(N__20255));
    LocalMux I__4707 (
            .O(N__20306),
            .I(N__20255));
    LocalMux I__4706 (
            .O(N__20301),
            .I(N__20252));
    Span4Mux_v I__4705 (
            .O(N__20298),
            .I(N__20245));
    LocalMux I__4704 (
            .O(N__20295),
            .I(N__20245));
    LocalMux I__4703 (
            .O(N__20290),
            .I(N__20245));
    InMux I__4702 (
            .O(N__20289),
            .I(N__20242));
    Span4Mux_h I__4701 (
            .O(N__20286),
            .I(N__20237));
    LocalMux I__4700 (
            .O(N__20283),
            .I(N__20237));
    LocalMux I__4699 (
            .O(N__20280),
            .I(N__20234));
    InMux I__4698 (
            .O(N__20279),
            .I(N__20229));
    InMux I__4697 (
            .O(N__20278),
            .I(N__20229));
    InMux I__4696 (
            .O(N__20277),
            .I(N__20216));
    InMux I__4695 (
            .O(N__20276),
            .I(N__20216));
    InMux I__4694 (
            .O(N__20275),
            .I(N__20216));
    InMux I__4693 (
            .O(N__20274),
            .I(N__20216));
    InMux I__4692 (
            .O(N__20271),
            .I(N__20216));
    InMux I__4691 (
            .O(N__20270),
            .I(N__20216));
    InMux I__4690 (
            .O(N__20267),
            .I(N__20211));
    InMux I__4689 (
            .O(N__20264),
            .I(N__20211));
    Span4Mux_v I__4688 (
            .O(N__20255),
            .I(N__20204));
    Span4Mux_v I__4687 (
            .O(N__20252),
            .I(N__20204));
    Span4Mux_h I__4686 (
            .O(N__20245),
            .I(N__20204));
    LocalMux I__4685 (
            .O(N__20242),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    Odrv4 I__4684 (
            .O(N__20237),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    Odrv4 I__4683 (
            .O(N__20234),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    LocalMux I__4682 (
            .O(N__20229),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    LocalMux I__4681 (
            .O(N__20216),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    LocalMux I__4680 (
            .O(N__20211),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    Odrv4 I__4679 (
            .O(N__20204),
            .I(\c0.byte_transmit_counter2Z0Z_2 ));
    InMux I__4678 (
            .O(N__20189),
            .I(N__20186));
    LocalMux I__4677 (
            .O(N__20186),
            .I(N__20183));
    Span4Mux_v I__4676 (
            .O(N__20183),
            .I(N__20180));
    Odrv4 I__4675 (
            .O(N__20180),
            .I(\c0.tx2_data_1_iv_5_5 ));
    InMux I__4674 (
            .O(N__20177),
            .I(N__20174));
    LocalMux I__4673 (
            .O(N__20174),
            .I(N__20171));
    Odrv4 I__4672 (
            .O(N__20171),
            .I(\c0.data_in_frame_6_Z0Z_5 ));
    InMux I__4671 (
            .O(N__20168),
            .I(N__20165));
    LocalMux I__4670 (
            .O(N__20165),
            .I(N__20162));
    Span4Mux_v I__4669 (
            .O(N__20162),
            .I(N__20153));
    InMux I__4668 (
            .O(N__20161),
            .I(N__20150));
    InMux I__4667 (
            .O(N__20160),
            .I(N__20145));
    InMux I__4666 (
            .O(N__20159),
            .I(N__20145));
    InMux I__4665 (
            .O(N__20158),
            .I(N__20142));
    InMux I__4664 (
            .O(N__20157),
            .I(N__20137));
    InMux I__4663 (
            .O(N__20156),
            .I(N__20137));
    Odrv4 I__4662 (
            .O(N__20153),
            .I(\c0.d_4_37 ));
    LocalMux I__4661 (
            .O(N__20150),
            .I(\c0.d_4_37 ));
    LocalMux I__4660 (
            .O(N__20145),
            .I(\c0.d_4_37 ));
    LocalMux I__4659 (
            .O(N__20142),
            .I(\c0.d_4_37 ));
    LocalMux I__4658 (
            .O(N__20137),
            .I(\c0.d_4_37 ));
    InMux I__4657 (
            .O(N__20126),
            .I(N__20123));
    LocalMux I__4656 (
            .O(N__20123),
            .I(\c0.tx2_data_1_iv_5_1_0_5 ));
    InMux I__4655 (
            .O(N__20120),
            .I(N__20117));
    LocalMux I__4654 (
            .O(N__20117),
            .I(N__20114));
    Span4Mux_h I__4653 (
            .O(N__20114),
            .I(N__20111));
    Odrv4 I__4652 (
            .O(N__20111),
            .I(\c0.rx.r_Rx_Bytece_1_6 ));
    InMux I__4651 (
            .O(N__20108),
            .I(N__20104));
    CascadeMux I__4650 (
            .O(N__20107),
            .I(N__20101));
    LocalMux I__4649 (
            .O(N__20104),
            .I(N__20098));
    InMux I__4648 (
            .O(N__20101),
            .I(N__20095));
    Odrv4 I__4647 (
            .O(N__20098),
            .I(\c0.rx_data_6 ));
    LocalMux I__4646 (
            .O(N__20095),
            .I(\c0.rx_data_6 ));
    CascadeMux I__4645 (
            .O(N__20090),
            .I(\c0.un1_byte_transmit_counter2_1_ac0_3_out_cascade_ ));
    CascadeMux I__4644 (
            .O(N__20087),
            .I(N__20079));
    InMux I__4643 (
            .O(N__20086),
            .I(N__20069));
    InMux I__4642 (
            .O(N__20085),
            .I(N__20069));
    InMux I__4641 (
            .O(N__20084),
            .I(N__20069));
    InMux I__4640 (
            .O(N__20083),
            .I(N__20069));
    InMux I__4639 (
            .O(N__20082),
            .I(N__20066));
    InMux I__4638 (
            .O(N__20079),
            .I(N__20061));
    InMux I__4637 (
            .O(N__20078),
            .I(N__20061));
    LocalMux I__4636 (
            .O(N__20069),
            .I(\c0.wait_for_transmission_RNI9PP5BZ0Z1 ));
    LocalMux I__4635 (
            .O(N__20066),
            .I(\c0.wait_for_transmission_RNI9PP5BZ0Z1 ));
    LocalMux I__4634 (
            .O(N__20061),
            .I(\c0.wait_for_transmission_RNI9PP5BZ0Z1 ));
    SRMux I__4633 (
            .O(N__20054),
            .I(N__20050));
    SRMux I__4632 (
            .O(N__20053),
            .I(N__20047));
    LocalMux I__4631 (
            .O(N__20050),
            .I(N__20042));
    LocalMux I__4630 (
            .O(N__20047),
            .I(N__20039));
    SRMux I__4629 (
            .O(N__20046),
            .I(N__20036));
    SRMux I__4628 (
            .O(N__20045),
            .I(N__20033));
    Span4Mux_h I__4627 (
            .O(N__20042),
            .I(N__20028));
    Span4Mux_v I__4626 (
            .O(N__20039),
            .I(N__20028));
    LocalMux I__4625 (
            .O(N__20036),
            .I(N__20025));
    LocalMux I__4624 (
            .O(N__20033),
            .I(N__20022));
    Sp12to4 I__4623 (
            .O(N__20028),
            .I(N__20019));
    Span12Mux_v I__4622 (
            .O(N__20025),
            .I(N__20016));
    Odrv4 I__4621 (
            .O(N__20022),
            .I(\c0.tx2_transmit_0_sqmuxa ));
    Odrv12 I__4620 (
            .O(N__20019),
            .I(\c0.tx2_transmit_0_sqmuxa ));
    Odrv12 I__4619 (
            .O(N__20016),
            .I(\c0.tx2_transmit_0_sqmuxa ));
    InMux I__4618 (
            .O(N__20009),
            .I(N__20006));
    LocalMux I__4617 (
            .O(N__20006),
            .I(N__20003));
    Span4Mux_v I__4616 (
            .O(N__20003),
            .I(N__19999));
    InMux I__4615 (
            .O(N__20002),
            .I(N__19996));
    Span4Mux_h I__4614 (
            .O(N__19999),
            .I(N__19993));
    LocalMux I__4613 (
            .O(N__19996),
            .I(N__19990));
    Odrv4 I__4612 (
            .O(N__19993),
            .I(\c0.data_in_4_Z0Z_5 ));
    Odrv4 I__4611 (
            .O(N__19990),
            .I(\c0.data_in_4_Z0Z_5 ));
    InMux I__4610 (
            .O(N__19985),
            .I(N__19982));
    LocalMux I__4609 (
            .O(N__19982),
            .I(N__19979));
    Span12Mux_h I__4608 (
            .O(N__19979),
            .I(N__19975));
    InMux I__4607 (
            .O(N__19978),
            .I(N__19972));
    Odrv12 I__4606 (
            .O(N__19975),
            .I(\c0.data_in_5_Z0Z_5 ));
    LocalMux I__4605 (
            .O(N__19972),
            .I(\c0.data_in_5_Z0Z_5 ));
    InMux I__4604 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__4603 (
            .O(N__19964),
            .I(N__19958));
    InMux I__4602 (
            .O(N__19963),
            .I(N__19955));
    CascadeMux I__4601 (
            .O(N__19962),
            .I(N__19951));
    CascadeMux I__4600 (
            .O(N__19961),
            .I(N__19948));
    Span4Mux_h I__4599 (
            .O(N__19958),
            .I(N__19945));
    LocalMux I__4598 (
            .O(N__19955),
            .I(N__19942));
    InMux I__4597 (
            .O(N__19954),
            .I(N__19935));
    InMux I__4596 (
            .O(N__19951),
            .I(N__19935));
    InMux I__4595 (
            .O(N__19948),
            .I(N__19935));
    Odrv4 I__4594 (
            .O(N__19945),
            .I(\c0.data_in_7_Z0Z_5 ));
    Odrv12 I__4593 (
            .O(N__19942),
            .I(\c0.data_in_7_Z0Z_5 ));
    LocalMux I__4592 (
            .O(N__19935),
            .I(\c0.data_in_7_Z0Z_5 ));
    CascadeMux I__4591 (
            .O(N__19928),
            .I(N__19924));
    InMux I__4590 (
            .O(N__19927),
            .I(N__19921));
    InMux I__4589 (
            .O(N__19924),
            .I(N__19918));
    LocalMux I__4588 (
            .O(N__19921),
            .I(N__19915));
    LocalMux I__4587 (
            .O(N__19918),
            .I(N__19911));
    Span4Mux_v I__4586 (
            .O(N__19915),
            .I(N__19908));
    InMux I__4585 (
            .O(N__19914),
            .I(N__19905));
    Span4Mux_h I__4584 (
            .O(N__19911),
            .I(N__19902));
    Odrv4 I__4583 (
            .O(N__19908),
            .I(\c0.data_in_6_Z0Z_5 ));
    LocalMux I__4582 (
            .O(N__19905),
            .I(\c0.data_in_6_Z0Z_5 ));
    Odrv4 I__4581 (
            .O(N__19902),
            .I(\c0.data_in_6_Z0Z_5 ));
    InMux I__4580 (
            .O(N__19895),
            .I(N__19892));
    LocalMux I__4579 (
            .O(N__19892),
            .I(N__19889));
    Span4Mux_v I__4578 (
            .O(N__19889),
            .I(N__19885));
    InMux I__4577 (
            .O(N__19888),
            .I(N__19882));
    Odrv4 I__4576 (
            .O(N__19885),
            .I(\c0.data_in_5_Z0Z_6 ));
    LocalMux I__4575 (
            .O(N__19882),
            .I(\c0.data_in_5_Z0Z_6 ));
    CascadeMux I__4574 (
            .O(N__19877),
            .I(N__19874));
    InMux I__4573 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__4572 (
            .O(N__19871),
            .I(N__19866));
    InMux I__4571 (
            .O(N__19870),
            .I(N__19863));
    InMux I__4570 (
            .O(N__19869),
            .I(N__19860));
    Span4Mux_h I__4569 (
            .O(N__19866),
            .I(N__19857));
    LocalMux I__4568 (
            .O(N__19863),
            .I(\c0.data_in_7_Z0Z_6 ));
    LocalMux I__4567 (
            .O(N__19860),
            .I(\c0.data_in_7_Z0Z_6 ));
    Odrv4 I__4566 (
            .O(N__19857),
            .I(\c0.data_in_7_Z0Z_6 ));
    InMux I__4565 (
            .O(N__19850),
            .I(N__19846));
    InMux I__4564 (
            .O(N__19849),
            .I(N__19843));
    LocalMux I__4563 (
            .O(N__19846),
            .I(N__19840));
    LocalMux I__4562 (
            .O(N__19843),
            .I(N__19837));
    Span12Mux_v I__4561 (
            .O(N__19840),
            .I(N__19834));
    Span4Mux_v I__4560 (
            .O(N__19837),
            .I(N__19831));
    Odrv12 I__4559 (
            .O(N__19834),
            .I(\c0.d_4_RNII9QU3Z0Z_14 ));
    Odrv4 I__4558 (
            .O(N__19831),
            .I(\c0.d_4_RNII9QU3Z0Z_14 ));
    InMux I__4557 (
            .O(N__19826),
            .I(N__19822));
    InMux I__4556 (
            .O(N__19825),
            .I(N__19819));
    LocalMux I__4555 (
            .O(N__19822),
            .I(N__19814));
    LocalMux I__4554 (
            .O(N__19819),
            .I(N__19814));
    Odrv12 I__4553 (
            .O(N__19814),
            .I(\c0.wait_for_transmission_RNI94LSZ0Z6 ));
    CascadeMux I__4552 (
            .O(N__19811),
            .I(N__19808));
    InMux I__4551 (
            .O(N__19808),
            .I(N__19804));
    InMux I__4550 (
            .O(N__19807),
            .I(N__19800));
    LocalMux I__4549 (
            .O(N__19804),
            .I(N__19797));
    InMux I__4548 (
            .O(N__19803),
            .I(N__19794));
    LocalMux I__4547 (
            .O(N__19800),
            .I(N__19789));
    Sp12to4 I__4546 (
            .O(N__19797),
            .I(N__19784));
    LocalMux I__4545 (
            .O(N__19794),
            .I(N__19784));
    InMux I__4544 (
            .O(N__19793),
            .I(N__19781));
    InMux I__4543 (
            .O(N__19792),
            .I(N__19778));
    Odrv4 I__4542 (
            .O(N__19789),
            .I(\c0.wait_for_transmissionZ0 ));
    Odrv12 I__4541 (
            .O(N__19784),
            .I(\c0.wait_for_transmissionZ0 ));
    LocalMux I__4540 (
            .O(N__19781),
            .I(\c0.wait_for_transmissionZ0 ));
    LocalMux I__4539 (
            .O(N__19778),
            .I(\c0.wait_for_transmissionZ0 ));
    InMux I__4538 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__4537 (
            .O(N__19766),
            .I(\c0.d_4_RNI9LFUVZ0Z_43 ));
    InMux I__4536 (
            .O(N__19763),
            .I(N__19760));
    LocalMux I__4535 (
            .O(N__19760),
            .I(N__19755));
    InMux I__4534 (
            .O(N__19759),
            .I(N__19750));
    InMux I__4533 (
            .O(N__19758),
            .I(N__19750));
    Span12Mux_h I__4532 (
            .O(N__19755),
            .I(N__19747));
    LocalMux I__4531 (
            .O(N__19750),
            .I(N__19744));
    Odrv12 I__4530 (
            .O(N__19747),
            .I(\c0.tx2_transmitZ0 ));
    Odrv12 I__4529 (
            .O(N__19744),
            .I(\c0.tx2_transmitZ0 ));
    InMux I__4528 (
            .O(N__19739),
            .I(N__19735));
    InMux I__4527 (
            .O(N__19738),
            .I(N__19732));
    LocalMux I__4526 (
            .O(N__19735),
            .I(\c0.m2_e_0_2 ));
    LocalMux I__4525 (
            .O(N__19732),
            .I(\c0.m2_e_0_2 ));
    InMux I__4524 (
            .O(N__19727),
            .I(N__19723));
    InMux I__4523 (
            .O(N__19726),
            .I(N__19720));
    LocalMux I__4522 (
            .O(N__19723),
            .I(N__19717));
    LocalMux I__4521 (
            .O(N__19720),
            .I(N__19714));
    Span4Mux_v I__4520 (
            .O(N__19717),
            .I(N__19707));
    Span4Mux_v I__4519 (
            .O(N__19714),
            .I(N__19707));
    InMux I__4518 (
            .O(N__19713),
            .I(N__19702));
    InMux I__4517 (
            .O(N__19712),
            .I(N__19702));
    Odrv4 I__4516 (
            .O(N__19707),
            .I(\c0.d_4_20 ));
    LocalMux I__4515 (
            .O(N__19702),
            .I(\c0.d_4_20 ));
    CascadeMux I__4514 (
            .O(N__19697),
            .I(\c0.N_203_cascade_ ));
    InMux I__4513 (
            .O(N__19694),
            .I(N__19691));
    LocalMux I__4512 (
            .O(N__19691),
            .I(N__19688));
    Span4Mux_h I__4511 (
            .O(N__19688),
            .I(N__19684));
    InMux I__4510 (
            .O(N__19687),
            .I(N__19681));
    Odrv4 I__4509 (
            .O(N__19684),
            .I(\c0.d_4_4 ));
    LocalMux I__4508 (
            .O(N__19681),
            .I(\c0.d_4_4 ));
    InMux I__4507 (
            .O(N__19676),
            .I(N__19673));
    LocalMux I__4506 (
            .O(N__19673),
            .I(\c0.tx2_data_1_iv_5_1_4 ));
    CascadeMux I__4505 (
            .O(N__19670),
            .I(\c0.un1_m4_0_a2_2_cascade_ ));
    InMux I__4504 (
            .O(N__19667),
            .I(N__19663));
    InMux I__4503 (
            .O(N__19666),
            .I(N__19660));
    LocalMux I__4502 (
            .O(N__19663),
            .I(\c0.byte_transmit_counter2Z0Z_7 ));
    LocalMux I__4501 (
            .O(N__19660),
            .I(\c0.byte_transmit_counter2Z0Z_7 ));
    InMux I__4500 (
            .O(N__19655),
            .I(N__19652));
    LocalMux I__4499 (
            .O(N__19652),
            .I(\c0.un1_m4_0_a2_1_0 ));
    CascadeMux I__4498 (
            .O(N__19649),
            .I(N__19644));
    CascadeMux I__4497 (
            .O(N__19648),
            .I(N__19641));
    CascadeMux I__4496 (
            .O(N__19647),
            .I(N__19638));
    InMux I__4495 (
            .O(N__19644),
            .I(N__19634));
    InMux I__4494 (
            .O(N__19641),
            .I(N__19631));
    InMux I__4493 (
            .O(N__19638),
            .I(N__19625));
    InMux I__4492 (
            .O(N__19637),
            .I(N__19625));
    LocalMux I__4491 (
            .O(N__19634),
            .I(N__19622));
    LocalMux I__4490 (
            .O(N__19631),
            .I(N__19619));
    InMux I__4489 (
            .O(N__19630),
            .I(N__19616));
    LocalMux I__4488 (
            .O(N__19625),
            .I(\c0.byte_transmit_counter2Z0Z_6 ));
    Odrv4 I__4487 (
            .O(N__19622),
            .I(\c0.byte_transmit_counter2Z0Z_6 ));
    Odrv4 I__4486 (
            .O(N__19619),
            .I(\c0.byte_transmit_counter2Z0Z_6 ));
    LocalMux I__4485 (
            .O(N__19616),
            .I(\c0.byte_transmit_counter2Z0Z_6 ));
    InMux I__4484 (
            .O(N__19607),
            .I(N__19601));
    InMux I__4483 (
            .O(N__19606),
            .I(N__19596));
    InMux I__4482 (
            .O(N__19605),
            .I(N__19591));
    InMux I__4481 (
            .O(N__19604),
            .I(N__19591));
    LocalMux I__4480 (
            .O(N__19601),
            .I(N__19588));
    InMux I__4479 (
            .O(N__19600),
            .I(N__19583));
    InMux I__4478 (
            .O(N__19599),
            .I(N__19583));
    LocalMux I__4477 (
            .O(N__19596),
            .I(\c0.byte_transmit_counter2Z0Z_5 ));
    LocalMux I__4476 (
            .O(N__19591),
            .I(\c0.byte_transmit_counter2Z0Z_5 ));
    Odrv4 I__4475 (
            .O(N__19588),
            .I(\c0.byte_transmit_counter2Z0Z_5 ));
    LocalMux I__4474 (
            .O(N__19583),
            .I(\c0.byte_transmit_counter2Z0Z_5 ));
    CascadeMux I__4473 (
            .O(N__19574),
            .I(N__19569));
    CascadeMux I__4472 (
            .O(N__19573),
            .I(N__19565));
    InMux I__4471 (
            .O(N__19572),
            .I(N__19560));
    InMux I__4470 (
            .O(N__19569),
            .I(N__19553));
    InMux I__4469 (
            .O(N__19568),
            .I(N__19553));
    InMux I__4468 (
            .O(N__19565),
            .I(N__19553));
    CascadeMux I__4467 (
            .O(N__19564),
            .I(N__19550));
    CascadeMux I__4466 (
            .O(N__19563),
            .I(N__19547));
    LocalMux I__4465 (
            .O(N__19560),
            .I(N__19542));
    LocalMux I__4464 (
            .O(N__19553),
            .I(N__19542));
    InMux I__4463 (
            .O(N__19550),
            .I(N__19536));
    InMux I__4462 (
            .O(N__19547),
            .I(N__19533));
    Span4Mux_h I__4461 (
            .O(N__19542),
            .I(N__19530));
    InMux I__4460 (
            .O(N__19541),
            .I(N__19527));
    CascadeMux I__4459 (
            .O(N__19540),
            .I(N__19524));
    CascadeMux I__4458 (
            .O(N__19539),
            .I(N__19520));
    LocalMux I__4457 (
            .O(N__19536),
            .I(N__19515));
    LocalMux I__4456 (
            .O(N__19533),
            .I(N__19515));
    Span4Mux_h I__4455 (
            .O(N__19530),
            .I(N__19510));
    LocalMux I__4454 (
            .O(N__19527),
            .I(N__19510));
    InMux I__4453 (
            .O(N__19524),
            .I(N__19503));
    InMux I__4452 (
            .O(N__19523),
            .I(N__19503));
    InMux I__4451 (
            .O(N__19520),
            .I(N__19503));
    Span4Mux_v I__4450 (
            .O(N__19515),
            .I(N__19497));
    Span4Mux_v I__4449 (
            .O(N__19510),
            .I(N__19497));
    LocalMux I__4448 (
            .O(N__19503),
            .I(N__19494));
    CascadeMux I__4447 (
            .O(N__19502),
            .I(N__19489));
    Span4Mux_h I__4446 (
            .O(N__19497),
            .I(N__19475));
    Span4Mux_v I__4445 (
            .O(N__19494),
            .I(N__19475));
    InMux I__4444 (
            .O(N__19493),
            .I(N__19466));
    InMux I__4443 (
            .O(N__19492),
            .I(N__19466));
    InMux I__4442 (
            .O(N__19489),
            .I(N__19466));
    InMux I__4441 (
            .O(N__19488),
            .I(N__19466));
    InMux I__4440 (
            .O(N__19487),
            .I(N__19459));
    InMux I__4439 (
            .O(N__19486),
            .I(N__19459));
    InMux I__4438 (
            .O(N__19485),
            .I(N__19459));
    InMux I__4437 (
            .O(N__19484),
            .I(N__19454));
    InMux I__4436 (
            .O(N__19483),
            .I(N__19454));
    InMux I__4435 (
            .O(N__19482),
            .I(N__19449));
    InMux I__4434 (
            .O(N__19481),
            .I(N__19449));
    InMux I__4433 (
            .O(N__19480),
            .I(N__19446));
    Sp12to4 I__4432 (
            .O(N__19475),
            .I(N__19441));
    LocalMux I__4431 (
            .O(N__19466),
            .I(N__19441));
    LocalMux I__4430 (
            .O(N__19459),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4429 (
            .O(N__19454),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4428 (
            .O(N__19449),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    LocalMux I__4427 (
            .O(N__19446),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    Odrv12 I__4426 (
            .O(N__19441),
            .I(\c0.byte_transmit_counter2Z0Z_0 ));
    InMux I__4425 (
            .O(N__19430),
            .I(N__19427));
    LocalMux I__4424 (
            .O(N__19427),
            .I(N__19424));
    Span4Mux_h I__4423 (
            .O(N__19424),
            .I(N__19420));
    InMux I__4422 (
            .O(N__19423),
            .I(N__19417));
    Odrv4 I__4421 (
            .O(N__19420),
            .I(\c0.N_201 ));
    LocalMux I__4420 (
            .O(N__19417),
            .I(\c0.N_201 ));
    InMux I__4419 (
            .O(N__19412),
            .I(N__19407));
    InMux I__4418 (
            .O(N__19411),
            .I(N__19404));
    InMux I__4417 (
            .O(N__19410),
            .I(N__19393));
    LocalMux I__4416 (
            .O(N__19407),
            .I(N__19388));
    LocalMux I__4415 (
            .O(N__19404),
            .I(N__19388));
    InMux I__4414 (
            .O(N__19403),
            .I(N__19381));
    InMux I__4413 (
            .O(N__19402),
            .I(N__19381));
    InMux I__4412 (
            .O(N__19401),
            .I(N__19381));
    InMux I__4411 (
            .O(N__19400),
            .I(N__19376));
    InMux I__4410 (
            .O(N__19399),
            .I(N__19376));
    InMux I__4409 (
            .O(N__19398),
            .I(N__19367));
    InMux I__4408 (
            .O(N__19397),
            .I(N__19364));
    InMux I__4407 (
            .O(N__19396),
            .I(N__19358));
    LocalMux I__4406 (
            .O(N__19393),
            .I(N__19351));
    Span4Mux_v I__4405 (
            .O(N__19388),
            .I(N__19351));
    LocalMux I__4404 (
            .O(N__19381),
            .I(N__19351));
    LocalMux I__4403 (
            .O(N__19376),
            .I(N__19348));
    InMux I__4402 (
            .O(N__19375),
            .I(N__19337));
    InMux I__4401 (
            .O(N__19374),
            .I(N__19337));
    InMux I__4400 (
            .O(N__19373),
            .I(N__19337));
    InMux I__4399 (
            .O(N__19372),
            .I(N__19337));
    InMux I__4398 (
            .O(N__19371),
            .I(N__19337));
    InMux I__4397 (
            .O(N__19370),
            .I(N__19334));
    LocalMux I__4396 (
            .O(N__19367),
            .I(N__19331));
    LocalMux I__4395 (
            .O(N__19364),
            .I(N__19328));
    InMux I__4394 (
            .O(N__19363),
            .I(N__19323));
    InMux I__4393 (
            .O(N__19362),
            .I(N__19323));
    InMux I__4392 (
            .O(N__19361),
            .I(N__19315));
    LocalMux I__4391 (
            .O(N__19358),
            .I(N__19302));
    Span4Mux_h I__4390 (
            .O(N__19351),
            .I(N__19302));
    Span4Mux_v I__4389 (
            .O(N__19348),
            .I(N__19302));
    LocalMux I__4388 (
            .O(N__19337),
            .I(N__19302));
    LocalMux I__4387 (
            .O(N__19334),
            .I(N__19293));
    Span4Mux_v I__4386 (
            .O(N__19331),
            .I(N__19293));
    Span4Mux_v I__4385 (
            .O(N__19328),
            .I(N__19293));
    LocalMux I__4384 (
            .O(N__19323),
            .I(N__19293));
    InMux I__4383 (
            .O(N__19322),
            .I(N__19288));
    InMux I__4382 (
            .O(N__19321),
            .I(N__19288));
    InMux I__4381 (
            .O(N__19320),
            .I(N__19283));
    InMux I__4380 (
            .O(N__19319),
            .I(N__19278));
    InMux I__4379 (
            .O(N__19318),
            .I(N__19278));
    LocalMux I__4378 (
            .O(N__19315),
            .I(N__19275));
    InMux I__4377 (
            .O(N__19314),
            .I(N__19266));
    InMux I__4376 (
            .O(N__19313),
            .I(N__19266));
    InMux I__4375 (
            .O(N__19312),
            .I(N__19266));
    InMux I__4374 (
            .O(N__19311),
            .I(N__19266));
    Span4Mux_h I__4373 (
            .O(N__19302),
            .I(N__19263));
    Span4Mux_h I__4372 (
            .O(N__19293),
            .I(N__19258));
    LocalMux I__4371 (
            .O(N__19288),
            .I(N__19258));
    InMux I__4370 (
            .O(N__19287),
            .I(N__19253));
    InMux I__4369 (
            .O(N__19286),
            .I(N__19253));
    LocalMux I__4368 (
            .O(N__19283),
            .I(\c0.N_129_mux ));
    LocalMux I__4367 (
            .O(N__19278),
            .I(\c0.N_129_mux ));
    Odrv12 I__4366 (
            .O(N__19275),
            .I(\c0.N_129_mux ));
    LocalMux I__4365 (
            .O(N__19266),
            .I(\c0.N_129_mux ));
    Odrv4 I__4364 (
            .O(N__19263),
            .I(\c0.N_129_mux ));
    Odrv4 I__4363 (
            .O(N__19258),
            .I(\c0.N_129_mux ));
    LocalMux I__4362 (
            .O(N__19253),
            .I(\c0.N_129_mux ));
    InMux I__4361 (
            .O(N__19238),
            .I(N__19229));
    CascadeMux I__4360 (
            .O(N__19237),
            .I(N__19226));
    CascadeMux I__4359 (
            .O(N__19236),
            .I(N__19223));
    CascadeMux I__4358 (
            .O(N__19235),
            .I(N__19219));
    CascadeMux I__4357 (
            .O(N__19234),
            .I(N__19215));
    CascadeMux I__4356 (
            .O(N__19233),
            .I(N__19210));
    CascadeMux I__4355 (
            .O(N__19232),
            .I(N__19206));
    LocalMux I__4354 (
            .O(N__19229),
            .I(N__19197));
    InMux I__4353 (
            .O(N__19226),
            .I(N__19186));
    InMux I__4352 (
            .O(N__19223),
            .I(N__19186));
    InMux I__4351 (
            .O(N__19222),
            .I(N__19186));
    InMux I__4350 (
            .O(N__19219),
            .I(N__19186));
    InMux I__4349 (
            .O(N__19218),
            .I(N__19186));
    InMux I__4348 (
            .O(N__19215),
            .I(N__19182));
    InMux I__4347 (
            .O(N__19214),
            .I(N__19179));
    InMux I__4346 (
            .O(N__19213),
            .I(N__19174));
    InMux I__4345 (
            .O(N__19210),
            .I(N__19174));
    InMux I__4344 (
            .O(N__19209),
            .I(N__19163));
    InMux I__4343 (
            .O(N__19206),
            .I(N__19163));
    InMux I__4342 (
            .O(N__19205),
            .I(N__19159));
    InMux I__4341 (
            .O(N__19204),
            .I(N__19153));
    InMux I__4340 (
            .O(N__19203),
            .I(N__19153));
    InMux I__4339 (
            .O(N__19202),
            .I(N__19146));
    InMux I__4338 (
            .O(N__19201),
            .I(N__19146));
    InMux I__4337 (
            .O(N__19200),
            .I(N__19146));
    Span4Mux_h I__4336 (
            .O(N__19197),
            .I(N__19143));
    LocalMux I__4335 (
            .O(N__19186),
            .I(N__19140));
    InMux I__4334 (
            .O(N__19185),
            .I(N__19137));
    LocalMux I__4333 (
            .O(N__19182),
            .I(N__19134));
    LocalMux I__4332 (
            .O(N__19179),
            .I(N__19129));
    LocalMux I__4331 (
            .O(N__19174),
            .I(N__19129));
    InMux I__4330 (
            .O(N__19173),
            .I(N__19120));
    InMux I__4329 (
            .O(N__19172),
            .I(N__19120));
    InMux I__4328 (
            .O(N__19171),
            .I(N__19120));
    InMux I__4327 (
            .O(N__19170),
            .I(N__19120));
    InMux I__4326 (
            .O(N__19169),
            .I(N__19115));
    InMux I__4325 (
            .O(N__19168),
            .I(N__19115));
    LocalMux I__4324 (
            .O(N__19163),
            .I(N__19110));
    InMux I__4323 (
            .O(N__19162),
            .I(N__19107));
    LocalMux I__4322 (
            .O(N__19159),
            .I(N__19104));
    InMux I__4321 (
            .O(N__19158),
            .I(N__19101));
    LocalMux I__4320 (
            .O(N__19153),
            .I(N__19096));
    LocalMux I__4319 (
            .O(N__19146),
            .I(N__19096));
    Span4Mux_h I__4318 (
            .O(N__19143),
            .I(N__19081));
    Span4Mux_v I__4317 (
            .O(N__19140),
            .I(N__19081));
    LocalMux I__4316 (
            .O(N__19137),
            .I(N__19081));
    Span4Mux_v I__4315 (
            .O(N__19134),
            .I(N__19081));
    Span4Mux_v I__4314 (
            .O(N__19129),
            .I(N__19081));
    LocalMux I__4313 (
            .O(N__19120),
            .I(N__19081));
    LocalMux I__4312 (
            .O(N__19115),
            .I(N__19081));
    CascadeMux I__4311 (
            .O(N__19114),
            .I(N__19078));
    InMux I__4310 (
            .O(N__19113),
            .I(N__19073));
    Span12Mux_h I__4309 (
            .O(N__19110),
            .I(N__19070));
    LocalMux I__4308 (
            .O(N__19107),
            .I(N__19061));
    Span12Mux_s8_h I__4307 (
            .O(N__19104),
            .I(N__19061));
    LocalMux I__4306 (
            .O(N__19101),
            .I(N__19061));
    Span12Mux_s9_v I__4305 (
            .O(N__19096),
            .I(N__19061));
    Span4Mux_h I__4304 (
            .O(N__19081),
            .I(N__19058));
    InMux I__4303 (
            .O(N__19078),
            .I(N__19051));
    InMux I__4302 (
            .O(N__19077),
            .I(N__19051));
    InMux I__4301 (
            .O(N__19076),
            .I(N__19051));
    LocalMux I__4300 (
            .O(N__19073),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    Odrv12 I__4299 (
            .O(N__19070),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    Odrv12 I__4298 (
            .O(N__19061),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    Odrv4 I__4297 (
            .O(N__19058),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    LocalMux I__4296 (
            .O(N__19051),
            .I(\c0.byte_transmit_counterZ0Z_2 ));
    InMux I__4295 (
            .O(N__19040),
            .I(N__19037));
    LocalMux I__4294 (
            .O(N__19037),
            .I(\c0.byte_transmit_counterZ0Z_7 ));
    CEMux I__4293 (
            .O(N__19034),
            .I(N__19031));
    LocalMux I__4292 (
            .O(N__19031),
            .I(N__19026));
    CEMux I__4291 (
            .O(N__19030),
            .I(N__19023));
    CEMux I__4290 (
            .O(N__19029),
            .I(N__19020));
    Span4Mux_h I__4289 (
            .O(N__19026),
            .I(N__19016));
    LocalMux I__4288 (
            .O(N__19023),
            .I(N__19013));
    LocalMux I__4287 (
            .O(N__19020),
            .I(N__19010));
    InMux I__4286 (
            .O(N__19019),
            .I(N__19007));
    Odrv4 I__4285 (
            .O(N__19016),
            .I(\c0.byte_transmit_counter15 ));
    Odrv4 I__4284 (
            .O(N__19013),
            .I(\c0.byte_transmit_counter15 ));
    Odrv12 I__4283 (
            .O(N__19010),
            .I(\c0.byte_transmit_counter15 ));
    LocalMux I__4282 (
            .O(N__19007),
            .I(\c0.byte_transmit_counter15 ));
    CascadeMux I__4281 (
            .O(N__18998),
            .I(N__18995));
    InMux I__4280 (
            .O(N__18995),
            .I(N__18992));
    LocalMux I__4279 (
            .O(N__18992),
            .I(N__18989));
    Odrv4 I__4278 (
            .O(N__18989),
            .I(\c0.tx2_data_1_iv_5_1_0_4 ));
    InMux I__4277 (
            .O(N__18986),
            .I(N__18982));
    InMux I__4276 (
            .O(N__18985),
            .I(N__18979));
    LocalMux I__4275 (
            .O(N__18982),
            .I(N__18976));
    LocalMux I__4274 (
            .O(N__18979),
            .I(\c0.N_207 ));
    Odrv4 I__4273 (
            .O(N__18976),
            .I(\c0.N_207 ));
    CascadeMux I__4272 (
            .O(N__18971),
            .I(\c0.N_207_cascade_ ));
    InMux I__4271 (
            .O(N__18968),
            .I(N__18964));
    InMux I__4270 (
            .O(N__18967),
            .I(N__18961));
    LocalMux I__4269 (
            .O(N__18964),
            .I(N__18958));
    LocalMux I__4268 (
            .O(N__18961),
            .I(N__18953));
    Span12Mux_h I__4267 (
            .O(N__18958),
            .I(N__18950));
    InMux I__4266 (
            .O(N__18957),
            .I(N__18947));
    InMux I__4265 (
            .O(N__18956),
            .I(N__18944));
    Span4Mux_h I__4264 (
            .O(N__18953),
            .I(N__18941));
    Odrv12 I__4263 (
            .O(N__18950),
            .I(\c0.d_4_28 ));
    LocalMux I__4262 (
            .O(N__18947),
            .I(\c0.d_4_28 ));
    LocalMux I__4261 (
            .O(N__18944),
            .I(\c0.d_4_28 ));
    Odrv4 I__4260 (
            .O(N__18941),
            .I(\c0.d_4_28 ));
    CascadeMux I__4259 (
            .O(N__18932),
            .I(\c0.m2_e_0_2_cascade_ ));
    InMux I__4258 (
            .O(N__18929),
            .I(N__18912));
    InMux I__4257 (
            .O(N__18928),
            .I(N__18912));
    InMux I__4256 (
            .O(N__18927),
            .I(N__18912));
    InMux I__4255 (
            .O(N__18926),
            .I(N__18912));
    InMux I__4254 (
            .O(N__18925),
            .I(N__18907));
    InMux I__4253 (
            .O(N__18924),
            .I(N__18898));
    InMux I__4252 (
            .O(N__18923),
            .I(N__18898));
    InMux I__4251 (
            .O(N__18922),
            .I(N__18898));
    InMux I__4250 (
            .O(N__18921),
            .I(N__18898));
    LocalMux I__4249 (
            .O(N__18912),
            .I(N__18892));
    InMux I__4248 (
            .O(N__18911),
            .I(N__18889));
    InMux I__4247 (
            .O(N__18910),
            .I(N__18886));
    LocalMux I__4246 (
            .O(N__18907),
            .I(N__18881));
    LocalMux I__4245 (
            .O(N__18898),
            .I(N__18881));
    InMux I__4244 (
            .O(N__18897),
            .I(N__18874));
    InMux I__4243 (
            .O(N__18896),
            .I(N__18874));
    InMux I__4242 (
            .O(N__18895),
            .I(N__18874));
    Span4Mux_h I__4241 (
            .O(N__18892),
            .I(N__18868));
    LocalMux I__4240 (
            .O(N__18889),
            .I(N__18868));
    LocalMux I__4239 (
            .O(N__18886),
            .I(N__18861));
    Span4Mux_v I__4238 (
            .O(N__18881),
            .I(N__18861));
    LocalMux I__4237 (
            .O(N__18874),
            .I(N__18861));
    InMux I__4236 (
            .O(N__18873),
            .I(N__18858));
    Span4Mux_v I__4235 (
            .O(N__18868),
            .I(N__18853));
    Span4Mux_h I__4234 (
            .O(N__18861),
            .I(N__18853));
    LocalMux I__4233 (
            .O(N__18858),
            .I(\c0.N_71_mux ));
    Odrv4 I__4232 (
            .O(N__18853),
            .I(\c0.N_71_mux ));
    InMux I__4231 (
            .O(N__18848),
            .I(N__18845));
    LocalMux I__4230 (
            .O(N__18845),
            .I(N__18842));
    Span4Mux_v I__4229 (
            .O(N__18842),
            .I(N__18838));
    InMux I__4228 (
            .O(N__18841),
            .I(N__18835));
    Span4Mux_h I__4227 (
            .O(N__18838),
            .I(N__18830));
    LocalMux I__4226 (
            .O(N__18835),
            .I(N__18830));
    Odrv4 I__4225 (
            .O(N__18830),
            .I(\c0.data_in_4_Z0Z_7 ));
    InMux I__4224 (
            .O(N__18827),
            .I(N__18823));
    CascadeMux I__4223 (
            .O(N__18826),
            .I(N__18820));
    LocalMux I__4222 (
            .O(N__18823),
            .I(N__18817));
    InMux I__4221 (
            .O(N__18820),
            .I(N__18814));
    Odrv12 I__4220 (
            .O(N__18817),
            .I(\c0.rx_data_7 ));
    LocalMux I__4219 (
            .O(N__18814),
            .I(\c0.rx_data_7 ));
    InMux I__4218 (
            .O(N__18809),
            .I(N__18806));
    LocalMux I__4217 (
            .O(N__18806),
            .I(N__18802));
    InMux I__4216 (
            .O(N__18805),
            .I(N__18798));
    Span4Mux_h I__4215 (
            .O(N__18802),
            .I(N__18795));
    InMux I__4214 (
            .O(N__18801),
            .I(N__18792));
    LocalMux I__4213 (
            .O(N__18798),
            .I(N__18789));
    Odrv4 I__4212 (
            .O(N__18795),
            .I(\c0.data_in_6_Z0Z_1 ));
    LocalMux I__4211 (
            .O(N__18792),
            .I(\c0.data_in_6_Z0Z_1 ));
    Odrv4 I__4210 (
            .O(N__18789),
            .I(\c0.data_in_6_Z0Z_1 ));
    InMux I__4209 (
            .O(N__18782),
            .I(N__18778));
    CascadeMux I__4208 (
            .O(N__18781),
            .I(N__18775));
    LocalMux I__4207 (
            .O(N__18778),
            .I(N__18772));
    InMux I__4206 (
            .O(N__18775),
            .I(N__18769));
    Span4Mux_h I__4205 (
            .O(N__18772),
            .I(N__18766));
    LocalMux I__4204 (
            .O(N__18769),
            .I(N__18762));
    Span4Mux_h I__4203 (
            .O(N__18766),
            .I(N__18759));
    InMux I__4202 (
            .O(N__18765),
            .I(N__18756));
    Span4Mux_h I__4201 (
            .O(N__18762),
            .I(N__18753));
    Odrv4 I__4200 (
            .O(N__18759),
            .I(\c0.data_in_6_Z0Z_0 ));
    LocalMux I__4199 (
            .O(N__18756),
            .I(\c0.data_in_6_Z0Z_0 ));
    Odrv4 I__4198 (
            .O(N__18753),
            .I(\c0.data_in_6_Z0Z_0 ));
    CascadeMux I__4197 (
            .O(N__18746),
            .I(N__18743));
    InMux I__4196 (
            .O(N__18743),
            .I(N__18739));
    InMux I__4195 (
            .O(N__18742),
            .I(N__18735));
    LocalMux I__4194 (
            .O(N__18739),
            .I(N__18732));
    InMux I__4193 (
            .O(N__18738),
            .I(N__18729));
    LocalMux I__4192 (
            .O(N__18735),
            .I(N__18724));
    Span4Mux_v I__4191 (
            .O(N__18732),
            .I(N__18724));
    LocalMux I__4190 (
            .O(N__18729),
            .I(\c0.data_in_7_Z0Z_0 ));
    Odrv4 I__4189 (
            .O(N__18724),
            .I(\c0.data_in_7_Z0Z_0 ));
    InMux I__4188 (
            .O(N__18719),
            .I(N__18715));
    InMux I__4187 (
            .O(N__18718),
            .I(N__18712));
    LocalMux I__4186 (
            .O(N__18715),
            .I(N__18709));
    LocalMux I__4185 (
            .O(N__18712),
            .I(N__18706));
    Span12Mux_h I__4184 (
            .O(N__18709),
            .I(N__18703));
    Span4Mux_h I__4183 (
            .O(N__18706),
            .I(N__18700));
    Odrv12 I__4182 (
            .O(N__18703),
            .I(\c0.data_in_5_Z0Z_4 ));
    Odrv4 I__4181 (
            .O(N__18700),
            .I(\c0.data_in_5_Z0Z_4 ));
    InMux I__4180 (
            .O(N__18695),
            .I(N__18692));
    LocalMux I__4179 (
            .O(N__18692),
            .I(\c0.byte_transmit_counterZ0Z_5 ));
    InMux I__4178 (
            .O(N__18689),
            .I(N__18686));
    LocalMux I__4177 (
            .O(N__18686),
            .I(\c0.d_4_RNIU6U8Z0Z_22 ));
    CascadeMux I__4176 (
            .O(N__18683),
            .I(\c0.d_4_RNIU6U8_0Z0Z_22_cascade_ ));
    InMux I__4175 (
            .O(N__18680),
            .I(N__18677));
    LocalMux I__4174 (
            .O(N__18677),
            .I(\c0.d_4_RNIMI4KZ0Z_37 ));
    InMux I__4173 (
            .O(N__18674),
            .I(N__18670));
    InMux I__4172 (
            .O(N__18673),
            .I(N__18667));
    LocalMux I__4171 (
            .O(N__18670),
            .I(N__18663));
    LocalMux I__4170 (
            .O(N__18667),
            .I(N__18660));
    InMux I__4169 (
            .O(N__18666),
            .I(N__18657));
    Odrv4 I__4168 (
            .O(N__18663),
            .I(\c0.data_in_3_Z0Z_0 ));
    Odrv12 I__4167 (
            .O(N__18660),
            .I(\c0.data_in_3_Z0Z_0 ));
    LocalMux I__4166 (
            .O(N__18657),
            .I(\c0.data_in_3_Z0Z_0 ));
    CascadeMux I__4165 (
            .O(N__18650),
            .I(N__18645));
    InMux I__4164 (
            .O(N__18649),
            .I(N__18641));
    InMux I__4163 (
            .O(N__18648),
            .I(N__18637));
    InMux I__4162 (
            .O(N__18645),
            .I(N__18634));
    CascadeMux I__4161 (
            .O(N__18644),
            .I(N__18631));
    LocalMux I__4160 (
            .O(N__18641),
            .I(N__18628));
    CascadeMux I__4159 (
            .O(N__18640),
            .I(N__18623));
    LocalMux I__4158 (
            .O(N__18637),
            .I(N__18620));
    LocalMux I__4157 (
            .O(N__18634),
            .I(N__18617));
    InMux I__4156 (
            .O(N__18631),
            .I(N__18614));
    Span4Mux_h I__4155 (
            .O(N__18628),
            .I(N__18611));
    InMux I__4154 (
            .O(N__18627),
            .I(N__18604));
    InMux I__4153 (
            .O(N__18626),
            .I(N__18604));
    InMux I__4152 (
            .O(N__18623),
            .I(N__18604));
    Span4Mux_h I__4151 (
            .O(N__18620),
            .I(N__18599));
    Span4Mux_h I__4150 (
            .O(N__18617),
            .I(N__18599));
    LocalMux I__4149 (
            .O(N__18614),
            .I(\c0.d_4_24 ));
    Odrv4 I__4148 (
            .O(N__18611),
            .I(\c0.d_4_24 ));
    LocalMux I__4147 (
            .O(N__18604),
            .I(\c0.d_4_24 ));
    Odrv4 I__4146 (
            .O(N__18599),
            .I(\c0.d_4_24 ));
    InMux I__4145 (
            .O(N__18590),
            .I(N__18586));
    CascadeMux I__4144 (
            .O(N__18589),
            .I(N__18583));
    LocalMux I__4143 (
            .O(N__18586),
            .I(N__18579));
    InMux I__4142 (
            .O(N__18583),
            .I(N__18576));
    InMux I__4141 (
            .O(N__18582),
            .I(N__18573));
    Span4Mux_v I__4140 (
            .O(N__18579),
            .I(N__18569));
    LocalMux I__4139 (
            .O(N__18576),
            .I(N__18564));
    LocalMux I__4138 (
            .O(N__18573),
            .I(N__18564));
    InMux I__4137 (
            .O(N__18572),
            .I(N__18561));
    Odrv4 I__4136 (
            .O(N__18569),
            .I(\c0.N_126 ));
    Odrv4 I__4135 (
            .O(N__18564),
            .I(\c0.N_126 ));
    LocalMux I__4134 (
            .O(N__18561),
            .I(\c0.N_126 ));
    InMux I__4133 (
            .O(N__18554),
            .I(N__18551));
    LocalMux I__4132 (
            .O(N__18551),
            .I(N__18546));
    InMux I__4131 (
            .O(N__18550),
            .I(N__18541));
    InMux I__4130 (
            .O(N__18549),
            .I(N__18541));
    Odrv4 I__4129 (
            .O(N__18546),
            .I(\c0.un1_data_in_6__1_0_a2_4_a2_1 ));
    LocalMux I__4128 (
            .O(N__18541),
            .I(\c0.un1_data_in_6__1_0_a2_4_a2_1 ));
    CascadeMux I__4127 (
            .O(N__18536),
            .I(N__18533));
    InMux I__4126 (
            .O(N__18533),
            .I(N__18530));
    LocalMux I__4125 (
            .O(N__18530),
            .I(N__18527));
    Span12Mux_v I__4124 (
            .O(N__18527),
            .I(N__18524));
    Odrv12 I__4123 (
            .O(N__18524),
            .I(\c0.un1_data_in_6__1_0 ));
    InMux I__4122 (
            .O(N__18521),
            .I(N__18518));
    LocalMux I__4121 (
            .O(N__18518),
            .I(N__18515));
    Span4Mux_v I__4120 (
            .O(N__18515),
            .I(N__18512));
    Span4Mux_h I__4119 (
            .O(N__18512),
            .I(N__18508));
    InMux I__4118 (
            .O(N__18511),
            .I(N__18505));
    Odrv4 I__4117 (
            .O(N__18508),
            .I(\c0.data_in_4_Z0Z_4 ));
    LocalMux I__4116 (
            .O(N__18505),
            .I(\c0.data_in_4_Z0Z_4 ));
    CascadeMux I__4115 (
            .O(N__18500),
            .I(N__18497));
    InMux I__4114 (
            .O(N__18497),
            .I(N__18487));
    InMux I__4113 (
            .O(N__18496),
            .I(N__18487));
    CascadeMux I__4112 (
            .O(N__18495),
            .I(N__18483));
    InMux I__4111 (
            .O(N__18494),
            .I(N__18477));
    InMux I__4110 (
            .O(N__18493),
            .I(N__18477));
    InMux I__4109 (
            .O(N__18492),
            .I(N__18474));
    LocalMux I__4108 (
            .O(N__18487),
            .I(N__18471));
    InMux I__4107 (
            .O(N__18486),
            .I(N__18464));
    InMux I__4106 (
            .O(N__18483),
            .I(N__18464));
    InMux I__4105 (
            .O(N__18482),
            .I(N__18464));
    LocalMux I__4104 (
            .O(N__18477),
            .I(\c0.d_4_36 ));
    LocalMux I__4103 (
            .O(N__18474),
            .I(\c0.d_4_36 ));
    Odrv4 I__4102 (
            .O(N__18471),
            .I(\c0.d_4_36 ));
    LocalMux I__4101 (
            .O(N__18464),
            .I(\c0.d_4_36 ));
    InMux I__4100 (
            .O(N__18455),
            .I(N__18452));
    LocalMux I__4099 (
            .O(N__18452),
            .I(\c0.data_in_frame_6_Z0Z_4 ));
    InMux I__4098 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__4097 (
            .O(N__18446),
            .I(N__18443));
    Span4Mux_v I__4096 (
            .O(N__18443),
            .I(N__18440));
    Odrv4 I__4095 (
            .O(N__18440),
            .I(\c0.tx2_data_1_iv_4_1_0_6 ));
    InMux I__4094 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__4093 (
            .O(N__18434),
            .I(\c0.data_in_frame_7_Z0Z_6 ));
    InMux I__4092 (
            .O(N__18431),
            .I(N__18424));
    InMux I__4091 (
            .O(N__18430),
            .I(N__18424));
    InMux I__4090 (
            .O(N__18429),
            .I(N__18420));
    LocalMux I__4089 (
            .O(N__18424),
            .I(N__18416));
    CascadeMux I__4088 (
            .O(N__18423),
            .I(N__18413));
    LocalMux I__4087 (
            .O(N__18420),
            .I(N__18408));
    InMux I__4086 (
            .O(N__18419),
            .I(N__18405));
    Span4Mux_h I__4085 (
            .O(N__18416),
            .I(N__18402));
    InMux I__4084 (
            .O(N__18413),
            .I(N__18397));
    InMux I__4083 (
            .O(N__18412),
            .I(N__18397));
    InMux I__4082 (
            .O(N__18411),
            .I(N__18394));
    Span4Mux_h I__4081 (
            .O(N__18408),
            .I(N__18391));
    LocalMux I__4080 (
            .O(N__18405),
            .I(N__18388));
    Span4Mux_h I__4079 (
            .O(N__18402),
            .I(N__18385));
    LocalMux I__4078 (
            .O(N__18397),
            .I(N__18382));
    LocalMux I__4077 (
            .O(N__18394),
            .I(\c0.d_4_42 ));
    Odrv4 I__4076 (
            .O(N__18391),
            .I(\c0.d_4_42 ));
    Odrv12 I__4075 (
            .O(N__18388),
            .I(\c0.d_4_42 ));
    Odrv4 I__4074 (
            .O(N__18385),
            .I(\c0.d_4_42 ));
    Odrv4 I__4073 (
            .O(N__18382),
            .I(\c0.d_4_42 ));
    CascadeMux I__4072 (
            .O(N__18371),
            .I(N__18365));
    CascadeMux I__4071 (
            .O(N__18370),
            .I(N__18362));
    InMux I__4070 (
            .O(N__18369),
            .I(N__18357));
    InMux I__4069 (
            .O(N__18368),
            .I(N__18357));
    InMux I__4068 (
            .O(N__18365),
            .I(N__18352));
    InMux I__4067 (
            .O(N__18362),
            .I(N__18352));
    LocalMux I__4066 (
            .O(N__18357),
            .I(\c0.d_4_46 ));
    LocalMux I__4065 (
            .O(N__18352),
            .I(\c0.d_4_46 ));
    InMux I__4064 (
            .O(N__18347),
            .I(N__18344));
    LocalMux I__4063 (
            .O(N__18344),
            .I(N__18341));
    Span4Mux_v I__4062 (
            .O(N__18341),
            .I(N__18338));
    Odrv4 I__4061 (
            .O(N__18338),
            .I(\c0.un1_data_in_7__2_0_a2_0_a2_4 ));
    InMux I__4060 (
            .O(N__18335),
            .I(N__18331));
    InMux I__4059 (
            .O(N__18334),
            .I(N__18328));
    LocalMux I__4058 (
            .O(N__18331),
            .I(N__18323));
    LocalMux I__4057 (
            .O(N__18328),
            .I(N__18323));
    Span4Mux_v I__4056 (
            .O(N__18323),
            .I(N__18318));
    InMux I__4055 (
            .O(N__18322),
            .I(N__18313));
    InMux I__4054 (
            .O(N__18321),
            .I(N__18313));
    Odrv4 I__4053 (
            .O(N__18318),
            .I(\c0.d_4_7 ));
    LocalMux I__4052 (
            .O(N__18313),
            .I(\c0.d_4_7 ));
    InMux I__4051 (
            .O(N__18308),
            .I(N__18305));
    LocalMux I__4050 (
            .O(N__18305),
            .I(N__18302));
    Span4Mux_v I__4049 (
            .O(N__18302),
            .I(N__18298));
    InMux I__4048 (
            .O(N__18301),
            .I(N__18294));
    Span4Mux_h I__4047 (
            .O(N__18298),
            .I(N__18291));
    InMux I__4046 (
            .O(N__18297),
            .I(N__18288));
    LocalMux I__4045 (
            .O(N__18294),
            .I(\c0.data_in_1_Z0Z_0 ));
    Odrv4 I__4044 (
            .O(N__18291),
            .I(\c0.data_in_1_Z0Z_0 ));
    LocalMux I__4043 (
            .O(N__18288),
            .I(\c0.data_in_1_Z0Z_0 ));
    InMux I__4042 (
            .O(N__18281),
            .I(N__18277));
    CascadeMux I__4041 (
            .O(N__18280),
            .I(N__18274));
    LocalMux I__4040 (
            .O(N__18277),
            .I(N__18269));
    InMux I__4039 (
            .O(N__18274),
            .I(N__18262));
    InMux I__4038 (
            .O(N__18273),
            .I(N__18262));
    InMux I__4037 (
            .O(N__18272),
            .I(N__18262));
    Odrv4 I__4036 (
            .O(N__18269),
            .I(\c0.d_4_8 ));
    LocalMux I__4035 (
            .O(N__18262),
            .I(\c0.d_4_8 ));
    InMux I__4034 (
            .O(N__18257),
            .I(N__18254));
    LocalMux I__4033 (
            .O(N__18254),
            .I(N__18249));
    InMux I__4032 (
            .O(N__18253),
            .I(N__18245));
    InMux I__4031 (
            .O(N__18252),
            .I(N__18242));
    Span4Mux_v I__4030 (
            .O(N__18249),
            .I(N__18238));
    InMux I__4029 (
            .O(N__18248),
            .I(N__18235));
    LocalMux I__4028 (
            .O(N__18245),
            .I(N__18230));
    LocalMux I__4027 (
            .O(N__18242),
            .I(N__18230));
    InMux I__4026 (
            .O(N__18241),
            .I(N__18227));
    Odrv4 I__4025 (
            .O(N__18238),
            .I(\c0.d_4_9 ));
    LocalMux I__4024 (
            .O(N__18235),
            .I(\c0.d_4_9 ));
    Odrv4 I__4023 (
            .O(N__18230),
            .I(\c0.d_4_9 ));
    LocalMux I__4022 (
            .O(N__18227),
            .I(\c0.d_4_9 ));
    InMux I__4021 (
            .O(N__18218),
            .I(N__18215));
    LocalMux I__4020 (
            .O(N__18215),
            .I(N__18212));
    Span4Mux_v I__4019 (
            .O(N__18212),
            .I(N__18206));
    InMux I__4018 (
            .O(N__18211),
            .I(N__18203));
    InMux I__4017 (
            .O(N__18210),
            .I(N__18200));
    InMux I__4016 (
            .O(N__18209),
            .I(N__18197));
    Odrv4 I__4015 (
            .O(N__18206),
            .I(\c0.d_4_39 ));
    LocalMux I__4014 (
            .O(N__18203),
            .I(\c0.d_4_39 ));
    LocalMux I__4013 (
            .O(N__18200),
            .I(\c0.d_4_39 ));
    LocalMux I__4012 (
            .O(N__18197),
            .I(\c0.d_4_39 ));
    InMux I__4011 (
            .O(N__18188),
            .I(N__18185));
    LocalMux I__4010 (
            .O(N__18185),
            .I(\c0.un1_data_in_6__2_0 ));
    InMux I__4009 (
            .O(N__18182),
            .I(N__18179));
    LocalMux I__4008 (
            .O(N__18179),
            .I(N__18174));
    InMux I__4007 (
            .O(N__18178),
            .I(N__18171));
    InMux I__4006 (
            .O(N__18177),
            .I(N__18168));
    Span4Mux_h I__4005 (
            .O(N__18174),
            .I(N__18165));
    LocalMux I__4004 (
            .O(N__18171),
            .I(N__18162));
    LocalMux I__4003 (
            .O(N__18168),
            .I(\c0.N_107 ));
    Odrv4 I__4002 (
            .O(N__18165),
            .I(\c0.N_107 ));
    Odrv4 I__4001 (
            .O(N__18162),
            .I(\c0.N_107 ));
    InMux I__4000 (
            .O(N__18155),
            .I(N__18149));
    InMux I__3999 (
            .O(N__18154),
            .I(N__18149));
    LocalMux I__3998 (
            .O(N__18149),
            .I(\c0.un1_data_in_6__2_0_a2_6_a2_2 ));
    CascadeMux I__3997 (
            .O(N__18146),
            .I(\c0.N_107_cascade_ ));
    InMux I__3996 (
            .O(N__18143),
            .I(N__18140));
    LocalMux I__3995 (
            .O(N__18140),
            .I(N__18136));
    InMux I__3994 (
            .O(N__18139),
            .I(N__18133));
    Span4Mux_h I__3993 (
            .O(N__18136),
            .I(N__18130));
    LocalMux I__3992 (
            .O(N__18133),
            .I(N__18127));
    Odrv4 I__3991 (
            .O(N__18130),
            .I(\c0.un1_data_in_6__2 ));
    Odrv4 I__3990 (
            .O(N__18127),
            .I(\c0.un1_data_in_6__2 ));
    InMux I__3989 (
            .O(N__18122),
            .I(N__18118));
    InMux I__3988 (
            .O(N__18121),
            .I(N__18115));
    LocalMux I__3987 (
            .O(N__18118),
            .I(N__18111));
    LocalMux I__3986 (
            .O(N__18115),
            .I(N__18108));
    InMux I__3985 (
            .O(N__18114),
            .I(N__18105));
    Span4Mux_h I__3984 (
            .O(N__18111),
            .I(N__18102));
    Span4Mux_h I__3983 (
            .O(N__18108),
            .I(N__18099));
    LocalMux I__3982 (
            .O(N__18105),
            .I(\c0.data_in_2_Z0Z_6 ));
    Odrv4 I__3981 (
            .O(N__18102),
            .I(\c0.data_in_2_Z0Z_6 ));
    Odrv4 I__3980 (
            .O(N__18099),
            .I(\c0.data_in_2_Z0Z_6 ));
    InMux I__3979 (
            .O(N__18092),
            .I(N__18089));
    LocalMux I__3978 (
            .O(N__18089),
            .I(N__18086));
    Span4Mux_h I__3977 (
            .O(N__18086),
            .I(N__18080));
    InMux I__3976 (
            .O(N__18085),
            .I(N__18073));
    InMux I__3975 (
            .O(N__18084),
            .I(N__18073));
    InMux I__3974 (
            .O(N__18083),
            .I(N__18073));
    Odrv4 I__3973 (
            .O(N__18080),
            .I(\c0.d_4_22 ));
    LocalMux I__3972 (
            .O(N__18073),
            .I(\c0.d_4_22 ));
    CascadeMux I__3971 (
            .O(N__18068),
            .I(\c0.d_4_RNI9LFUVZ0Z_43_cascade_ ));
    CascadeMux I__3970 (
            .O(N__18065),
            .I(\c0.wait_for_transmission_RNI9PP5BZ0Z1_cascade_ ));
    InMux I__3969 (
            .O(N__18062),
            .I(N__18059));
    LocalMux I__3968 (
            .O(N__18059),
            .I(N__18056));
    Span4Mux_v I__3967 (
            .O(N__18056),
            .I(N__18053));
    Odrv4 I__3966 (
            .O(N__18053),
            .I(\c0.un1_data_in_6__1_1 ));
    InMux I__3965 (
            .O(N__18050),
            .I(N__18047));
    LocalMux I__3964 (
            .O(N__18047),
            .I(\c0.g0_2_3 ));
    InMux I__3963 (
            .O(N__18044),
            .I(N__18041));
    LocalMux I__3962 (
            .O(N__18041),
            .I(N__18037));
    CascadeMux I__3961 (
            .O(N__18040),
            .I(N__18032));
    Span4Mux_v I__3960 (
            .O(N__18037),
            .I(N__18029));
    InMux I__3959 (
            .O(N__18036),
            .I(N__18026));
    InMux I__3958 (
            .O(N__18035),
            .I(N__18021));
    InMux I__3957 (
            .O(N__18032),
            .I(N__18021));
    Odrv4 I__3956 (
            .O(N__18029),
            .I(\c0.d_4_23 ));
    LocalMux I__3955 (
            .O(N__18026),
            .I(\c0.d_4_23 ));
    LocalMux I__3954 (
            .O(N__18021),
            .I(\c0.d_4_23 ));
    CascadeMux I__3953 (
            .O(N__18014),
            .I(\c0.N_126_cascade_ ));
    InMux I__3952 (
            .O(N__18011),
            .I(N__18008));
    LocalMux I__3951 (
            .O(N__18008),
            .I(\c0.un1_data_in_6__1 ));
    InMux I__3950 (
            .O(N__18005),
            .I(N__18000));
    InMux I__3949 (
            .O(N__18004),
            .I(N__17996));
    InMux I__3948 (
            .O(N__18003),
            .I(N__17992));
    LocalMux I__3947 (
            .O(N__18000),
            .I(N__17988));
    InMux I__3946 (
            .O(N__17999),
            .I(N__17985));
    LocalMux I__3945 (
            .O(N__17996),
            .I(N__17982));
    InMux I__3944 (
            .O(N__17995),
            .I(N__17979));
    LocalMux I__3943 (
            .O(N__17992),
            .I(N__17976));
    InMux I__3942 (
            .O(N__17991),
            .I(N__17973));
    Odrv4 I__3941 (
            .O(N__17988),
            .I(\c0.d_4_35 ));
    LocalMux I__3940 (
            .O(N__17985),
            .I(\c0.d_4_35 ));
    Odrv4 I__3939 (
            .O(N__17982),
            .I(\c0.d_4_35 ));
    LocalMux I__3938 (
            .O(N__17979),
            .I(\c0.d_4_35 ));
    Odrv4 I__3937 (
            .O(N__17976),
            .I(\c0.d_4_35 ));
    LocalMux I__3936 (
            .O(N__17973),
            .I(\c0.d_4_35 ));
    InMux I__3935 (
            .O(N__17960),
            .I(N__17957));
    LocalMux I__3934 (
            .O(N__17957),
            .I(N__17953));
    InMux I__3933 (
            .O(N__17956),
            .I(N__17950));
    Odrv12 I__3932 (
            .O(N__17953),
            .I(\c0.data_in_0_Z0Z_7 ));
    LocalMux I__3931 (
            .O(N__17950),
            .I(\c0.data_in_0_Z0Z_7 ));
    InMux I__3930 (
            .O(N__17945),
            .I(N__17942));
    LocalMux I__3929 (
            .O(N__17942),
            .I(N__17938));
    CascadeMux I__3928 (
            .O(N__17941),
            .I(N__17934));
    Span4Mux_v I__3927 (
            .O(N__17938),
            .I(N__17931));
    InMux I__3926 (
            .O(N__17937),
            .I(N__17926));
    InMux I__3925 (
            .O(N__17934),
            .I(N__17926));
    Odrv4 I__3924 (
            .O(N__17931),
            .I(\c0.d_4_15 ));
    LocalMux I__3923 (
            .O(N__17926),
            .I(\c0.d_4_15 ));
    CascadeMux I__3922 (
            .O(N__17921),
            .I(\c0.data_in_frame_1__m_7_cascade_ ));
    InMux I__3921 (
            .O(N__17918),
            .I(N__17914));
    InMux I__3920 (
            .O(N__17917),
            .I(N__17911));
    LocalMux I__3919 (
            .O(N__17914),
            .I(N__17906));
    LocalMux I__3918 (
            .O(N__17911),
            .I(N__17906));
    Span4Mux_h I__3917 (
            .O(N__17906),
            .I(N__17897));
    InMux I__3916 (
            .O(N__17905),
            .I(N__17890));
    InMux I__3915 (
            .O(N__17904),
            .I(N__17890));
    InMux I__3914 (
            .O(N__17903),
            .I(N__17890));
    InMux I__3913 (
            .O(N__17902),
            .I(N__17883));
    InMux I__3912 (
            .O(N__17901),
            .I(N__17883));
    InMux I__3911 (
            .O(N__17900),
            .I(N__17883));
    Odrv4 I__3910 (
            .O(N__17897),
            .I(\c0.d_4_31 ));
    LocalMux I__3909 (
            .O(N__17890),
            .I(\c0.d_4_31 ));
    LocalMux I__3908 (
            .O(N__17883),
            .I(\c0.d_4_31 ));
    InMux I__3907 (
            .O(N__17876),
            .I(N__17873));
    LocalMux I__3906 (
            .O(N__17873),
            .I(\c0.tx2_data_1_iv_1_7 ));
    InMux I__3905 (
            .O(N__17870),
            .I(N__17866));
    CascadeMux I__3904 (
            .O(N__17869),
            .I(N__17862));
    LocalMux I__3903 (
            .O(N__17866),
            .I(N__17859));
    InMux I__3902 (
            .O(N__17865),
            .I(N__17851));
    InMux I__3901 (
            .O(N__17862),
            .I(N__17851));
    Span4Mux_h I__3900 (
            .O(N__17859),
            .I(N__17847));
    CascadeMux I__3899 (
            .O(N__17858),
            .I(N__17844));
    InMux I__3898 (
            .O(N__17857),
            .I(N__17839));
    InMux I__3897 (
            .O(N__17856),
            .I(N__17839));
    LocalMux I__3896 (
            .O(N__17851),
            .I(N__17836));
    CascadeMux I__3895 (
            .O(N__17850),
            .I(N__17832));
    Span4Mux_h I__3894 (
            .O(N__17847),
            .I(N__17829));
    InMux I__3893 (
            .O(N__17844),
            .I(N__17826));
    LocalMux I__3892 (
            .O(N__17839),
            .I(N__17821));
    Span12Mux_v I__3891 (
            .O(N__17836),
            .I(N__17821));
    InMux I__3890 (
            .O(N__17835),
            .I(N__17816));
    InMux I__3889 (
            .O(N__17832),
            .I(N__17816));
    Odrv4 I__3888 (
            .O(N__17829),
            .I(\c0.N_205 ));
    LocalMux I__3887 (
            .O(N__17826),
            .I(\c0.N_205 ));
    Odrv12 I__3886 (
            .O(N__17821),
            .I(\c0.N_205 ));
    LocalMux I__3885 (
            .O(N__17816),
            .I(\c0.N_205 ));
    InMux I__3884 (
            .O(N__17807),
            .I(N__17804));
    LocalMux I__3883 (
            .O(N__17804),
            .I(N__17801));
    Span4Mux_h I__3882 (
            .O(N__17801),
            .I(N__17795));
    InMux I__3881 (
            .O(N__17800),
            .I(N__17790));
    InMux I__3880 (
            .O(N__17799),
            .I(N__17790));
    InMux I__3879 (
            .O(N__17798),
            .I(N__17787));
    Odrv4 I__3878 (
            .O(N__17795),
            .I(\c0.d_4_27 ));
    LocalMux I__3877 (
            .O(N__17790),
            .I(\c0.d_4_27 ));
    LocalMux I__3876 (
            .O(N__17787),
            .I(\c0.d_4_27 ));
    CascadeMux I__3875 (
            .O(N__17780),
            .I(\c0.N_205_cascade_ ));
    InMux I__3874 (
            .O(N__17777),
            .I(N__17774));
    LocalMux I__3873 (
            .O(N__17774),
            .I(N__17771));
    Span4Mux_h I__3872 (
            .O(N__17771),
            .I(N__17767));
    InMux I__3871 (
            .O(N__17770),
            .I(N__17764));
    Odrv4 I__3870 (
            .O(N__17767),
            .I(\c0.d_4_11 ));
    LocalMux I__3869 (
            .O(N__17764),
            .I(\c0.d_4_11 ));
    InMux I__3868 (
            .O(N__17759),
            .I(N__17756));
    LocalMux I__3867 (
            .O(N__17756),
            .I(N__17753));
    Span4Mux_h I__3866 (
            .O(N__17753),
            .I(N__17750));
    Span4Mux_h I__3865 (
            .O(N__17750),
            .I(N__17747));
    Odrv4 I__3864 (
            .O(N__17747),
            .I(\c0.tx2_data_1_iv_4_1_3 ));
    InMux I__3863 (
            .O(N__17744),
            .I(N__17740));
    CascadeMux I__3862 (
            .O(N__17743),
            .I(N__17737));
    LocalMux I__3861 (
            .O(N__17740),
            .I(N__17734));
    InMux I__3860 (
            .O(N__17737),
            .I(N__17731));
    Odrv4 I__3859 (
            .O(N__17734),
            .I(\c0.un1_data_in_6__5 ));
    LocalMux I__3858 (
            .O(N__17731),
            .I(\c0.un1_data_in_6__5 ));
    InMux I__3857 (
            .O(N__17726),
            .I(N__17721));
    InMux I__3856 (
            .O(N__17725),
            .I(N__17718));
    InMux I__3855 (
            .O(N__17724),
            .I(N__17715));
    LocalMux I__3854 (
            .O(N__17721),
            .I(N__17712));
    LocalMux I__3853 (
            .O(N__17718),
            .I(\c0.i12_THRU_CO ));
    LocalMux I__3852 (
            .O(N__17715),
            .I(\c0.i12_THRU_CO ));
    Odrv12 I__3851 (
            .O(N__17712),
            .I(\c0.i12_THRU_CO ));
    InMux I__3850 (
            .O(N__17705),
            .I(N__17701));
    InMux I__3849 (
            .O(N__17704),
            .I(N__17698));
    LocalMux I__3848 (
            .O(N__17701),
            .I(\c0.N_136 ));
    LocalMux I__3847 (
            .O(N__17698),
            .I(\c0.N_136 ));
    InMux I__3846 (
            .O(N__17693),
            .I(N__17688));
    InMux I__3845 (
            .O(N__17692),
            .I(N__17685));
    InMux I__3844 (
            .O(N__17691),
            .I(N__17682));
    LocalMux I__3843 (
            .O(N__17688),
            .I(N__17679));
    LocalMux I__3842 (
            .O(N__17685),
            .I(N__17676));
    LocalMux I__3841 (
            .O(N__17682),
            .I(N__17673));
    Span4Mux_v I__3840 (
            .O(N__17679),
            .I(N__17670));
    Odrv4 I__3839 (
            .O(N__17676),
            .I(\c0.wait_for_transmission4_13_1 ));
    Odrv4 I__3838 (
            .O(N__17673),
            .I(\c0.wait_for_transmission4_13_1 ));
    Odrv4 I__3837 (
            .O(N__17670),
            .I(\c0.wait_for_transmission4_13_1 ));
    CascadeMux I__3836 (
            .O(N__17663),
            .I(\c0.g1_3_cascade_ ));
    InMux I__3835 (
            .O(N__17660),
            .I(N__17657));
    LocalMux I__3834 (
            .O(N__17657),
            .I(N__17654));
    Span4Mux_v I__3833 (
            .O(N__17654),
            .I(N__17650));
    InMux I__3832 (
            .O(N__17653),
            .I(N__17647));
    Span4Mux_h I__3831 (
            .O(N__17650),
            .I(N__17642));
    LocalMux I__3830 (
            .O(N__17647),
            .I(N__17642));
    Sp12to4 I__3829 (
            .O(N__17642),
            .I(N__17639));
    Odrv12 I__3828 (
            .O(N__17639),
            .I(\c0.un1_data_in_7__0_0_a2_1_a2_5_0 ));
    CascadeMux I__3827 (
            .O(N__17636),
            .I(\c0.i12_7_c_RNIP740G_cascade_ ));
    InMux I__3826 (
            .O(N__17633),
            .I(N__17630));
    LocalMux I__3825 (
            .O(N__17630),
            .I(\c0.g1_2 ));
    InMux I__3824 (
            .O(N__17627),
            .I(N__17624));
    LocalMux I__3823 (
            .O(N__17624),
            .I(N__17621));
    Span4Mux_v I__3822 (
            .O(N__17621),
            .I(N__17617));
    InMux I__3821 (
            .O(N__17620),
            .I(N__17614));
    Odrv4 I__3820 (
            .O(N__17617),
            .I(\c0.wait_for_transmission4_12_5 ));
    LocalMux I__3819 (
            .O(N__17614),
            .I(\c0.wait_for_transmission4_12_5 ));
    InMux I__3818 (
            .O(N__17609),
            .I(N__17606));
    LocalMux I__3817 (
            .O(N__17606),
            .I(N__17602));
    InMux I__3816 (
            .O(N__17605),
            .I(N__17599));
    Span4Mux_v I__3815 (
            .O(N__17602),
            .I(N__17596));
    LocalMux I__3814 (
            .O(N__17599),
            .I(\c0.un1_data_in_7__3_i ));
    Odrv4 I__3813 (
            .O(N__17596),
            .I(\c0.un1_data_in_7__3_i ));
    CascadeMux I__3812 (
            .O(N__17591),
            .I(\c0.g1_5_cascade_ ));
    InMux I__3811 (
            .O(N__17588),
            .I(N__17584));
    InMux I__3810 (
            .O(N__17587),
            .I(N__17581));
    LocalMux I__3809 (
            .O(N__17584),
            .I(N__17578));
    LocalMux I__3808 (
            .O(N__17581),
            .I(\c0.wait_for_transmission4_12_4 ));
    Odrv4 I__3807 (
            .O(N__17578),
            .I(\c0.wait_for_transmission4_12_4 ));
    InMux I__3806 (
            .O(N__17573),
            .I(N__17570));
    LocalMux I__3805 (
            .O(N__17570),
            .I(\c0.byte_transmit_counterZ0Z_4 ));
    InMux I__3804 (
            .O(N__17567),
            .I(N__17558));
    InMux I__3803 (
            .O(N__17566),
            .I(N__17555));
    InMux I__3802 (
            .O(N__17565),
            .I(N__17550));
    InMux I__3801 (
            .O(N__17564),
            .I(N__17547));
    InMux I__3800 (
            .O(N__17563),
            .I(N__17544));
    InMux I__3799 (
            .O(N__17562),
            .I(N__17541));
    InMux I__3798 (
            .O(N__17561),
            .I(N__17537));
    LocalMux I__3797 (
            .O(N__17558),
            .I(N__17534));
    LocalMux I__3796 (
            .O(N__17555),
            .I(N__17531));
    InMux I__3795 (
            .O(N__17554),
            .I(N__17528));
    InMux I__3794 (
            .O(N__17553),
            .I(N__17525));
    LocalMux I__3793 (
            .O(N__17550),
            .I(N__17522));
    LocalMux I__3792 (
            .O(N__17547),
            .I(N__17517));
    LocalMux I__3791 (
            .O(N__17544),
            .I(N__17512));
    LocalMux I__3790 (
            .O(N__17541),
            .I(N__17512));
    InMux I__3789 (
            .O(N__17540),
            .I(N__17509));
    LocalMux I__3788 (
            .O(N__17537),
            .I(N__17506));
    Span4Mux_v I__3787 (
            .O(N__17534),
            .I(N__17492));
    Span4Mux_v I__3786 (
            .O(N__17531),
            .I(N__17492));
    LocalMux I__3785 (
            .O(N__17528),
            .I(N__17492));
    LocalMux I__3784 (
            .O(N__17525),
            .I(N__17492));
    Span4Mux_v I__3783 (
            .O(N__17522),
            .I(N__17492));
    InMux I__3782 (
            .O(N__17521),
            .I(N__17489));
    InMux I__3781 (
            .O(N__17520),
            .I(N__17486));
    Span4Mux_v I__3780 (
            .O(N__17517),
            .I(N__17483));
    Span4Mux_v I__3779 (
            .O(N__17512),
            .I(N__17476));
    LocalMux I__3778 (
            .O(N__17509),
            .I(N__17476));
    Span4Mux_h I__3777 (
            .O(N__17506),
            .I(N__17476));
    InMux I__3776 (
            .O(N__17505),
            .I(N__17470));
    InMux I__3775 (
            .O(N__17504),
            .I(N__17470));
    InMux I__3774 (
            .O(N__17503),
            .I(N__17467));
    Span4Mux_h I__3773 (
            .O(N__17492),
            .I(N__17462));
    LocalMux I__3772 (
            .O(N__17489),
            .I(N__17462));
    LocalMux I__3771 (
            .O(N__17486),
            .I(N__17455));
    Span4Mux_h I__3770 (
            .O(N__17483),
            .I(N__17455));
    Span4Mux_h I__3769 (
            .O(N__17476),
            .I(N__17455));
    InMux I__3768 (
            .O(N__17475),
            .I(N__17452));
    LocalMux I__3767 (
            .O(N__17470),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    LocalMux I__3766 (
            .O(N__17467),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    Odrv4 I__3765 (
            .O(N__17462),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    Odrv4 I__3764 (
            .O(N__17455),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    LocalMux I__3763 (
            .O(N__17452),
            .I(\c0.byte_transmit_counterZ0Z_0 ));
    InMux I__3762 (
            .O(N__17441),
            .I(N__17438));
    LocalMux I__3761 (
            .O(N__17438),
            .I(\c0.un144_newcrc_3 ));
    InMux I__3760 (
            .O(N__17435),
            .I(N__17430));
    InMux I__3759 (
            .O(N__17434),
            .I(N__17427));
    InMux I__3758 (
            .O(N__17433),
            .I(N__17424));
    LocalMux I__3757 (
            .O(N__17430),
            .I(N__17419));
    LocalMux I__3756 (
            .O(N__17427),
            .I(N__17419));
    LocalMux I__3755 (
            .O(N__17424),
            .I(N__17415));
    Span4Mux_h I__3754 (
            .O(N__17419),
            .I(N__17412));
    InMux I__3753 (
            .O(N__17418),
            .I(N__17409));
    Odrv12 I__3752 (
            .O(N__17415),
            .I(\c0.d_2_34 ));
    Odrv4 I__3751 (
            .O(N__17412),
            .I(\c0.d_2_34 ));
    LocalMux I__3750 (
            .O(N__17409),
            .I(\c0.d_2_34 ));
    CascadeMux I__3749 (
            .O(N__17402),
            .I(N__17399));
    InMux I__3748 (
            .O(N__17399),
            .I(N__17396));
    LocalMux I__3747 (
            .O(N__17396),
            .I(\c0.un144_newcrc_4 ));
    InMux I__3746 (
            .O(N__17393),
            .I(N__17389));
    CascadeMux I__3745 (
            .O(N__17392),
            .I(N__17386));
    LocalMux I__3744 (
            .O(N__17389),
            .I(N__17383));
    InMux I__3743 (
            .O(N__17386),
            .I(N__17380));
    Span4Mux_v I__3742 (
            .O(N__17383),
            .I(N__17373));
    LocalMux I__3741 (
            .O(N__17380),
            .I(N__17373));
    InMux I__3740 (
            .O(N__17379),
            .I(N__17370));
    InMux I__3739 (
            .O(N__17378),
            .I(N__17367));
    Span4Mux_h I__3738 (
            .O(N__17373),
            .I(N__17362));
    LocalMux I__3737 (
            .O(N__17370),
            .I(N__17362));
    LocalMux I__3736 (
            .O(N__17367),
            .I(\c0.d_2_33 ));
    Odrv4 I__3735 (
            .O(N__17362),
            .I(\c0.d_2_33 ));
    InMux I__3734 (
            .O(N__17357),
            .I(N__17354));
    LocalMux I__3733 (
            .O(N__17354),
            .I(N__17351));
    Odrv4 I__3732 (
            .O(N__17351),
            .I(\c0.data_out_7_Z0Z_6 ));
    SRMux I__3731 (
            .O(N__17348),
            .I(N__17334));
    SRMux I__3730 (
            .O(N__17347),
            .I(N__17331));
    SRMux I__3729 (
            .O(N__17346),
            .I(N__17328));
    SRMux I__3728 (
            .O(N__17345),
            .I(N__17325));
    SRMux I__3727 (
            .O(N__17344),
            .I(N__17322));
    SRMux I__3726 (
            .O(N__17343),
            .I(N__17319));
    SRMux I__3725 (
            .O(N__17342),
            .I(N__17316));
    SRMux I__3724 (
            .O(N__17341),
            .I(N__17313));
    SRMux I__3723 (
            .O(N__17340),
            .I(N__17310));
    SRMux I__3722 (
            .O(N__17339),
            .I(N__17307));
    SRMux I__3721 (
            .O(N__17338),
            .I(N__17304));
    SRMux I__3720 (
            .O(N__17337),
            .I(N__17301));
    LocalMux I__3719 (
            .O(N__17334),
            .I(N__17284));
    LocalMux I__3718 (
            .O(N__17331),
            .I(N__17281));
    LocalMux I__3717 (
            .O(N__17328),
            .I(N__17278));
    LocalMux I__3716 (
            .O(N__17325),
            .I(N__17275));
    LocalMux I__3715 (
            .O(N__17322),
            .I(N__17272));
    LocalMux I__3714 (
            .O(N__17319),
            .I(N__17269));
    LocalMux I__3713 (
            .O(N__17316),
            .I(N__17266));
    LocalMux I__3712 (
            .O(N__17313),
            .I(N__17263));
    LocalMux I__3711 (
            .O(N__17310),
            .I(N__17260));
    LocalMux I__3710 (
            .O(N__17307),
            .I(N__17257));
    LocalMux I__3709 (
            .O(N__17304),
            .I(N__17254));
    LocalMux I__3708 (
            .O(N__17301),
            .I(N__17251));
    CEMux I__3707 (
            .O(N__17300),
            .I(N__17198));
    CEMux I__3706 (
            .O(N__17299),
            .I(N__17198));
    CEMux I__3705 (
            .O(N__17298),
            .I(N__17198));
    CEMux I__3704 (
            .O(N__17297),
            .I(N__17198));
    CEMux I__3703 (
            .O(N__17296),
            .I(N__17198));
    CEMux I__3702 (
            .O(N__17295),
            .I(N__17198));
    CEMux I__3701 (
            .O(N__17294),
            .I(N__17198));
    CEMux I__3700 (
            .O(N__17293),
            .I(N__17198));
    CEMux I__3699 (
            .O(N__17292),
            .I(N__17198));
    CEMux I__3698 (
            .O(N__17291),
            .I(N__17198));
    CEMux I__3697 (
            .O(N__17290),
            .I(N__17198));
    CEMux I__3696 (
            .O(N__17289),
            .I(N__17198));
    CEMux I__3695 (
            .O(N__17288),
            .I(N__17198));
    CEMux I__3694 (
            .O(N__17287),
            .I(N__17198));
    Glb2LocalMux I__3693 (
            .O(N__17284),
            .I(N__17198));
    Glb2LocalMux I__3692 (
            .O(N__17281),
            .I(N__17198));
    Glb2LocalMux I__3691 (
            .O(N__17278),
            .I(N__17198));
    Glb2LocalMux I__3690 (
            .O(N__17275),
            .I(N__17198));
    Glb2LocalMux I__3689 (
            .O(N__17272),
            .I(N__17198));
    Glb2LocalMux I__3688 (
            .O(N__17269),
            .I(N__17198));
    Glb2LocalMux I__3687 (
            .O(N__17266),
            .I(N__17198));
    Glb2LocalMux I__3686 (
            .O(N__17263),
            .I(N__17198));
    Glb2LocalMux I__3685 (
            .O(N__17260),
            .I(N__17198));
    Glb2LocalMux I__3684 (
            .O(N__17257),
            .I(N__17198));
    Glb2LocalMux I__3683 (
            .O(N__17254),
            .I(N__17198));
    Glb2LocalMux I__3682 (
            .O(N__17251),
            .I(N__17198));
    GlobalMux I__3681 (
            .O(N__17198),
            .I(N__17195));
    gio2CtrlBuf I__3680 (
            .O(N__17195),
            .I(\c0.data_out_0__1_sqmuxa_g ));
    InMux I__3679 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__3678 (
            .O(N__17189),
            .I(N__17185));
    InMux I__3677 (
            .O(N__17188),
            .I(N__17181));
    Span4Mux_v I__3676 (
            .O(N__17185),
            .I(N__17175));
    InMux I__3675 (
            .O(N__17184),
            .I(N__17172));
    LocalMux I__3674 (
            .O(N__17181),
            .I(N__17168));
    InMux I__3673 (
            .O(N__17180),
            .I(N__17161));
    InMux I__3672 (
            .O(N__17179),
            .I(N__17161));
    InMux I__3671 (
            .O(N__17178),
            .I(N__17161));
    Span4Mux_v I__3670 (
            .O(N__17175),
            .I(N__17158));
    LocalMux I__3669 (
            .O(N__17172),
            .I(N__17155));
    InMux I__3668 (
            .O(N__17171),
            .I(N__17152));
    Span4Mux_h I__3667 (
            .O(N__17168),
            .I(N__17147));
    LocalMux I__3666 (
            .O(N__17161),
            .I(N__17147));
    Odrv4 I__3665 (
            .O(N__17158),
            .I(\c0.d_4_12 ));
    Odrv4 I__3664 (
            .O(N__17155),
            .I(\c0.d_4_12 ));
    LocalMux I__3663 (
            .O(N__17152),
            .I(\c0.d_4_12 ));
    Odrv4 I__3662 (
            .O(N__17147),
            .I(\c0.d_4_12 ));
    InMux I__3661 (
            .O(N__17138),
            .I(N__17135));
    LocalMux I__3660 (
            .O(N__17135),
            .I(N__17132));
    Span4Mux_h I__3659 (
            .O(N__17132),
            .I(N__17129));
    Span4Mux_v I__3658 (
            .O(N__17129),
            .I(N__17122));
    InMux I__3657 (
            .O(N__17128),
            .I(N__17119));
    InMux I__3656 (
            .O(N__17127),
            .I(N__17116));
    InMux I__3655 (
            .O(N__17126),
            .I(N__17111));
    InMux I__3654 (
            .O(N__17125),
            .I(N__17111));
    Odrv4 I__3653 (
            .O(N__17122),
            .I(\c0.d_4_44 ));
    LocalMux I__3652 (
            .O(N__17119),
            .I(\c0.d_4_44 ));
    LocalMux I__3651 (
            .O(N__17116),
            .I(\c0.d_4_44 ));
    LocalMux I__3650 (
            .O(N__17111),
            .I(\c0.d_4_44 ));
    InMux I__3649 (
            .O(N__17102),
            .I(N__17099));
    LocalMux I__3648 (
            .O(N__17099),
            .I(N__17096));
    Odrv12 I__3647 (
            .O(N__17096),
            .I(\c0.tx2_data_1_iv_5_7 ));
    CascadeMux I__3646 (
            .O(N__17093),
            .I(N__17090));
    InMux I__3645 (
            .O(N__17090),
            .I(N__17087));
    LocalMux I__3644 (
            .O(N__17087),
            .I(N__17084));
    Odrv12 I__3643 (
            .O(N__17084),
            .I(\c0.tx2_data_1_0_i_1_7 ));
    InMux I__3642 (
            .O(N__17081),
            .I(N__17078));
    LocalMux I__3641 (
            .O(N__17078),
            .I(N__17075));
    Span4Mux_h I__3640 (
            .O(N__17075),
            .I(N__17072));
    Span4Mux_v I__3639 (
            .O(N__17072),
            .I(N__17069));
    Odrv4 I__3638 (
            .O(N__17069),
            .I(\c0.tx2.r_Tx_DataZ0Z_7 ));
    InMux I__3637 (
            .O(N__17066),
            .I(N__17063));
    LocalMux I__3636 (
            .O(N__17063),
            .I(N__17059));
    InMux I__3635 (
            .O(N__17062),
            .I(N__17056));
    Span4Mux_h I__3634 (
            .O(N__17059),
            .I(N__17050));
    LocalMux I__3633 (
            .O(N__17056),
            .I(N__17050));
    InMux I__3632 (
            .O(N__17055),
            .I(N__17047));
    Odrv4 I__3631 (
            .O(N__17050),
            .I(\c0.d_4_13 ));
    LocalMux I__3630 (
            .O(N__17047),
            .I(\c0.d_4_13 ));
    InMux I__3629 (
            .O(N__17042),
            .I(N__17039));
    LocalMux I__3628 (
            .O(N__17039),
            .I(N__17036));
    Span4Mux_h I__3627 (
            .O(N__17036),
            .I(N__17032));
    InMux I__3626 (
            .O(N__17035),
            .I(N__17029));
    Span4Mux_h I__3625 (
            .O(N__17032),
            .I(N__17024));
    LocalMux I__3624 (
            .O(N__17029),
            .I(N__17024));
    Span4Mux_v I__3623 (
            .O(N__17024),
            .I(N__17019));
    CascadeMux I__3622 (
            .O(N__17023),
            .I(N__17016));
    InMux I__3621 (
            .O(N__17022),
            .I(N__17012));
    Span4Mux_h I__3620 (
            .O(N__17019),
            .I(N__17009));
    InMux I__3619 (
            .O(N__17016),
            .I(N__17004));
    InMux I__3618 (
            .O(N__17015),
            .I(N__17004));
    LocalMux I__3617 (
            .O(N__17012),
            .I(\c0.d_4_29 ));
    Odrv4 I__3616 (
            .O(N__17009),
            .I(\c0.d_4_29 ));
    LocalMux I__3615 (
            .O(N__17004),
            .I(\c0.d_4_29 ));
    CascadeMux I__3614 (
            .O(N__16997),
            .I(\c0.data_in_frame_1__m_5_cascade_ ));
    InMux I__3613 (
            .O(N__16994),
            .I(N__16991));
    LocalMux I__3612 (
            .O(N__16991),
            .I(N__16988));
    Odrv4 I__3611 (
            .O(N__16988),
            .I(\c0.tx2_data_1_0_i_1_5 ));
    CascadeMux I__3610 (
            .O(N__16985),
            .I(\c0.tx2_data_1_iv_1_5_cascade_ ));
    InMux I__3609 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__3608 (
            .O(N__16979),
            .I(N__16976));
    Span4Mux_v I__3607 (
            .O(N__16976),
            .I(N__16973));
    Span4Mux_v I__3606 (
            .O(N__16973),
            .I(N__16970));
    Odrv4 I__3605 (
            .O(N__16970),
            .I(\c0.tx2.r_Tx_DataZ0Z_5 ));
    InMux I__3604 (
            .O(N__16967),
            .I(N__16964));
    LocalMux I__3603 (
            .O(N__16964),
            .I(\c0.data_out_6_Z0Z_6 ));
    CascadeMux I__3602 (
            .O(N__16961),
            .I(\c0.N_4_0_cascade_ ));
    InMux I__3601 (
            .O(N__16958),
            .I(N__16955));
    LocalMux I__3600 (
            .O(N__16955),
            .I(N__16952));
    Odrv12 I__3599 (
            .O(N__16952),
            .I(\c0.N_197 ));
    IoInMux I__3598 (
            .O(N__16949),
            .I(N__16946));
    LocalMux I__3597 (
            .O(N__16946),
            .I(N__16943));
    IoSpan4Mux I__3596 (
            .O(N__16943),
            .I(N__16940));
    Span4Mux_s1_v I__3595 (
            .O(N__16940),
            .I(N__16937));
    Span4Mux_v I__3594 (
            .O(N__16937),
            .I(N__16934));
    Odrv4 I__3593 (
            .O(N__16934),
            .I(\c0.data_out_0__1_sqmuxa ));
    InMux I__3592 (
            .O(N__16931),
            .I(N__16928));
    LocalMux I__3591 (
            .O(N__16928),
            .I(\c0.byte_transmit_counterZ0Z_6 ));
    InMux I__3590 (
            .O(N__16925),
            .I(N__16922));
    LocalMux I__3589 (
            .O(N__16922),
            .I(\c0.byte_transmit_counterZ0Z_3 ));
    CascadeMux I__3588 (
            .O(N__16919),
            .I(\c0.m2_e_1_cascade_ ));
    CascadeMux I__3587 (
            .O(N__16916),
            .I(\c0.N_129_mux_cascade_ ));
    InMux I__3586 (
            .O(N__16913),
            .I(N__16910));
    LocalMux I__3585 (
            .O(N__16910),
            .I(N__16905));
    InMux I__3584 (
            .O(N__16909),
            .I(N__16902));
    InMux I__3583 (
            .O(N__16908),
            .I(N__16899));
    Span4Mux_h I__3582 (
            .O(N__16905),
            .I(N__16894));
    LocalMux I__3581 (
            .O(N__16902),
            .I(N__16894));
    LocalMux I__3580 (
            .O(N__16899),
            .I(N__16891));
    Span4Mux_h I__3579 (
            .O(N__16894),
            .I(N__16888));
    Odrv12 I__3578 (
            .O(N__16891),
            .I(\c0.N_86 ));
    Odrv4 I__3577 (
            .O(N__16888),
            .I(\c0.N_86 ));
    InMux I__3576 (
            .O(N__16883),
            .I(N__16878));
    CascadeMux I__3575 (
            .O(N__16882),
            .I(N__16872));
    InMux I__3574 (
            .O(N__16881),
            .I(N__16864));
    LocalMux I__3573 (
            .O(N__16878),
            .I(N__16861));
    InMux I__3572 (
            .O(N__16877),
            .I(N__16856));
    InMux I__3571 (
            .O(N__16876),
            .I(N__16856));
    InMux I__3570 (
            .O(N__16875),
            .I(N__16851));
    InMux I__3569 (
            .O(N__16872),
            .I(N__16851));
    InMux I__3568 (
            .O(N__16871),
            .I(N__16844));
    InMux I__3567 (
            .O(N__16870),
            .I(N__16844));
    InMux I__3566 (
            .O(N__16869),
            .I(N__16844));
    InMux I__3565 (
            .O(N__16868),
            .I(N__16839));
    InMux I__3564 (
            .O(N__16867),
            .I(N__16836));
    LocalMux I__3563 (
            .O(N__16864),
            .I(N__16833));
    Span4Mux_v I__3562 (
            .O(N__16861),
            .I(N__16828));
    LocalMux I__3561 (
            .O(N__16856),
            .I(N__16828));
    LocalMux I__3560 (
            .O(N__16851),
            .I(N__16825));
    LocalMux I__3559 (
            .O(N__16844),
            .I(N__16822));
    InMux I__3558 (
            .O(N__16843),
            .I(N__16819));
    InMux I__3557 (
            .O(N__16842),
            .I(N__16816));
    LocalMux I__3556 (
            .O(N__16839),
            .I(N__16813));
    LocalMux I__3555 (
            .O(N__16836),
            .I(N__16810));
    Span4Mux_v I__3554 (
            .O(N__16833),
            .I(N__16800));
    Span4Mux_v I__3553 (
            .O(N__16828),
            .I(N__16800));
    Span4Mux_v I__3552 (
            .O(N__16825),
            .I(N__16800));
    Sp12to4 I__3551 (
            .O(N__16822),
            .I(N__16795));
    LocalMux I__3550 (
            .O(N__16819),
            .I(N__16795));
    LocalMux I__3549 (
            .O(N__16816),
            .I(N__16788));
    Span4Mux_h I__3548 (
            .O(N__16813),
            .I(N__16788));
    Span4Mux_v I__3547 (
            .O(N__16810),
            .I(N__16788));
    InMux I__3546 (
            .O(N__16809),
            .I(N__16783));
    InMux I__3545 (
            .O(N__16808),
            .I(N__16783));
    InMux I__3544 (
            .O(N__16807),
            .I(N__16778));
    Span4Mux_h I__3543 (
            .O(N__16800),
            .I(N__16775));
    Span12Mux_s7_v I__3542 (
            .O(N__16795),
            .I(N__16768));
    Sp12to4 I__3541 (
            .O(N__16788),
            .I(N__16768));
    LocalMux I__3540 (
            .O(N__16783),
            .I(N__16768));
    InMux I__3539 (
            .O(N__16782),
            .I(N__16763));
    InMux I__3538 (
            .O(N__16781),
            .I(N__16763));
    LocalMux I__3537 (
            .O(N__16778),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    Odrv4 I__3536 (
            .O(N__16775),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    Odrv12 I__3535 (
            .O(N__16768),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    LocalMux I__3534 (
            .O(N__16763),
            .I(\c0.byte_transmit_counterZ0Z_1 ));
    InMux I__3533 (
            .O(N__16754),
            .I(N__16751));
    LocalMux I__3532 (
            .O(N__16751),
            .I(N__16748));
    Odrv4 I__3531 (
            .O(N__16748),
            .I(\c0.data_in_frame_6_Z0Z_0 ));
    InMux I__3530 (
            .O(N__16745),
            .I(N__16742));
    LocalMux I__3529 (
            .O(N__16742),
            .I(N__16738));
    CascadeMux I__3528 (
            .O(N__16741),
            .I(N__16734));
    Span4Mux_v I__3527 (
            .O(N__16738),
            .I(N__16731));
    InMux I__3526 (
            .O(N__16737),
            .I(N__16726));
    InMux I__3525 (
            .O(N__16734),
            .I(N__16726));
    Odrv4 I__3524 (
            .O(N__16731),
            .I(\c0.data_in_3_Z0Z_2 ));
    LocalMux I__3523 (
            .O(N__16726),
            .I(\c0.data_in_3_Z0Z_2 ));
    InMux I__3522 (
            .O(N__16721),
            .I(N__16718));
    LocalMux I__3521 (
            .O(N__16718),
            .I(N__16712));
    InMux I__3520 (
            .O(N__16717),
            .I(N__16709));
    InMux I__3519 (
            .O(N__16716),
            .I(N__16703));
    InMux I__3518 (
            .O(N__16715),
            .I(N__16703));
    Span4Mux_v I__3517 (
            .O(N__16712),
            .I(N__16698));
    LocalMux I__3516 (
            .O(N__16709),
            .I(N__16698));
    InMux I__3515 (
            .O(N__16708),
            .I(N__16695));
    LocalMux I__3514 (
            .O(N__16703),
            .I(N__16692));
    Span4Mux_h I__3513 (
            .O(N__16698),
            .I(N__16688));
    LocalMux I__3512 (
            .O(N__16695),
            .I(N__16685));
    Span4Mux_h I__3511 (
            .O(N__16692),
            .I(N__16682));
    InMux I__3510 (
            .O(N__16691),
            .I(N__16679));
    Odrv4 I__3509 (
            .O(N__16688),
            .I(\c0.d_4_26 ));
    Odrv12 I__3508 (
            .O(N__16685),
            .I(\c0.d_4_26 ));
    Odrv4 I__3507 (
            .O(N__16682),
            .I(\c0.d_4_26 ));
    LocalMux I__3506 (
            .O(N__16679),
            .I(\c0.d_4_26 ));
    InMux I__3505 (
            .O(N__16670),
            .I(N__16667));
    LocalMux I__3504 (
            .O(N__16667),
            .I(N__16664));
    Span4Mux_h I__3503 (
            .O(N__16664),
            .I(N__16661));
    Span4Mux_h I__3502 (
            .O(N__16661),
            .I(N__16658));
    Odrv4 I__3501 (
            .O(N__16658),
            .I(\c0.data_in_frame_6_Z0Z_1 ));
    InMux I__3500 (
            .O(N__16655),
            .I(N__16652));
    LocalMux I__3499 (
            .O(N__16652),
            .I(N__16649));
    Span4Mux_h I__3498 (
            .O(N__16649),
            .I(N__16646));
    Span4Mux_h I__3497 (
            .O(N__16646),
            .I(N__16641));
    InMux I__3496 (
            .O(N__16645),
            .I(N__16638));
    InMux I__3495 (
            .O(N__16644),
            .I(N__16635));
    Odrv4 I__3494 (
            .O(N__16641),
            .I(\c0.data_in_1_Z0Z_2 ));
    LocalMux I__3493 (
            .O(N__16638),
            .I(\c0.data_in_1_Z0Z_2 ));
    LocalMux I__3492 (
            .O(N__16635),
            .I(\c0.data_in_1_Z0Z_2 ));
    InMux I__3491 (
            .O(N__16628),
            .I(N__16624));
    CascadeMux I__3490 (
            .O(N__16627),
            .I(N__16621));
    LocalMux I__3489 (
            .O(N__16624),
            .I(N__16616));
    InMux I__3488 (
            .O(N__16621),
            .I(N__16612));
    InMux I__3487 (
            .O(N__16620),
            .I(N__16607));
    InMux I__3486 (
            .O(N__16619),
            .I(N__16607));
    Span4Mux_v I__3485 (
            .O(N__16616),
            .I(N__16604));
    InMux I__3484 (
            .O(N__16615),
            .I(N__16601));
    LocalMux I__3483 (
            .O(N__16612),
            .I(N__16598));
    LocalMux I__3482 (
            .O(N__16607),
            .I(N__16595));
    Span4Mux_h I__3481 (
            .O(N__16604),
            .I(N__16588));
    LocalMux I__3480 (
            .O(N__16601),
            .I(N__16588));
    Span4Mux_h I__3479 (
            .O(N__16598),
            .I(N__16588));
    Odrv12 I__3478 (
            .O(N__16595),
            .I(\c0.d_4_10 ));
    Odrv4 I__3477 (
            .O(N__16588),
            .I(\c0.d_4_10 ));
    CascadeMux I__3476 (
            .O(N__16583),
            .I(N__16580));
    InMux I__3475 (
            .O(N__16580),
            .I(N__16577));
    LocalMux I__3474 (
            .O(N__16577),
            .I(N__16574));
    Span4Mux_h I__3473 (
            .O(N__16574),
            .I(N__16571));
    Odrv4 I__3472 (
            .O(N__16571),
            .I(\c0.data_in_frame_7_Z0Z_0 ));
    InMux I__3471 (
            .O(N__16568),
            .I(N__16563));
    InMux I__3470 (
            .O(N__16567),
            .I(N__16560));
    InMux I__3469 (
            .O(N__16566),
            .I(N__16557));
    LocalMux I__3468 (
            .O(N__16563),
            .I(N__16554));
    LocalMux I__3467 (
            .O(N__16560),
            .I(N__16551));
    LocalMux I__3466 (
            .O(N__16557),
            .I(N__16548));
    Span4Mux_v I__3465 (
            .O(N__16554),
            .I(N__16545));
    Sp12to4 I__3464 (
            .O(N__16551),
            .I(N__16542));
    Span4Mux_h I__3463 (
            .O(N__16548),
            .I(N__16538));
    Sp12to4 I__3462 (
            .O(N__16545),
            .I(N__16533));
    Span12Mux_v I__3461 (
            .O(N__16542),
            .I(N__16533));
    InMux I__3460 (
            .O(N__16541),
            .I(N__16530));
    Odrv4 I__3459 (
            .O(N__16538),
            .I(\c0.d_2_36 ));
    Odrv12 I__3458 (
            .O(N__16533),
            .I(\c0.d_2_36 ));
    LocalMux I__3457 (
            .O(N__16530),
            .I(\c0.d_2_36 ));
    InMux I__3456 (
            .O(N__16523),
            .I(N__16520));
    LocalMux I__3455 (
            .O(N__16520),
            .I(N__16517));
    Span4Mux_v I__3454 (
            .O(N__16517),
            .I(N__16512));
    InMux I__3453 (
            .O(N__16516),
            .I(N__16509));
    InMux I__3452 (
            .O(N__16515),
            .I(N__16506));
    Span4Mux_h I__3451 (
            .O(N__16512),
            .I(N__16501));
    LocalMux I__3450 (
            .O(N__16509),
            .I(N__16501));
    LocalMux I__3449 (
            .O(N__16506),
            .I(N__16498));
    Span4Mux_h I__3448 (
            .O(N__16501),
            .I(N__16495));
    Span4Mux_h I__3447 (
            .O(N__16498),
            .I(N__16491));
    Span4Mux_v I__3446 (
            .O(N__16495),
            .I(N__16488));
    InMux I__3445 (
            .O(N__16494),
            .I(N__16485));
    Odrv4 I__3444 (
            .O(N__16491),
            .I(\c0.d_2_35 ));
    Odrv4 I__3443 (
            .O(N__16488),
            .I(\c0.d_2_35 ));
    LocalMux I__3442 (
            .O(N__16485),
            .I(\c0.d_2_35 ));
    CascadeMux I__3441 (
            .O(N__16478),
            .I(N__16475));
    InMux I__3440 (
            .O(N__16475),
            .I(N__16472));
    LocalMux I__3439 (
            .O(N__16472),
            .I(N__16469));
    Span4Mux_h I__3438 (
            .O(N__16469),
            .I(N__16466));
    Odrv4 I__3437 (
            .O(N__16466),
            .I(\c0.N_71 ));
    CascadeMux I__3436 (
            .O(N__16463),
            .I(N__16458));
    InMux I__3435 (
            .O(N__16462),
            .I(N__16454));
    InMux I__3434 (
            .O(N__16461),
            .I(N__16451));
    InMux I__3433 (
            .O(N__16458),
            .I(N__16446));
    InMux I__3432 (
            .O(N__16457),
            .I(N__16446));
    LocalMux I__3431 (
            .O(N__16454),
            .I(\c0.tx2.r_Bit_IndexZ0Z_0 ));
    LocalMux I__3430 (
            .O(N__16451),
            .I(\c0.tx2.r_Bit_IndexZ0Z_0 ));
    LocalMux I__3429 (
            .O(N__16446),
            .I(\c0.tx2.r_Bit_IndexZ0Z_0 ));
    InMux I__3428 (
            .O(N__16439),
            .I(N__16429));
    InMux I__3427 (
            .O(N__16438),
            .I(N__16424));
    InMux I__3426 (
            .O(N__16437),
            .I(N__16424));
    InMux I__3425 (
            .O(N__16436),
            .I(N__16415));
    InMux I__3424 (
            .O(N__16435),
            .I(N__16415));
    InMux I__3423 (
            .O(N__16434),
            .I(N__16408));
    InMux I__3422 (
            .O(N__16433),
            .I(N__16408));
    InMux I__3421 (
            .O(N__16432),
            .I(N__16408));
    LocalMux I__3420 (
            .O(N__16429),
            .I(N__16403));
    LocalMux I__3419 (
            .O(N__16424),
            .I(N__16403));
    InMux I__3418 (
            .O(N__16423),
            .I(N__16400));
    InMux I__3417 (
            .O(N__16422),
            .I(N__16393));
    InMux I__3416 (
            .O(N__16421),
            .I(N__16393));
    InMux I__3415 (
            .O(N__16420),
            .I(N__16393));
    LocalMux I__3414 (
            .O(N__16415),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    LocalMux I__3413 (
            .O(N__16408),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    Odrv4 I__3412 (
            .O(N__16403),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    LocalMux I__3411 (
            .O(N__16400),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    LocalMux I__3410 (
            .O(N__16393),
            .I(\c0.tx2.r_Clock_Count12_THRU_CO ));
    InMux I__3409 (
            .O(N__16382),
            .I(N__16378));
    InMux I__3408 (
            .O(N__16381),
            .I(N__16375));
    LocalMux I__3407 (
            .O(N__16378),
            .I(\c0.tx2.N_257 ));
    LocalMux I__3406 (
            .O(N__16375),
            .I(\c0.tx2.N_257 ));
    CascadeMux I__3405 (
            .O(N__16370),
            .I(\c0.tx2.N_258_cascade_ ));
    InMux I__3404 (
            .O(N__16367),
            .I(N__16362));
    InMux I__3403 (
            .O(N__16366),
            .I(N__16359));
    InMux I__3402 (
            .O(N__16365),
            .I(N__16356));
    LocalMux I__3401 (
            .O(N__16362),
            .I(N__16353));
    LocalMux I__3400 (
            .O(N__16359),
            .I(N__16341));
    LocalMux I__3399 (
            .O(N__16356),
            .I(N__16341));
    Span4Mux_h I__3398 (
            .O(N__16353),
            .I(N__16338));
    InMux I__3397 (
            .O(N__16352),
            .I(N__16331));
    InMux I__3396 (
            .O(N__16351),
            .I(N__16331));
    InMux I__3395 (
            .O(N__16350),
            .I(N__16331));
    InMux I__3394 (
            .O(N__16349),
            .I(N__16326));
    InMux I__3393 (
            .O(N__16348),
            .I(N__16326));
    InMux I__3392 (
            .O(N__16347),
            .I(N__16321));
    InMux I__3391 (
            .O(N__16346),
            .I(N__16321));
    Span4Mux_h I__3390 (
            .O(N__16341),
            .I(N__16318));
    Odrv4 I__3389 (
            .O(N__16338),
            .I(\c0.tx2.r_SM_MainZ0Z_1 ));
    LocalMux I__3388 (
            .O(N__16331),
            .I(\c0.tx2.r_SM_MainZ0Z_1 ));
    LocalMux I__3387 (
            .O(N__16326),
            .I(\c0.tx2.r_SM_MainZ0Z_1 ));
    LocalMux I__3386 (
            .O(N__16321),
            .I(\c0.tx2.r_SM_MainZ0Z_1 ));
    Odrv4 I__3385 (
            .O(N__16318),
            .I(\c0.tx2.r_SM_MainZ0Z_1 ));
    InMux I__3384 (
            .O(N__16307),
            .I(N__16293));
    InMux I__3383 (
            .O(N__16306),
            .I(N__16293));
    InMux I__3382 (
            .O(N__16305),
            .I(N__16293));
    InMux I__3381 (
            .O(N__16304),
            .I(N__16293));
    InMux I__3380 (
            .O(N__16303),
            .I(N__16290));
    InMux I__3379 (
            .O(N__16302),
            .I(N__16287));
    LocalMux I__3378 (
            .O(N__16293),
            .I(N__16284));
    LocalMux I__3377 (
            .O(N__16290),
            .I(\c0.tx2.r_Bit_IndexZ0Z_1 ));
    LocalMux I__3376 (
            .O(N__16287),
            .I(\c0.tx2.r_Bit_IndexZ0Z_1 ));
    Odrv4 I__3375 (
            .O(N__16284),
            .I(\c0.tx2.r_Bit_IndexZ0Z_1 ));
    CascadeMux I__3374 (
            .O(N__16277),
            .I(N__16274));
    InMux I__3373 (
            .O(N__16274),
            .I(N__16271));
    LocalMux I__3372 (
            .O(N__16271),
            .I(\c0.un1_data_in_7__7_0_a2_0_a2_2 ));
    InMux I__3371 (
            .O(N__16268),
            .I(N__16265));
    LocalMux I__3370 (
            .O(N__16265),
            .I(N__16262));
    Span4Mux_h I__3369 (
            .O(N__16262),
            .I(N__16259));
    Span4Mux_h I__3368 (
            .O(N__16259),
            .I(N__16255));
    InMux I__3367 (
            .O(N__16258),
            .I(N__16252));
    Odrv4 I__3366 (
            .O(N__16255),
            .I(\c0.data_in_0_Z0Z_5 ));
    LocalMux I__3365 (
            .O(N__16252),
            .I(\c0.data_in_0_Z0Z_5 ));
    InMux I__3364 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__3363 (
            .O(N__16244),
            .I(N__16241));
    Span4Mux_h I__3362 (
            .O(N__16241),
            .I(N__16238));
    Odrv4 I__3361 (
            .O(N__16238),
            .I(\c0.wait_for_transmission_RNOZ0Z_9 ));
    InMux I__3360 (
            .O(N__16235),
            .I(N__16232));
    LocalMux I__3359 (
            .O(N__16232),
            .I(N__16228));
    CascadeMux I__3358 (
            .O(N__16231),
            .I(N__16224));
    Span4Mux_h I__3357 (
            .O(N__16228),
            .I(N__16221));
    InMux I__3356 (
            .O(N__16227),
            .I(N__16218));
    InMux I__3355 (
            .O(N__16224),
            .I(N__16215));
    Odrv4 I__3354 (
            .O(N__16221),
            .I(\c0.data_in_2_Z0Z_2 ));
    LocalMux I__3353 (
            .O(N__16218),
            .I(\c0.data_in_2_Z0Z_2 ));
    LocalMux I__3352 (
            .O(N__16215),
            .I(\c0.data_in_2_Z0Z_2 ));
    InMux I__3351 (
            .O(N__16208),
            .I(N__16205));
    LocalMux I__3350 (
            .O(N__16205),
            .I(N__16202));
    Span4Mux_h I__3349 (
            .O(N__16202),
            .I(N__16198));
    CascadeMux I__3348 (
            .O(N__16201),
            .I(N__16194));
    Span4Mux_v I__3347 (
            .O(N__16198),
            .I(N__16191));
    InMux I__3346 (
            .O(N__16197),
            .I(N__16186));
    InMux I__3345 (
            .O(N__16194),
            .I(N__16186));
    Odrv4 I__3344 (
            .O(N__16191),
            .I(\c0.data_in_2_Z0Z_4 ));
    LocalMux I__3343 (
            .O(N__16186),
            .I(\c0.data_in_2_Z0Z_4 ));
    InMux I__3342 (
            .O(N__16181),
            .I(N__16177));
    InMux I__3341 (
            .O(N__16180),
            .I(N__16174));
    LocalMux I__3340 (
            .O(N__16177),
            .I(N__16171));
    LocalMux I__3339 (
            .O(N__16174),
            .I(N__16168));
    Span4Mux_h I__3338 (
            .O(N__16171),
            .I(N__16161));
    Span4Mux_v I__3337 (
            .O(N__16168),
            .I(N__16161));
    InMux I__3336 (
            .O(N__16167),
            .I(N__16156));
    InMux I__3335 (
            .O(N__16166),
            .I(N__16156));
    Odrv4 I__3334 (
            .O(N__16161),
            .I(\c0.d_4_18 ));
    LocalMux I__3333 (
            .O(N__16156),
            .I(\c0.d_4_18 ));
    InMux I__3332 (
            .O(N__16151),
            .I(N__16147));
    InMux I__3331 (
            .O(N__16150),
            .I(N__16144));
    LocalMux I__3330 (
            .O(N__16147),
            .I(N__16139));
    LocalMux I__3329 (
            .O(N__16144),
            .I(N__16139));
    Odrv12 I__3328 (
            .O(N__16139),
            .I(\c0.N_124 ));
    CascadeMux I__3327 (
            .O(N__16136),
            .I(\c0.N_124_cascade_ ));
    InMux I__3326 (
            .O(N__16133),
            .I(N__16129));
    InMux I__3325 (
            .O(N__16132),
            .I(N__16126));
    LocalMux I__3324 (
            .O(N__16129),
            .I(N__16121));
    LocalMux I__3323 (
            .O(N__16126),
            .I(N__16118));
    InMux I__3322 (
            .O(N__16125),
            .I(N__16115));
    InMux I__3321 (
            .O(N__16124),
            .I(N__16112));
    Odrv4 I__3320 (
            .O(N__16121),
            .I(\c0.d_4_RNI21N6Z0Z_11 ));
    Odrv4 I__3319 (
            .O(N__16118),
            .I(\c0.d_4_RNI21N6Z0Z_11 ));
    LocalMux I__3318 (
            .O(N__16115),
            .I(\c0.d_4_RNI21N6Z0Z_11 ));
    LocalMux I__3317 (
            .O(N__16112),
            .I(\c0.d_4_RNI21N6Z0Z_11 ));
    InMux I__3316 (
            .O(N__16103),
            .I(N__16100));
    LocalMux I__3315 (
            .O(N__16100),
            .I(N__16096));
    InMux I__3314 (
            .O(N__16099),
            .I(N__16093));
    Span4Mux_h I__3313 (
            .O(N__16096),
            .I(N__16090));
    LocalMux I__3312 (
            .O(N__16093),
            .I(\c0.d_4_RNIPF9J2Z0Z_37 ));
    Odrv4 I__3311 (
            .O(N__16090),
            .I(\c0.d_4_RNIPF9J2Z0Z_37 ));
    InMux I__3310 (
            .O(N__16085),
            .I(N__16082));
    LocalMux I__3309 (
            .O(N__16082),
            .I(N__16079));
    Span4Mux_v I__3308 (
            .O(N__16079),
            .I(N__16075));
    InMux I__3307 (
            .O(N__16078),
            .I(N__16072));
    Odrv4 I__3306 (
            .O(N__16075),
            .I(\c0.data_in_4_Z0Z_1 ));
    LocalMux I__3305 (
            .O(N__16072),
            .I(\c0.data_in_4_Z0Z_1 ));
    CascadeMux I__3304 (
            .O(N__16067),
            .I(N__16064));
    InMux I__3303 (
            .O(N__16064),
            .I(N__16060));
    InMux I__3302 (
            .O(N__16063),
            .I(N__16057));
    LocalMux I__3301 (
            .O(N__16060),
            .I(N__16054));
    LocalMux I__3300 (
            .O(N__16057),
            .I(N__16051));
    Span4Mux_h I__3299 (
            .O(N__16054),
            .I(N__16044));
    Span4Mux_h I__3298 (
            .O(N__16051),
            .I(N__16044));
    InMux I__3297 (
            .O(N__16050),
            .I(N__16039));
    InMux I__3296 (
            .O(N__16049),
            .I(N__16039));
    Odrv4 I__3295 (
            .O(N__16044),
            .I(\c0.d_4_33 ));
    LocalMux I__3294 (
            .O(N__16039),
            .I(\c0.d_4_33 ));
    CascadeMux I__3293 (
            .O(N__16034),
            .I(\c0.un1_data_in_6__3_0_a2_5_a2_2_cascade_ ));
    InMux I__3292 (
            .O(N__16031),
            .I(N__16026));
    InMux I__3291 (
            .O(N__16030),
            .I(N__16022));
    InMux I__3290 (
            .O(N__16029),
            .I(N__16019));
    LocalMux I__3289 (
            .O(N__16026),
            .I(N__16015));
    InMux I__3288 (
            .O(N__16025),
            .I(N__16012));
    LocalMux I__3287 (
            .O(N__16022),
            .I(N__16007));
    LocalMux I__3286 (
            .O(N__16019),
            .I(N__16007));
    InMux I__3285 (
            .O(N__16018),
            .I(N__16004));
    Odrv4 I__3284 (
            .O(N__16015),
            .I(\c0.d_4_25 ));
    LocalMux I__3283 (
            .O(N__16012),
            .I(\c0.d_4_25 ));
    Odrv4 I__3282 (
            .O(N__16007),
            .I(\c0.d_4_25 ));
    LocalMux I__3281 (
            .O(N__16004),
            .I(\c0.d_4_25 ));
    InMux I__3280 (
            .O(N__15995),
            .I(N__15992));
    LocalMux I__3279 (
            .O(N__15992),
            .I(N__15989));
    Span4Mux_v I__3278 (
            .O(N__15989),
            .I(N__15986));
    Odrv4 I__3277 (
            .O(N__15986),
            .I(\c0.un1_data_in_6__3 ));
    InMux I__3276 (
            .O(N__15983),
            .I(N__15980));
    LocalMux I__3275 (
            .O(N__15980),
            .I(\c0.un1_data_in_6__3_0_a2_5_a2_1 ));
    InMux I__3274 (
            .O(N__15977),
            .I(N__15973));
    InMux I__3273 (
            .O(N__15976),
            .I(N__15970));
    LocalMux I__3272 (
            .O(N__15973),
            .I(N__15967));
    LocalMux I__3271 (
            .O(N__15970),
            .I(N__15964));
    Span4Mux_h I__3270 (
            .O(N__15967),
            .I(N__15961));
    Span4Mux_h I__3269 (
            .O(N__15964),
            .I(N__15955));
    Span4Mux_h I__3268 (
            .O(N__15961),
            .I(N__15955));
    InMux I__3267 (
            .O(N__15960),
            .I(N__15952));
    Odrv4 I__3266 (
            .O(N__15955),
            .I(\c0.data_in_1_Z0Z_1 ));
    LocalMux I__3265 (
            .O(N__15952),
            .I(\c0.data_in_1_Z0Z_1 ));
    InMux I__3264 (
            .O(N__15947),
            .I(N__15943));
    InMux I__3263 (
            .O(N__15946),
            .I(N__15940));
    LocalMux I__3262 (
            .O(N__15943),
            .I(N__15936));
    LocalMux I__3261 (
            .O(N__15940),
            .I(N__15933));
    InMux I__3260 (
            .O(N__15939),
            .I(N__15930));
    Span12Mux_v I__3259 (
            .O(N__15936),
            .I(N__15927));
    Span4Mux_h I__3258 (
            .O(N__15933),
            .I(N__15922));
    LocalMux I__3257 (
            .O(N__15930),
            .I(N__15922));
    Odrv12 I__3256 (
            .O(N__15927),
            .I(\c0.data_in_2_Z0Z_7 ));
    Odrv4 I__3255 (
            .O(N__15922),
            .I(\c0.data_in_2_Z0Z_7 ));
    InMux I__3254 (
            .O(N__15917),
            .I(N__15914));
    LocalMux I__3253 (
            .O(N__15914),
            .I(N__15910));
    InMux I__3252 (
            .O(N__15913),
            .I(N__15907));
    Odrv12 I__3251 (
            .O(N__15910),
            .I(\c0.data_in_5_Z0Z_0 ));
    LocalMux I__3250 (
            .O(N__15907),
            .I(\c0.data_in_5_Z0Z_0 ));
    InMux I__3249 (
            .O(N__15902),
            .I(N__15899));
    LocalMux I__3248 (
            .O(N__15899),
            .I(N__15895));
    CascadeMux I__3247 (
            .O(N__15898),
            .I(N__15892));
    Span4Mux_h I__3246 (
            .O(N__15895),
            .I(N__15887));
    InMux I__3245 (
            .O(N__15892),
            .I(N__15884));
    InMux I__3244 (
            .O(N__15891),
            .I(N__15881));
    InMux I__3243 (
            .O(N__15890),
            .I(N__15878));
    Odrv4 I__3242 (
            .O(N__15887),
            .I(\c0.d_4_40 ));
    LocalMux I__3241 (
            .O(N__15884),
            .I(\c0.d_4_40 ));
    LocalMux I__3240 (
            .O(N__15881),
            .I(\c0.d_4_40 ));
    LocalMux I__3239 (
            .O(N__15878),
            .I(\c0.d_4_40 ));
    InMux I__3238 (
            .O(N__15869),
            .I(N__15866));
    LocalMux I__3237 (
            .O(N__15866),
            .I(N__15863));
    Span4Mux_h I__3236 (
            .O(N__15863),
            .I(N__15859));
    InMux I__3235 (
            .O(N__15862),
            .I(N__15856));
    Odrv4 I__3234 (
            .O(N__15859),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_4_1_0 ));
    LocalMux I__3233 (
            .O(N__15856),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_4_1_0 ));
    InMux I__3232 (
            .O(N__15851),
            .I(N__15848));
    LocalMux I__3231 (
            .O(N__15848),
            .I(N__15845));
    Span4Mux_h I__3230 (
            .O(N__15845),
            .I(N__15841));
    InMux I__3229 (
            .O(N__15844),
            .I(N__15838));
    Odrv4 I__3228 (
            .O(N__15841),
            .I(\c0.data_in_4_Z0Z_3 ));
    LocalMux I__3227 (
            .O(N__15838),
            .I(\c0.data_in_4_Z0Z_3 ));
    CascadeMux I__3226 (
            .O(N__15833),
            .I(\c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_ ));
    InMux I__3225 (
            .O(N__15830),
            .I(N__15827));
    LocalMux I__3224 (
            .O(N__15827),
            .I(N__15824));
    Odrv12 I__3223 (
            .O(N__15824),
            .I(\c0.g3_2 ));
    CascadeMux I__3222 (
            .O(N__15821),
            .I(\c0.un1_data_in_6__6_0_a2_0_a2_3_cascade_ ));
    InMux I__3221 (
            .O(N__15818),
            .I(N__15815));
    LocalMux I__3220 (
            .O(N__15815),
            .I(N__15812));
    Span4Mux_h I__3219 (
            .O(N__15812),
            .I(N__15804));
    InMux I__3218 (
            .O(N__15811),
            .I(N__15801));
    InMux I__3217 (
            .O(N__15810),
            .I(N__15798));
    InMux I__3216 (
            .O(N__15809),
            .I(N__15791));
    InMux I__3215 (
            .O(N__15808),
            .I(N__15791));
    InMux I__3214 (
            .O(N__15807),
            .I(N__15791));
    Odrv4 I__3213 (
            .O(N__15804),
            .I(\c0.N_128 ));
    LocalMux I__3212 (
            .O(N__15801),
            .I(\c0.N_128 ));
    LocalMux I__3211 (
            .O(N__15798),
            .I(\c0.N_128 ));
    LocalMux I__3210 (
            .O(N__15791),
            .I(\c0.N_128 ));
    InMux I__3209 (
            .O(N__15782),
            .I(N__15777));
    InMux I__3208 (
            .O(N__15781),
            .I(N__15774));
    CascadeMux I__3207 (
            .O(N__15780),
            .I(N__15771));
    LocalMux I__3206 (
            .O(N__15777),
            .I(N__15768));
    LocalMux I__3205 (
            .O(N__15774),
            .I(N__15765));
    InMux I__3204 (
            .O(N__15771),
            .I(N__15762));
    Span4Mux_h I__3203 (
            .O(N__15768),
            .I(N__15757));
    Span4Mux_h I__3202 (
            .O(N__15765),
            .I(N__15752));
    LocalMux I__3201 (
            .O(N__15762),
            .I(N__15752));
    InMux I__3200 (
            .O(N__15761),
            .I(N__15749));
    InMux I__3199 (
            .O(N__15760),
            .I(N__15746));
    Odrv4 I__3198 (
            .O(N__15757),
            .I(\c0.d_4_41 ));
    Odrv4 I__3197 (
            .O(N__15752),
            .I(\c0.d_4_41 ));
    LocalMux I__3196 (
            .O(N__15749),
            .I(\c0.d_4_41 ));
    LocalMux I__3195 (
            .O(N__15746),
            .I(\c0.d_4_41 ));
    CascadeMux I__3194 (
            .O(N__15737),
            .I(\c0.un1_data_in_6__5_0_a2_5_a2_2_cascade_ ));
    InMux I__3193 (
            .O(N__15734),
            .I(N__15729));
    InMux I__3192 (
            .O(N__15733),
            .I(N__15724));
    InMux I__3191 (
            .O(N__15732),
            .I(N__15724));
    LocalMux I__3190 (
            .O(N__15729),
            .I(N__15720));
    LocalMux I__3189 (
            .O(N__15724),
            .I(N__15717));
    CascadeMux I__3188 (
            .O(N__15723),
            .I(N__15714));
    Span4Mux_v I__3187 (
            .O(N__15720),
            .I(N__15711));
    Span4Mux_v I__3186 (
            .O(N__15717),
            .I(N__15708));
    InMux I__3185 (
            .O(N__15714),
            .I(N__15705));
    Odrv4 I__3184 (
            .O(N__15711),
            .I(\c0.N_132 ));
    Odrv4 I__3183 (
            .O(N__15708),
            .I(\c0.N_132 ));
    LocalMux I__3182 (
            .O(N__15705),
            .I(\c0.N_132 ));
    InMux I__3181 (
            .O(N__15698),
            .I(N__15695));
    LocalMux I__3180 (
            .O(N__15695),
            .I(N__15691));
    InMux I__3179 (
            .O(N__15694),
            .I(N__15688));
    Odrv12 I__3178 (
            .O(N__15691),
            .I(\c0.un1_data_in_6__6_0_a2_0_a2_3 ));
    LocalMux I__3177 (
            .O(N__15688),
            .I(\c0.un1_data_in_6__6_0_a2_0_a2_3 ));
    CascadeMux I__3176 (
            .O(N__15683),
            .I(\c0.un1_data_in_6__5_cascade_ ));
    InMux I__3175 (
            .O(N__15680),
            .I(N__15677));
    LocalMux I__3174 (
            .O(N__15677),
            .I(N__15674));
    Odrv4 I__3173 (
            .O(N__15674),
            .I(\c0.g0_2_0 ));
    InMux I__3172 (
            .O(N__15671),
            .I(N__15666));
    InMux I__3171 (
            .O(N__15670),
            .I(N__15661));
    InMux I__3170 (
            .O(N__15669),
            .I(N__15661));
    LocalMux I__3169 (
            .O(N__15666),
            .I(N__15655));
    LocalMux I__3168 (
            .O(N__15661),
            .I(N__15655));
    InMux I__3167 (
            .O(N__15660),
            .I(N__15652));
    Span4Mux_h I__3166 (
            .O(N__15655),
            .I(N__15649));
    LocalMux I__3165 (
            .O(N__15652),
            .I(\c0.d_4_43 ));
    Odrv4 I__3164 (
            .O(N__15649),
            .I(\c0.d_4_43 ));
    InMux I__3163 (
            .O(N__15644),
            .I(N__15641));
    LocalMux I__3162 (
            .O(N__15641),
            .I(\c0.un1_data_in_7__0_0_a2_1_a2_2 ));
    InMux I__3161 (
            .O(N__15638),
            .I(N__15635));
    LocalMux I__3160 (
            .O(N__15635),
            .I(\c0.un1_data_in_6__4 ));
    CascadeMux I__3159 (
            .O(N__15632),
            .I(\c0.wait_for_transmission4_12_5_1_cascade_ ));
    InMux I__3158 (
            .O(N__15629),
            .I(N__15625));
    InMux I__3157 (
            .O(N__15628),
            .I(N__15622));
    LocalMux I__3156 (
            .O(N__15625),
            .I(N__15619));
    LocalMux I__3155 (
            .O(N__15622),
            .I(N__15613));
    Span4Mux_h I__3154 (
            .O(N__15619),
            .I(N__15613));
    InMux I__3153 (
            .O(N__15618),
            .I(N__15610));
    Odrv4 I__3152 (
            .O(N__15613),
            .I(\c0.N_108 ));
    LocalMux I__3151 (
            .O(N__15610),
            .I(\c0.N_108 ));
    InMux I__3150 (
            .O(N__15605),
            .I(N__15602));
    LocalMux I__3149 (
            .O(N__15602),
            .I(N__15598));
    InMux I__3148 (
            .O(N__15601),
            .I(N__15590));
    Span4Mux_h I__3147 (
            .O(N__15598),
            .I(N__15587));
    InMux I__3146 (
            .O(N__15597),
            .I(N__15580));
    InMux I__3145 (
            .O(N__15596),
            .I(N__15580));
    InMux I__3144 (
            .O(N__15595),
            .I(N__15580));
    InMux I__3143 (
            .O(N__15594),
            .I(N__15577));
    InMux I__3142 (
            .O(N__15593),
            .I(N__15574));
    LocalMux I__3141 (
            .O(N__15590),
            .I(\c0.d_4_32 ));
    Odrv4 I__3140 (
            .O(N__15587),
            .I(\c0.d_4_32 ));
    LocalMux I__3139 (
            .O(N__15580),
            .I(\c0.d_4_32 ));
    LocalMux I__3138 (
            .O(N__15577),
            .I(\c0.d_4_32 ));
    LocalMux I__3137 (
            .O(N__15574),
            .I(\c0.d_4_32 ));
    InMux I__3136 (
            .O(N__15563),
            .I(N__15560));
    LocalMux I__3135 (
            .O(N__15560),
            .I(\c0.un1_data_in_7__6_0_a2_5_a2_2 ));
    InMux I__3134 (
            .O(N__15557),
            .I(N__15554));
    LocalMux I__3133 (
            .O(N__15554),
            .I(\c0.wait_for_transmission_RNOZ0Z_11 ));
    InMux I__3132 (
            .O(N__15551),
            .I(N__15547));
    InMux I__3131 (
            .O(N__15550),
            .I(N__15544));
    LocalMux I__3130 (
            .O(N__15547),
            .I(N__15541));
    LocalMux I__3129 (
            .O(N__15544),
            .I(N__15538));
    Span4Mux_v I__3128 (
            .O(N__15541),
            .I(N__15533));
    Span4Mux_h I__3127 (
            .O(N__15538),
            .I(N__15533));
    Odrv4 I__3126 (
            .O(N__15533),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_4_1 ));
    CascadeMux I__3125 (
            .O(N__15530),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_4_1_cascade_ ));
    CascadeMux I__3124 (
            .O(N__15527),
            .I(N__15521));
    InMux I__3123 (
            .O(N__15526),
            .I(N__15518));
    CascadeMux I__3122 (
            .O(N__15525),
            .I(N__15515));
    InMux I__3121 (
            .O(N__15524),
            .I(N__15510));
    InMux I__3120 (
            .O(N__15521),
            .I(N__15510));
    LocalMux I__3119 (
            .O(N__15518),
            .I(N__15507));
    InMux I__3118 (
            .O(N__15515),
            .I(N__15504));
    LocalMux I__3117 (
            .O(N__15510),
            .I(\c0.d_4_47 ));
    Odrv4 I__3116 (
            .O(N__15507),
            .I(\c0.d_4_47 ));
    LocalMux I__3115 (
            .O(N__15504),
            .I(\c0.d_4_47 ));
    InMux I__3114 (
            .O(N__15497),
            .I(N__15494));
    LocalMux I__3113 (
            .O(N__15494),
            .I(N__15491));
    Span4Mux_h I__3112 (
            .O(N__15491),
            .I(N__15487));
    InMux I__3111 (
            .O(N__15490),
            .I(N__15484));
    Odrv4 I__3110 (
            .O(N__15487),
            .I(\c0.N_125 ));
    LocalMux I__3109 (
            .O(N__15484),
            .I(\c0.N_125 ));
    InMux I__3108 (
            .O(N__15479),
            .I(N__15476));
    LocalMux I__3107 (
            .O(N__15476),
            .I(N__15473));
    Span4Mux_h I__3106 (
            .O(N__15473),
            .I(N__15469));
    InMux I__3105 (
            .O(N__15472),
            .I(N__15466));
    Odrv4 I__3104 (
            .O(N__15469),
            .I(\c0.data_in_0_Z0Z_6 ));
    LocalMux I__3103 (
            .O(N__15466),
            .I(\c0.data_in_0_Z0Z_6 ));
    InMux I__3102 (
            .O(N__15461),
            .I(N__15457));
    InMux I__3101 (
            .O(N__15460),
            .I(N__15453));
    LocalMux I__3100 (
            .O(N__15457),
            .I(N__15449));
    InMux I__3099 (
            .O(N__15456),
            .I(N__15446));
    LocalMux I__3098 (
            .O(N__15453),
            .I(N__15443));
    InMux I__3097 (
            .O(N__15452),
            .I(N__15440));
    Odrv4 I__3096 (
            .O(N__15449),
            .I(\c0.d_4_6 ));
    LocalMux I__3095 (
            .O(N__15446),
            .I(\c0.d_4_6 ));
    Odrv4 I__3094 (
            .O(N__15443),
            .I(\c0.d_4_6 ));
    LocalMux I__3093 (
            .O(N__15440),
            .I(\c0.d_4_6 ));
    InMux I__3092 (
            .O(N__15431),
            .I(N__15428));
    LocalMux I__3091 (
            .O(N__15428),
            .I(N__15425));
    Span4Mux_h I__3090 (
            .O(N__15425),
            .I(N__15420));
    InMux I__3089 (
            .O(N__15424),
            .I(N__15417));
    InMux I__3088 (
            .O(N__15423),
            .I(N__15414));
    Odrv4 I__3087 (
            .O(N__15420),
            .I(\c0.data_in_2_Z0Z_3 ));
    LocalMux I__3086 (
            .O(N__15417),
            .I(\c0.data_in_2_Z0Z_3 ));
    LocalMux I__3085 (
            .O(N__15414),
            .I(\c0.data_in_2_Z0Z_3 ));
    CascadeMux I__3084 (
            .O(N__15407),
            .I(N__15403));
    InMux I__3083 (
            .O(N__15406),
            .I(N__15398));
    InMux I__3082 (
            .O(N__15403),
            .I(N__15391));
    InMux I__3081 (
            .O(N__15402),
            .I(N__15391));
    InMux I__3080 (
            .O(N__15401),
            .I(N__15391));
    LocalMux I__3079 (
            .O(N__15398),
            .I(N__15387));
    LocalMux I__3078 (
            .O(N__15391),
            .I(N__15384));
    InMux I__3077 (
            .O(N__15390),
            .I(N__15380));
    Span4Mux_h I__3076 (
            .O(N__15387),
            .I(N__15375));
    Span4Mux_v I__3075 (
            .O(N__15384),
            .I(N__15375));
    InMux I__3074 (
            .O(N__15383),
            .I(N__15372));
    LocalMux I__3073 (
            .O(N__15380),
            .I(\c0.d_4_19 ));
    Odrv4 I__3072 (
            .O(N__15375),
            .I(\c0.d_4_19 ));
    LocalMux I__3071 (
            .O(N__15372),
            .I(\c0.d_4_19 ));
    InMux I__3070 (
            .O(N__15365),
            .I(N__15362));
    LocalMux I__3069 (
            .O(N__15362),
            .I(N__15357));
    InMux I__3068 (
            .O(N__15361),
            .I(N__15354));
    InMux I__3067 (
            .O(N__15360),
            .I(N__15351));
    Span4Mux_v I__3066 (
            .O(N__15357),
            .I(N__15345));
    LocalMux I__3065 (
            .O(N__15354),
            .I(N__15345));
    LocalMux I__3064 (
            .O(N__15351),
            .I(N__15342));
    InMux I__3063 (
            .O(N__15350),
            .I(N__15339));
    Odrv4 I__3062 (
            .O(N__15345),
            .I(\c0.d_2_31 ));
    Odrv4 I__3061 (
            .O(N__15342),
            .I(\c0.d_2_31 ));
    LocalMux I__3060 (
            .O(N__15339),
            .I(\c0.d_2_31 ));
    InMux I__3059 (
            .O(N__15332),
            .I(N__15327));
    InMux I__3058 (
            .O(N__15331),
            .I(N__15324));
    CascadeMux I__3057 (
            .O(N__15330),
            .I(N__15321));
    LocalMux I__3056 (
            .O(N__15327),
            .I(N__15318));
    LocalMux I__3055 (
            .O(N__15324),
            .I(N__15315));
    InMux I__3054 (
            .O(N__15321),
            .I(N__15312));
    Span4Mux_v I__3053 (
            .O(N__15318),
            .I(N__15309));
    Span4Mux_v I__3052 (
            .O(N__15315),
            .I(N__15303));
    LocalMux I__3051 (
            .O(N__15312),
            .I(N__15303));
    Span4Mux_h I__3050 (
            .O(N__15309),
            .I(N__15300));
    InMux I__3049 (
            .O(N__15308),
            .I(N__15297));
    Span4Mux_h I__3048 (
            .O(N__15303),
            .I(N__15294));
    Odrv4 I__3047 (
            .O(N__15300),
            .I(\c0.d_2_43 ));
    LocalMux I__3046 (
            .O(N__15297),
            .I(\c0.d_2_43 ));
    Odrv4 I__3045 (
            .O(N__15294),
            .I(\c0.d_2_43 ));
    InMux I__3044 (
            .O(N__15287),
            .I(N__15283));
    InMux I__3043 (
            .O(N__15286),
            .I(N__15279));
    LocalMux I__3042 (
            .O(N__15283),
            .I(N__15276));
    InMux I__3041 (
            .O(N__15282),
            .I(N__15273));
    LocalMux I__3040 (
            .O(N__15279),
            .I(N__15270));
    Span4Mux_h I__3039 (
            .O(N__15276),
            .I(N__15265));
    LocalMux I__3038 (
            .O(N__15273),
            .I(N__15265));
    Span4Mux_v I__3037 (
            .O(N__15270),
            .I(N__15260));
    Span4Mux_h I__3036 (
            .O(N__15265),
            .I(N__15260));
    Odrv4 I__3035 (
            .O(N__15260),
            .I(\c0.d_2_15 ));
    CascadeMux I__3034 (
            .O(N__15257),
            .I(N__15254));
    InMux I__3033 (
            .O(N__15254),
            .I(N__15251));
    LocalMux I__3032 (
            .O(N__15251),
            .I(N__15248));
    Span4Mux_v I__3031 (
            .O(N__15248),
            .I(N__15243));
    InMux I__3030 (
            .O(N__15247),
            .I(N__15240));
    CascadeMux I__3029 (
            .O(N__15246),
            .I(N__15236));
    Span4Mux_h I__3028 (
            .O(N__15243),
            .I(N__15231));
    LocalMux I__3027 (
            .O(N__15240),
            .I(N__15231));
    InMux I__3026 (
            .O(N__15239),
            .I(N__15228));
    InMux I__3025 (
            .O(N__15236),
            .I(N__15225));
    Span4Mux_h I__3024 (
            .O(N__15231),
            .I(N__15222));
    LocalMux I__3023 (
            .O(N__15228),
            .I(N__15217));
    LocalMux I__3022 (
            .O(N__15225),
            .I(N__15217));
    Span4Mux_h I__3021 (
            .O(N__15222),
            .I(N__15214));
    Odrv12 I__3020 (
            .O(N__15217),
            .I(\c0.d_2_2 ));
    Odrv4 I__3019 (
            .O(N__15214),
            .I(\c0.d_2_2 ));
    InMux I__3018 (
            .O(N__15209),
            .I(N__15205));
    CascadeMux I__3017 (
            .O(N__15208),
            .I(N__15202));
    LocalMux I__3016 (
            .O(N__15205),
            .I(N__15199));
    InMux I__3015 (
            .O(N__15202),
            .I(N__15196));
    Span4Mux_v I__3014 (
            .O(N__15199),
            .I(N__15192));
    LocalMux I__3013 (
            .O(N__15196),
            .I(N__15189));
    InMux I__3012 (
            .O(N__15195),
            .I(N__15186));
    Odrv4 I__3011 (
            .O(N__15192),
            .I(\c0.d_2_47 ));
    Odrv4 I__3010 (
            .O(N__15189),
            .I(\c0.d_2_47 ));
    LocalMux I__3009 (
            .O(N__15186),
            .I(\c0.d_2_47 ));
    CascadeMux I__3008 (
            .O(N__15179),
            .I(\c0.un105_newcrc_0_a2_3_cascade_ ));
    InMux I__3007 (
            .O(N__15176),
            .I(N__15173));
    LocalMux I__3006 (
            .O(N__15173),
            .I(\c0.un105_newcrc_0_a2_4 ));
    InMux I__3005 (
            .O(N__15170),
            .I(N__15167));
    LocalMux I__3004 (
            .O(N__15167),
            .I(N__15163));
    InMux I__3003 (
            .O(N__15166),
            .I(N__15160));
    Span4Mux_v I__3002 (
            .O(N__15163),
            .I(N__15154));
    LocalMux I__3001 (
            .O(N__15160),
            .I(N__15154));
    InMux I__3000 (
            .O(N__15159),
            .I(N__15151));
    Span4Mux_h I__2999 (
            .O(N__15154),
            .I(N__15148));
    LocalMux I__2998 (
            .O(N__15151),
            .I(\c0.d_2_5 ));
    Odrv4 I__2997 (
            .O(N__15148),
            .I(\c0.d_2_5 ));
    InMux I__2996 (
            .O(N__15143),
            .I(N__15139));
    InMux I__2995 (
            .O(N__15142),
            .I(N__15136));
    LocalMux I__2994 (
            .O(N__15139),
            .I(N__15130));
    LocalMux I__2993 (
            .O(N__15136),
            .I(N__15130));
    InMux I__2992 (
            .O(N__15135),
            .I(N__15127));
    Span4Mux_v I__2991 (
            .O(N__15130),
            .I(N__15123));
    LocalMux I__2990 (
            .O(N__15127),
            .I(N__15120));
    InMux I__2989 (
            .O(N__15126),
            .I(N__15117));
    Odrv4 I__2988 (
            .O(N__15123),
            .I(\c0.d_2_32 ));
    Odrv12 I__2987 (
            .O(N__15120),
            .I(\c0.d_2_32 ));
    LocalMux I__2986 (
            .O(N__15117),
            .I(\c0.d_2_32 ));
    CascadeMux I__2985 (
            .O(N__15110),
            .I(N__15107));
    InMux I__2984 (
            .O(N__15107),
            .I(N__15102));
    InMux I__2983 (
            .O(N__15106),
            .I(N__15099));
    InMux I__2982 (
            .O(N__15105),
            .I(N__15095));
    LocalMux I__2981 (
            .O(N__15102),
            .I(N__15092));
    LocalMux I__2980 (
            .O(N__15099),
            .I(N__15089));
    InMux I__2979 (
            .O(N__15098),
            .I(N__15086));
    LocalMux I__2978 (
            .O(N__15095),
            .I(N__15083));
    Span4Mux_v I__2977 (
            .O(N__15092),
            .I(N__15080));
    Span4Mux_v I__2976 (
            .O(N__15089),
            .I(N__15073));
    LocalMux I__2975 (
            .O(N__15086),
            .I(N__15073));
    Span4Mux_v I__2974 (
            .O(N__15083),
            .I(N__15073));
    Span4Mux_h I__2973 (
            .O(N__15080),
            .I(N__15070));
    Span4Mux_h I__2972 (
            .O(N__15073),
            .I(N__15067));
    Odrv4 I__2971 (
            .O(N__15070),
            .I(\c0.d_2_18 ));
    Odrv4 I__2970 (
            .O(N__15067),
            .I(\c0.d_2_18 ));
    CascadeMux I__2969 (
            .O(N__15062),
            .I(N__15057));
    InMux I__2968 (
            .O(N__15061),
            .I(N__15052));
    InMux I__2967 (
            .O(N__15060),
            .I(N__15049));
    InMux I__2966 (
            .O(N__15057),
            .I(N__15046));
    InMux I__2965 (
            .O(N__15056),
            .I(N__15041));
    InMux I__2964 (
            .O(N__15055),
            .I(N__15041));
    LocalMux I__2963 (
            .O(N__15052),
            .I(N__15038));
    LocalMux I__2962 (
            .O(N__15049),
            .I(N__15035));
    LocalMux I__2961 (
            .O(N__15046),
            .I(N__15032));
    LocalMux I__2960 (
            .O(N__15041),
            .I(\c0.d_2_46 ));
    Odrv12 I__2959 (
            .O(N__15038),
            .I(\c0.d_2_46 ));
    Odrv12 I__2958 (
            .O(N__15035),
            .I(\c0.d_2_46 ));
    Odrv4 I__2957 (
            .O(N__15032),
            .I(\c0.d_2_46 ));
    InMux I__2956 (
            .O(N__15023),
            .I(N__15018));
    InMux I__2955 (
            .O(N__15022),
            .I(N__15014));
    InMux I__2954 (
            .O(N__15021),
            .I(N__15011));
    LocalMux I__2953 (
            .O(N__15018),
            .I(N__15008));
    CascadeMux I__2952 (
            .O(N__15017),
            .I(N__15005));
    LocalMux I__2951 (
            .O(N__15014),
            .I(N__15002));
    LocalMux I__2950 (
            .O(N__15011),
            .I(N__14999));
    Span4Mux_v I__2949 (
            .O(N__15008),
            .I(N__14996));
    InMux I__2948 (
            .O(N__15005),
            .I(N__14993));
    Span4Mux_v I__2947 (
            .O(N__15002),
            .I(N__14990));
    Span4Mux_h I__2946 (
            .O(N__14999),
            .I(N__14987));
    Odrv4 I__2945 (
            .O(N__14996),
            .I(\c0.d_2_20 ));
    LocalMux I__2944 (
            .O(N__14993),
            .I(\c0.d_2_20 ));
    Odrv4 I__2943 (
            .O(N__14990),
            .I(\c0.d_2_20 ));
    Odrv4 I__2942 (
            .O(N__14987),
            .I(\c0.d_2_20 ));
    InMux I__2941 (
            .O(N__14978),
            .I(N__14975));
    LocalMux I__2940 (
            .O(N__14975),
            .I(N__14971));
    InMux I__2939 (
            .O(N__14974),
            .I(N__14968));
    Span4Mux_v I__2938 (
            .O(N__14971),
            .I(N__14965));
    LocalMux I__2937 (
            .O(N__14968),
            .I(\c0.nextCRC16_3_3_1 ));
    Odrv4 I__2936 (
            .O(N__14965),
            .I(\c0.nextCRC16_3_3_1 ));
    InMux I__2935 (
            .O(N__14960),
            .I(N__14956));
    InMux I__2934 (
            .O(N__14959),
            .I(N__14953));
    LocalMux I__2933 (
            .O(N__14956),
            .I(N__14950));
    LocalMux I__2932 (
            .O(N__14953),
            .I(N__14947));
    Span4Mux_h I__2931 (
            .O(N__14950),
            .I(N__14944));
    Span4Mux_v I__2930 (
            .O(N__14947),
            .I(N__14941));
    Span4Mux_v I__2929 (
            .O(N__14944),
            .I(N__14934));
    Span4Mux_h I__2928 (
            .O(N__14941),
            .I(N__14934));
    InMux I__2927 (
            .O(N__14940),
            .I(N__14931));
    InMux I__2926 (
            .O(N__14939),
            .I(N__14928));
    Odrv4 I__2925 (
            .O(N__14934),
            .I(\c0.d_2_17 ));
    LocalMux I__2924 (
            .O(N__14931),
            .I(\c0.d_2_17 ));
    LocalMux I__2923 (
            .O(N__14928),
            .I(\c0.d_2_17 ));
    CascadeMux I__2922 (
            .O(N__14921),
            .I(N__14917));
    CascadeMux I__2921 (
            .O(N__14920),
            .I(N__14913));
    InMux I__2920 (
            .O(N__14917),
            .I(N__14909));
    InMux I__2919 (
            .O(N__14916),
            .I(N__14906));
    InMux I__2918 (
            .O(N__14913),
            .I(N__14903));
    CascadeMux I__2917 (
            .O(N__14912),
            .I(N__14900));
    LocalMux I__2916 (
            .O(N__14909),
            .I(N__14896));
    LocalMux I__2915 (
            .O(N__14906),
            .I(N__14893));
    LocalMux I__2914 (
            .O(N__14903),
            .I(N__14890));
    InMux I__2913 (
            .O(N__14900),
            .I(N__14886));
    InMux I__2912 (
            .O(N__14899),
            .I(N__14883));
    Span4Mux_h I__2911 (
            .O(N__14896),
            .I(N__14880));
    Span4Mux_v I__2910 (
            .O(N__14893),
            .I(N__14875));
    Span4Mux_v I__2909 (
            .O(N__14890),
            .I(N__14875));
    InMux I__2908 (
            .O(N__14889),
            .I(N__14872));
    LocalMux I__2907 (
            .O(N__14886),
            .I(\c0.d_2_1 ));
    LocalMux I__2906 (
            .O(N__14883),
            .I(\c0.d_2_1 ));
    Odrv4 I__2905 (
            .O(N__14880),
            .I(\c0.d_2_1 ));
    Odrv4 I__2904 (
            .O(N__14875),
            .I(\c0.d_2_1 ));
    LocalMux I__2903 (
            .O(N__14872),
            .I(\c0.d_2_1 ));
    InMux I__2902 (
            .O(N__14861),
            .I(N__14857));
    InMux I__2901 (
            .O(N__14860),
            .I(N__14853));
    LocalMux I__2900 (
            .O(N__14857),
            .I(N__14850));
    InMux I__2899 (
            .O(N__14856),
            .I(N__14847));
    LocalMux I__2898 (
            .O(N__14853),
            .I(N__14844));
    Span4Mux_v I__2897 (
            .O(N__14850),
            .I(N__14838));
    LocalMux I__2896 (
            .O(N__14847),
            .I(N__14838));
    Span4Mux_h I__2895 (
            .O(N__14844),
            .I(N__14835));
    InMux I__2894 (
            .O(N__14843),
            .I(N__14832));
    Odrv4 I__2893 (
            .O(N__14838),
            .I(\c0.d_2_4 ));
    Odrv4 I__2892 (
            .O(N__14835),
            .I(\c0.d_2_4 ));
    LocalMux I__2891 (
            .O(N__14832),
            .I(\c0.d_2_4 ));
    CascadeMux I__2890 (
            .O(N__14825),
            .I(N__14822));
    InMux I__2889 (
            .O(N__14822),
            .I(N__14819));
    LocalMux I__2888 (
            .O(N__14819),
            .I(\c0.nextCRC16_3_0_a2_1_1 ));
    CascadeMux I__2887 (
            .O(N__14816),
            .I(N__14813));
    InMux I__2886 (
            .O(N__14813),
            .I(N__14810));
    LocalMux I__2885 (
            .O(N__14810),
            .I(\c0.un1_data_in_6__4_0_a2_5_a2_1 ));
    InMux I__2884 (
            .O(N__14807),
            .I(N__14804));
    LocalMux I__2883 (
            .O(N__14804),
            .I(N__14800));
    InMux I__2882 (
            .O(N__14803),
            .I(N__14795));
    Span4Mux_v I__2881 (
            .O(N__14800),
            .I(N__14792));
    InMux I__2880 (
            .O(N__14799),
            .I(N__14787));
    InMux I__2879 (
            .O(N__14798),
            .I(N__14787));
    LocalMux I__2878 (
            .O(N__14795),
            .I(\c0.N_133 ));
    Odrv4 I__2877 (
            .O(N__14792),
            .I(\c0.N_133 ));
    LocalMux I__2876 (
            .O(N__14787),
            .I(\c0.N_133 ));
    CascadeMux I__2875 (
            .O(N__14780),
            .I(N__14777));
    InMux I__2874 (
            .O(N__14777),
            .I(N__14774));
    LocalMux I__2873 (
            .O(N__14774),
            .I(N__14771));
    Span4Mux_h I__2872 (
            .O(N__14771),
            .I(N__14768));
    Odrv4 I__2871 (
            .O(N__14768),
            .I(\c0.un1_data_in_7__2_0_a2_0_a2_5 ));
    InMux I__2870 (
            .O(N__14765),
            .I(N__14762));
    LocalMux I__2869 (
            .O(N__14762),
            .I(N__14759));
    Odrv4 I__2868 (
            .O(N__14759),
            .I(\c0.tx2_data_1_iv_4_6 ));
    CascadeMux I__2867 (
            .O(N__14756),
            .I(N__14753));
    InMux I__2866 (
            .O(N__14753),
            .I(N__14750));
    LocalMux I__2865 (
            .O(N__14750),
            .I(N__14747));
    Odrv4 I__2864 (
            .O(N__14747),
            .I(\c0.tx2_data_1_iv_3_6 ));
    CascadeMux I__2863 (
            .O(N__14744),
            .I(N__14741));
    InMux I__2862 (
            .O(N__14741),
            .I(N__14738));
    LocalMux I__2861 (
            .O(N__14738),
            .I(\c0.tx2.r_Tx_DataZ0Z_6 ));
    CascadeMux I__2860 (
            .O(N__14735),
            .I(N__14732));
    InMux I__2859 (
            .O(N__14732),
            .I(N__14728));
    CascadeMux I__2858 (
            .O(N__14731),
            .I(N__14725));
    LocalMux I__2857 (
            .O(N__14728),
            .I(N__14722));
    InMux I__2856 (
            .O(N__14725),
            .I(N__14719));
    Span4Mux_v I__2855 (
            .O(N__14722),
            .I(N__14714));
    LocalMux I__2854 (
            .O(N__14719),
            .I(N__14714));
    Span4Mux_h I__2853 (
            .O(N__14714),
            .I(N__14711));
    Span4Mux_h I__2852 (
            .O(N__14711),
            .I(N__14708));
    Odrv4 I__2851 (
            .O(N__14708),
            .I(\c0.d_2_27 ));
    InMux I__2850 (
            .O(N__14705),
            .I(N__14702));
    LocalMux I__2849 (
            .O(N__14702),
            .I(N__14699));
    Span4Mux_h I__2848 (
            .O(N__14699),
            .I(N__14696));
    Odrv4 I__2847 (
            .O(N__14696),
            .I(\c0.tx_data_RNO_1Z0Z_3 ));
    CascadeMux I__2846 (
            .O(N__14693),
            .I(N__14690));
    InMux I__2845 (
            .O(N__14690),
            .I(N__14687));
    LocalMux I__2844 (
            .O(N__14687),
            .I(N__14684));
    Odrv12 I__2843 (
            .O(N__14684),
            .I(\c0.data_out_7_Z0Z_7 ));
    CascadeMux I__2842 (
            .O(N__14681),
            .I(N__14678));
    InMux I__2841 (
            .O(N__14678),
            .I(N__14675));
    LocalMux I__2840 (
            .O(N__14675),
            .I(N__14672));
    Odrv12 I__2839 (
            .O(N__14672),
            .I(\c0.tx_data_RNO_1Z0Z_7 ));
    CascadeMux I__2838 (
            .O(N__14669),
            .I(\c0.tx_data_RNO_3Z0Z_2_cascade_ ));
    InMux I__2837 (
            .O(N__14666),
            .I(N__14663));
    LocalMux I__2836 (
            .O(N__14663),
            .I(N__14660));
    Odrv4 I__2835 (
            .O(N__14660),
            .I(\c0.tx_data_1_0_i_ns_1_2 ));
    InMux I__2834 (
            .O(N__14657),
            .I(N__14654));
    LocalMux I__2833 (
            .O(N__14654),
            .I(N__14650));
    InMux I__2832 (
            .O(N__14653),
            .I(N__14647));
    Span4Mux_h I__2831 (
            .O(N__14650),
            .I(N__14642));
    LocalMux I__2830 (
            .O(N__14647),
            .I(N__14642));
    Span4Mux_h I__2829 (
            .O(N__14642),
            .I(N__14638));
    InMux I__2828 (
            .O(N__14641),
            .I(N__14635));
    Odrv4 I__2827 (
            .O(N__14638),
            .I(\c0.d_2_10 ));
    LocalMux I__2826 (
            .O(N__14635),
            .I(\c0.d_2_10 ));
    CascadeMux I__2825 (
            .O(N__14630),
            .I(N__14625));
    CascadeMux I__2824 (
            .O(N__14629),
            .I(N__14622));
    CascadeMux I__2823 (
            .O(N__14628),
            .I(N__14619));
    InMux I__2822 (
            .O(N__14625),
            .I(N__14615));
    InMux I__2821 (
            .O(N__14622),
            .I(N__14610));
    InMux I__2820 (
            .O(N__14619),
            .I(N__14610));
    InMux I__2819 (
            .O(N__14618),
            .I(N__14607));
    LocalMux I__2818 (
            .O(N__14615),
            .I(N__14604));
    LocalMux I__2817 (
            .O(N__14610),
            .I(N__14600));
    LocalMux I__2816 (
            .O(N__14607),
            .I(N__14595));
    Span4Mux_v I__2815 (
            .O(N__14604),
            .I(N__14595));
    InMux I__2814 (
            .O(N__14603),
            .I(N__14592));
    Span4Mux_h I__2813 (
            .O(N__14600),
            .I(N__14589));
    Odrv4 I__2812 (
            .O(N__14595),
            .I(\c0.d_2_42 ));
    LocalMux I__2811 (
            .O(N__14592),
            .I(\c0.d_2_42 ));
    Odrv4 I__2810 (
            .O(N__14589),
            .I(\c0.d_2_42 ));
    InMux I__2809 (
            .O(N__14582),
            .I(N__14579));
    LocalMux I__2808 (
            .O(N__14579),
            .I(\c0.tx_data_RNO_4Z0Z_2 ));
    InMux I__2807 (
            .O(N__14576),
            .I(N__14573));
    LocalMux I__2806 (
            .O(N__14573),
            .I(N__14570));
    Span4Mux_h I__2805 (
            .O(N__14570),
            .I(N__14566));
    InMux I__2804 (
            .O(N__14569),
            .I(N__14563));
    Odrv4 I__2803 (
            .O(N__14566),
            .I(\c0.N_81 ));
    LocalMux I__2802 (
            .O(N__14563),
            .I(\c0.N_81 ));
    InMux I__2801 (
            .O(N__14558),
            .I(N__14554));
    InMux I__2800 (
            .O(N__14557),
            .I(N__14551));
    LocalMux I__2799 (
            .O(N__14554),
            .I(N__14547));
    LocalMux I__2798 (
            .O(N__14551),
            .I(N__14543));
    InMux I__2797 (
            .O(N__14550),
            .I(N__14540));
    Span4Mux_h I__2796 (
            .O(N__14547),
            .I(N__14537));
    InMux I__2795 (
            .O(N__14546),
            .I(N__14534));
    Span4Mux_h I__2794 (
            .O(N__14543),
            .I(N__14529));
    LocalMux I__2793 (
            .O(N__14540),
            .I(N__14529));
    Span4Mux_h I__2792 (
            .O(N__14537),
            .I(N__14526));
    LocalMux I__2791 (
            .O(N__14534),
            .I(\c0.d_2_29 ));
    Odrv4 I__2790 (
            .O(N__14529),
            .I(\c0.d_2_29 ));
    Odrv4 I__2789 (
            .O(N__14526),
            .I(\c0.d_2_29 ));
    CascadeMux I__2788 (
            .O(N__14519),
            .I(N__14515));
    CascadeMux I__2787 (
            .O(N__14518),
            .I(N__14512));
    InMux I__2786 (
            .O(N__14515),
            .I(N__14506));
    InMux I__2785 (
            .O(N__14512),
            .I(N__14506));
    InMux I__2784 (
            .O(N__14511),
            .I(N__14502));
    LocalMux I__2783 (
            .O(N__14506),
            .I(N__14497));
    CascadeMux I__2782 (
            .O(N__14505),
            .I(N__14494));
    LocalMux I__2781 (
            .O(N__14502),
            .I(N__14491));
    InMux I__2780 (
            .O(N__14501),
            .I(N__14488));
    InMux I__2779 (
            .O(N__14500),
            .I(N__14485));
    Span4Mux_h I__2778 (
            .O(N__14497),
            .I(N__14482));
    InMux I__2777 (
            .O(N__14494),
            .I(N__14479));
    Span4Mux_h I__2776 (
            .O(N__14491),
            .I(N__14474));
    LocalMux I__2775 (
            .O(N__14488),
            .I(N__14474));
    LocalMux I__2774 (
            .O(N__14485),
            .I(\c0.d_2_30 ));
    Odrv4 I__2773 (
            .O(N__14482),
            .I(\c0.d_2_30 ));
    LocalMux I__2772 (
            .O(N__14479),
            .I(\c0.d_2_30 ));
    Odrv4 I__2771 (
            .O(N__14474),
            .I(\c0.d_2_30 ));
    InMux I__2770 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__2769 (
            .O(N__14462),
            .I(N__14459));
    Odrv12 I__2768 (
            .O(N__14459),
            .I(\c0.data_out_7_Z0Z_3 ));
    CascadeMux I__2767 (
            .O(N__14456),
            .I(\c0.tx2_data_1_iv_4_1_6_cascade_ ));
    InMux I__2766 (
            .O(N__14453),
            .I(N__14450));
    LocalMux I__2765 (
            .O(N__14450),
            .I(N__14447));
    Span4Mux_h I__2764 (
            .O(N__14447),
            .I(N__14443));
    InMux I__2763 (
            .O(N__14446),
            .I(N__14440));
    Odrv4 I__2762 (
            .O(N__14443),
            .I(\c0.data_in_5_Z0Z_3 ));
    LocalMux I__2761 (
            .O(N__14440),
            .I(\c0.data_in_5_Z0Z_3 ));
    InMux I__2760 (
            .O(N__14435),
            .I(N__14422));
    InMux I__2759 (
            .O(N__14434),
            .I(N__14422));
    InMux I__2758 (
            .O(N__14433),
            .I(N__14422));
    CascadeMux I__2757 (
            .O(N__14432),
            .I(N__14416));
    CascadeMux I__2756 (
            .O(N__14431),
            .I(N__14413));
    CascadeMux I__2755 (
            .O(N__14430),
            .I(N__14410));
    CascadeMux I__2754 (
            .O(N__14429),
            .I(N__14405));
    LocalMux I__2753 (
            .O(N__14422),
            .I(N__14402));
    CascadeMux I__2752 (
            .O(N__14421),
            .I(N__14399));
    InMux I__2751 (
            .O(N__14420),
            .I(N__14391));
    InMux I__2750 (
            .O(N__14419),
            .I(N__14391));
    InMux I__2749 (
            .O(N__14416),
            .I(N__14391));
    InMux I__2748 (
            .O(N__14413),
            .I(N__14384));
    InMux I__2747 (
            .O(N__14410),
            .I(N__14384));
    InMux I__2746 (
            .O(N__14409),
            .I(N__14384));
    InMux I__2745 (
            .O(N__14408),
            .I(N__14379));
    InMux I__2744 (
            .O(N__14405),
            .I(N__14379));
    Span4Mux_h I__2743 (
            .O(N__14402),
            .I(N__14376));
    InMux I__2742 (
            .O(N__14399),
            .I(N__14373));
    InMux I__2741 (
            .O(N__14398),
            .I(N__14370));
    LocalMux I__2740 (
            .O(N__14391),
            .I(N__14367));
    LocalMux I__2739 (
            .O(N__14384),
            .I(\c0.tx2.r_SM_MainZ0Z_2 ));
    LocalMux I__2738 (
            .O(N__14379),
            .I(\c0.tx2.r_SM_MainZ0Z_2 ));
    Odrv4 I__2737 (
            .O(N__14376),
            .I(\c0.tx2.r_SM_MainZ0Z_2 ));
    LocalMux I__2736 (
            .O(N__14373),
            .I(\c0.tx2.r_SM_MainZ0Z_2 ));
    LocalMux I__2735 (
            .O(N__14370),
            .I(\c0.tx2.r_SM_MainZ0Z_2 ));
    Odrv4 I__2734 (
            .O(N__14367),
            .I(\c0.tx2.r_SM_MainZ0Z_2 ));
    InMux I__2733 (
            .O(N__14354),
            .I(N__14351));
    LocalMux I__2732 (
            .O(N__14351),
            .I(N__14344));
    InMux I__2731 (
            .O(N__14350),
            .I(N__14337));
    InMux I__2730 (
            .O(N__14349),
            .I(N__14330));
    InMux I__2729 (
            .O(N__14348),
            .I(N__14330));
    InMux I__2728 (
            .O(N__14347),
            .I(N__14330));
    Span4Mux_h I__2727 (
            .O(N__14344),
            .I(N__14327));
    InMux I__2726 (
            .O(N__14343),
            .I(N__14322));
    InMux I__2725 (
            .O(N__14342),
            .I(N__14322));
    InMux I__2724 (
            .O(N__14341),
            .I(N__14317));
    InMux I__2723 (
            .O(N__14340),
            .I(N__14317));
    LocalMux I__2722 (
            .O(N__14337),
            .I(N__14314));
    LocalMux I__2721 (
            .O(N__14330),
            .I(\c0.tx2.r_SM_MainZ0Z_0 ));
    Odrv4 I__2720 (
            .O(N__14327),
            .I(\c0.tx2.r_SM_MainZ0Z_0 ));
    LocalMux I__2719 (
            .O(N__14322),
            .I(\c0.tx2.r_SM_MainZ0Z_0 ));
    LocalMux I__2718 (
            .O(N__14317),
            .I(\c0.tx2.r_SM_MainZ0Z_0 ));
    Odrv4 I__2717 (
            .O(N__14314),
            .I(\c0.tx2.r_SM_MainZ0Z_0 ));
    CascadeMux I__2716 (
            .O(N__14303),
            .I(\c0.tx2.N_257_cascade_ ));
    InMux I__2715 (
            .O(N__14300),
            .I(N__14297));
    LocalMux I__2714 (
            .O(N__14297),
            .I(\c0.tx2.N_261 ));
    InMux I__2713 (
            .O(N__14294),
            .I(N__14288));
    CascadeMux I__2712 (
            .O(N__14293),
            .I(N__14284));
    CascadeMux I__2711 (
            .O(N__14292),
            .I(N__14281));
    CascadeMux I__2710 (
            .O(N__14291),
            .I(N__14278));
    LocalMux I__2709 (
            .O(N__14288),
            .I(N__14275));
    SRMux I__2708 (
            .O(N__14287),
            .I(N__14272));
    InMux I__2707 (
            .O(N__14284),
            .I(N__14269));
    InMux I__2706 (
            .O(N__14281),
            .I(N__14266));
    InMux I__2705 (
            .O(N__14278),
            .I(N__14263));
    Span4Mux_v I__2704 (
            .O(N__14275),
            .I(N__14260));
    LocalMux I__2703 (
            .O(N__14272),
            .I(N__14257));
    LocalMux I__2702 (
            .O(N__14269),
            .I(N__14246));
    LocalMux I__2701 (
            .O(N__14266),
            .I(N__14246));
    LocalMux I__2700 (
            .O(N__14263),
            .I(N__14246));
    Span4Mux_h I__2699 (
            .O(N__14260),
            .I(N__14246));
    Span4Mux_v I__2698 (
            .O(N__14257),
            .I(N__14246));
    Span4Mux_h I__2697 (
            .O(N__14246),
            .I(N__14243));
    Sp12to4 I__2696 (
            .O(N__14243),
            .I(N__14240));
    Odrv12 I__2695 (
            .O(N__14240),
            .I(\c0.tx2.o_Tx_Serial12 ));
    CascadeMux I__2694 (
            .O(N__14237),
            .I(\c0.tx2.N_261_cascade_ ));
    InMux I__2693 (
            .O(N__14234),
            .I(N__14229));
    CascadeMux I__2692 (
            .O(N__14233),
            .I(N__14226));
    InMux I__2691 (
            .O(N__14232),
            .I(N__14222));
    LocalMux I__2690 (
            .O(N__14229),
            .I(N__14219));
    InMux I__2689 (
            .O(N__14226),
            .I(N__14214));
    InMux I__2688 (
            .O(N__14225),
            .I(N__14214));
    LocalMux I__2687 (
            .O(N__14222),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    Odrv4 I__2686 (
            .O(N__14219),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    LocalMux I__2685 (
            .O(N__14214),
            .I(\c0.tx2.r_Bit_IndexZ0Z_2 ));
    InMux I__2684 (
            .O(N__14207),
            .I(N__14204));
    LocalMux I__2683 (
            .O(N__14204),
            .I(N__14201));
    Span4Mux_h I__2682 (
            .O(N__14201),
            .I(N__14196));
    InMux I__2681 (
            .O(N__14200),
            .I(N__14191));
    InMux I__2680 (
            .O(N__14199),
            .I(N__14191));
    Odrv4 I__2679 (
            .O(N__14196),
            .I(\c0.tx_transmitZ0 ));
    LocalMux I__2678 (
            .O(N__14191),
            .I(\c0.tx_transmitZ0 ));
    InMux I__2677 (
            .O(N__14186),
            .I(N__14179));
    InMux I__2676 (
            .O(N__14185),
            .I(N__14179));
    InMux I__2675 (
            .O(N__14184),
            .I(N__14176));
    LocalMux I__2674 (
            .O(N__14179),
            .I(N__14173));
    LocalMux I__2673 (
            .O(N__14176),
            .I(N__14168));
    Span4Mux_h I__2672 (
            .O(N__14173),
            .I(N__14168));
    Odrv4 I__2671 (
            .O(N__14168),
            .I(\c0.tx_active ));
    InMux I__2670 (
            .O(N__14165),
            .I(N__14162));
    LocalMux I__2669 (
            .O(N__14162),
            .I(N__14159));
    Span4Mux_h I__2668 (
            .O(N__14159),
            .I(N__14155));
    InMux I__2667 (
            .O(N__14158),
            .I(N__14152));
    Span4Mux_v I__2666 (
            .O(N__14155),
            .I(N__14147));
    LocalMux I__2665 (
            .O(N__14152),
            .I(N__14144));
    InMux I__2664 (
            .O(N__14151),
            .I(N__14139));
    InMux I__2663 (
            .O(N__14150),
            .I(N__14139));
    Odrv4 I__2662 (
            .O(N__14147),
            .I(\c0.d_4_34 ));
    Odrv4 I__2661 (
            .O(N__14144),
            .I(\c0.d_4_34 ));
    LocalMux I__2660 (
            .O(N__14139),
            .I(\c0.d_4_34 ));
    InMux I__2659 (
            .O(N__14132),
            .I(N__14129));
    LocalMux I__2658 (
            .O(N__14129),
            .I(N__14126));
    Span4Mux_h I__2657 (
            .O(N__14126),
            .I(N__14123));
    Odrv4 I__2656 (
            .O(N__14123),
            .I(\c0.un1_data_in_7__7_i ));
    InMux I__2655 (
            .O(N__14120),
            .I(N__14117));
    LocalMux I__2654 (
            .O(N__14117),
            .I(N__14114));
    Odrv12 I__2653 (
            .O(N__14114),
            .I(\c0.tx2_data_1_0_i_1_3 ));
    CascadeMux I__2652 (
            .O(N__14111),
            .I(N__14108));
    InMux I__2651 (
            .O(N__14108),
            .I(N__14105));
    LocalMux I__2650 (
            .O(N__14105),
            .I(N__14102));
    Span4Mux_h I__2649 (
            .O(N__14102),
            .I(N__14099));
    Span4Mux_h I__2648 (
            .O(N__14099),
            .I(N__14096));
    Odrv4 I__2647 (
            .O(N__14096),
            .I(\c0.tx2_data_1_iv_4_1_0_3 ));
    InMux I__2646 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__2645 (
            .O(N__14090),
            .I(N__14087));
    Span4Mux_v I__2644 (
            .O(N__14087),
            .I(N__14083));
    InMux I__2643 (
            .O(N__14086),
            .I(N__14079));
    Span4Mux_h I__2642 (
            .O(N__14083),
            .I(N__14076));
    InMux I__2641 (
            .O(N__14082),
            .I(N__14073));
    LocalMux I__2640 (
            .O(N__14079),
            .I(\c0.data_in_1_Z0Z_4 ));
    Odrv4 I__2639 (
            .O(N__14076),
            .I(\c0.data_in_1_Z0Z_4 ));
    LocalMux I__2638 (
            .O(N__14073),
            .I(\c0.data_in_1_Z0Z_4 ));
    InMux I__2637 (
            .O(N__14066),
            .I(N__14061));
    InMux I__2636 (
            .O(N__14065),
            .I(N__14058));
    CascadeMux I__2635 (
            .O(N__14064),
            .I(N__14055));
    LocalMux I__2634 (
            .O(N__14061),
            .I(N__14052));
    LocalMux I__2633 (
            .O(N__14058),
            .I(N__14049));
    InMux I__2632 (
            .O(N__14055),
            .I(N__14046));
    Span4Mux_h I__2631 (
            .O(N__14052),
            .I(N__14043));
    Span4Mux_v I__2630 (
            .O(N__14049),
            .I(N__14040));
    LocalMux I__2629 (
            .O(N__14046),
            .I(N__14037));
    Odrv4 I__2628 (
            .O(N__14043),
            .I(\c0.data_in_7_Z0Z_3 ));
    Odrv4 I__2627 (
            .O(N__14040),
            .I(\c0.data_in_7_Z0Z_3 ));
    Odrv12 I__2626 (
            .O(N__14037),
            .I(\c0.data_in_7_Z0Z_3 ));
    InMux I__2625 (
            .O(N__14030),
            .I(N__14027));
    LocalMux I__2624 (
            .O(N__14027),
            .I(\c0.data_in_frame_7_Z0Z_3 ));
    CascadeMux I__2623 (
            .O(N__14024),
            .I(N__14019));
    InMux I__2622 (
            .O(N__14023),
            .I(N__14016));
    InMux I__2621 (
            .O(N__14022),
            .I(N__14013));
    InMux I__2620 (
            .O(N__14019),
            .I(N__14010));
    LocalMux I__2619 (
            .O(N__14016),
            .I(N__14005));
    LocalMux I__2618 (
            .O(N__14013),
            .I(N__14002));
    LocalMux I__2617 (
            .O(N__14010),
            .I(N__13999));
    InMux I__2616 (
            .O(N__14009),
            .I(N__13996));
    CascadeMux I__2615 (
            .O(N__14008),
            .I(N__13993));
    Span4Mux_h I__2614 (
            .O(N__14005),
            .I(N__13990));
    Span4Mux_h I__2613 (
            .O(N__14002),
            .I(N__13987));
    Span4Mux_v I__2612 (
            .O(N__13999),
            .I(N__13982));
    LocalMux I__2611 (
            .O(N__13996),
            .I(N__13982));
    InMux I__2610 (
            .O(N__13993),
            .I(N__13979));
    Odrv4 I__2609 (
            .O(N__13990),
            .I(\c0.d_4_14 ));
    Odrv4 I__2608 (
            .O(N__13987),
            .I(\c0.d_4_14 ));
    Odrv4 I__2607 (
            .O(N__13982),
            .I(\c0.d_4_14 ));
    LocalMux I__2606 (
            .O(N__13979),
            .I(\c0.d_4_14 ));
    InMux I__2605 (
            .O(N__13970),
            .I(N__13966));
    CascadeMux I__2604 (
            .O(N__13969),
            .I(N__13963));
    LocalMux I__2603 (
            .O(N__13966),
            .I(N__13958));
    InMux I__2602 (
            .O(N__13963),
            .I(N__13955));
    InMux I__2601 (
            .O(N__13962),
            .I(N__13950));
    InMux I__2600 (
            .O(N__13961),
            .I(N__13950));
    Odrv4 I__2599 (
            .O(N__13958),
            .I(\c0.d_4_30 ));
    LocalMux I__2598 (
            .O(N__13955),
            .I(\c0.d_4_30 ));
    LocalMux I__2597 (
            .O(N__13950),
            .I(\c0.d_4_30 ));
    InMux I__2596 (
            .O(N__13943),
            .I(N__13940));
    LocalMux I__2595 (
            .O(N__13940),
            .I(N__13936));
    InMux I__2594 (
            .O(N__13939),
            .I(N__13933));
    Odrv4 I__2593 (
            .O(N__13936),
            .I(\c0.data_in_4_Z0Z_2 ));
    LocalMux I__2592 (
            .O(N__13933),
            .I(\c0.data_in_4_Z0Z_2 ));
    InMux I__2591 (
            .O(N__13928),
            .I(N__13924));
    InMux I__2590 (
            .O(N__13927),
            .I(N__13920));
    LocalMux I__2589 (
            .O(N__13924),
            .I(N__13917));
    CascadeMux I__2588 (
            .O(N__13923),
            .I(N__13914));
    LocalMux I__2587 (
            .O(N__13920),
            .I(N__13911));
    Span4Mux_v I__2586 (
            .O(N__13917),
            .I(N__13908));
    InMux I__2585 (
            .O(N__13914),
            .I(N__13905));
    Odrv4 I__2584 (
            .O(N__13911),
            .I(\c0.data_in_1_Z0Z_3 ));
    Odrv4 I__2583 (
            .O(N__13908),
            .I(\c0.data_in_1_Z0Z_3 ));
    LocalMux I__2582 (
            .O(N__13905),
            .I(\c0.data_in_1_Z0Z_3 ));
    InMux I__2581 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__2580 (
            .O(N__13895),
            .I(N__13892));
    Span4Mux_v I__2579 (
            .O(N__13892),
            .I(N__13888));
    InMux I__2578 (
            .O(N__13891),
            .I(N__13884));
    Span4Mux_h I__2577 (
            .O(N__13888),
            .I(N__13881));
    InMux I__2576 (
            .O(N__13887),
            .I(N__13878));
    LocalMux I__2575 (
            .O(N__13884),
            .I(\c0.data_in_1_Z0Z_5 ));
    Odrv4 I__2574 (
            .O(N__13881),
            .I(\c0.data_in_1_Z0Z_5 ));
    LocalMux I__2573 (
            .O(N__13878),
            .I(\c0.data_in_1_Z0Z_5 ));
    InMux I__2572 (
            .O(N__13871),
            .I(N__13868));
    LocalMux I__2571 (
            .O(N__13868),
            .I(N__13864));
    InMux I__2570 (
            .O(N__13867),
            .I(N__13860));
    Span4Mux_h I__2569 (
            .O(N__13864),
            .I(N__13857));
    InMux I__2568 (
            .O(N__13863),
            .I(N__13854));
    LocalMux I__2567 (
            .O(N__13860),
            .I(\c0.data_in_2_Z0Z_5 ));
    Odrv4 I__2566 (
            .O(N__13857),
            .I(\c0.data_in_2_Z0Z_5 ));
    LocalMux I__2565 (
            .O(N__13854),
            .I(\c0.data_in_2_Z0Z_5 ));
    InMux I__2564 (
            .O(N__13847),
            .I(N__13843));
    InMux I__2563 (
            .O(N__13846),
            .I(N__13840));
    LocalMux I__2562 (
            .O(N__13843),
            .I(N__13836));
    LocalMux I__2561 (
            .O(N__13840),
            .I(N__13833));
    InMux I__2560 (
            .O(N__13839),
            .I(N__13830));
    Odrv4 I__2559 (
            .O(N__13836),
            .I(\c0.data_in_3_Z0Z_1 ));
    Odrv4 I__2558 (
            .O(N__13833),
            .I(\c0.data_in_3_Z0Z_1 ));
    LocalMux I__2557 (
            .O(N__13830),
            .I(\c0.data_in_3_Z0Z_1 ));
    InMux I__2556 (
            .O(N__13823),
            .I(N__13820));
    LocalMux I__2555 (
            .O(N__13820),
            .I(N__13816));
    InMux I__2554 (
            .O(N__13819),
            .I(N__13813));
    Odrv4 I__2553 (
            .O(N__13816),
            .I(\c0.data_in_5_Z0Z_1 ));
    LocalMux I__2552 (
            .O(N__13813),
            .I(\c0.data_in_5_Z0Z_1 ));
    InMux I__2551 (
            .O(N__13808),
            .I(N__13805));
    LocalMux I__2550 (
            .O(N__13805),
            .I(N__13800));
    InMux I__2549 (
            .O(N__13804),
            .I(N__13795));
    InMux I__2548 (
            .O(N__13803),
            .I(N__13795));
    Odrv4 I__2547 (
            .O(N__13800),
            .I(\c0.data_in_3_Z0Z_3 ));
    LocalMux I__2546 (
            .O(N__13795),
            .I(\c0.data_in_3_Z0Z_3 ));
    CascadeMux I__2545 (
            .O(N__13790),
            .I(\c0.tx2_data_1_iv_3_1_6_cascade_ ));
    CascadeMux I__2544 (
            .O(N__13787),
            .I(\c0.un1_data_in_7__3_0_a2_0_a2_3_cascade_ ));
    InMux I__2543 (
            .O(N__13784),
            .I(N__13778));
    InMux I__2542 (
            .O(N__13783),
            .I(N__13775));
    InMux I__2541 (
            .O(N__13782),
            .I(N__13770));
    InMux I__2540 (
            .O(N__13781),
            .I(N__13770));
    LocalMux I__2539 (
            .O(N__13778),
            .I(\c0.N_129 ));
    LocalMux I__2538 (
            .O(N__13775),
            .I(\c0.N_129 ));
    LocalMux I__2537 (
            .O(N__13770),
            .I(\c0.N_129 ));
    InMux I__2536 (
            .O(N__13763),
            .I(N__13760));
    LocalMux I__2535 (
            .O(N__13760),
            .I(N__13757));
    Span4Mux_h I__2534 (
            .O(N__13757),
            .I(N__13752));
    InMux I__2533 (
            .O(N__13756),
            .I(N__13749));
    InMux I__2532 (
            .O(N__13755),
            .I(N__13746));
    Odrv4 I__2531 (
            .O(N__13752),
            .I(\c0.data_in_2_Z0Z_1 ));
    LocalMux I__2530 (
            .O(N__13749),
            .I(\c0.data_in_2_Z0Z_1 ));
    LocalMux I__2529 (
            .O(N__13746),
            .I(\c0.data_in_2_Z0Z_1 ));
    InMux I__2528 (
            .O(N__13739),
            .I(N__13735));
    InMux I__2527 (
            .O(N__13738),
            .I(N__13732));
    LocalMux I__2526 (
            .O(N__13735),
            .I(N__13726));
    LocalMux I__2525 (
            .O(N__13732),
            .I(N__13726));
    InMux I__2524 (
            .O(N__13731),
            .I(N__13722));
    Span4Mux_v I__2523 (
            .O(N__13726),
            .I(N__13719));
    InMux I__2522 (
            .O(N__13725),
            .I(N__13716));
    LocalMux I__2521 (
            .O(N__13722),
            .I(\c0.d_4_17 ));
    Odrv4 I__2520 (
            .O(N__13719),
            .I(\c0.d_4_17 ));
    LocalMux I__2519 (
            .O(N__13716),
            .I(\c0.d_4_17 ));
    InMux I__2518 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__2517 (
            .O(N__13706),
            .I(N__13702));
    CascadeMux I__2516 (
            .O(N__13705),
            .I(N__13698));
    Span4Mux_v I__2515 (
            .O(N__13702),
            .I(N__13695));
    InMux I__2514 (
            .O(N__13701),
            .I(N__13690));
    InMux I__2513 (
            .O(N__13698),
            .I(N__13690));
    Odrv4 I__2512 (
            .O(N__13695),
            .I(\c0.data_in_3_Z0Z_6 ));
    LocalMux I__2511 (
            .O(N__13690),
            .I(\c0.data_in_3_Z0Z_6 ));
    InMux I__2510 (
            .O(N__13685),
            .I(N__13682));
    LocalMux I__2509 (
            .O(N__13682),
            .I(N__13679));
    Span4Mux_h I__2508 (
            .O(N__13679),
            .I(N__13675));
    InMux I__2507 (
            .O(N__13678),
            .I(N__13672));
    Odrv4 I__2506 (
            .O(N__13675),
            .I(\c0.data_in_0_Z0Z_0 ));
    LocalMux I__2505 (
            .O(N__13672),
            .I(\c0.data_in_0_Z0Z_0 ));
    InMux I__2504 (
            .O(N__13667),
            .I(N__13664));
    LocalMux I__2503 (
            .O(N__13664),
            .I(N__13661));
    Span4Mux_h I__2502 (
            .O(N__13661),
            .I(N__13656));
    InMux I__2501 (
            .O(N__13660),
            .I(N__13653));
    InMux I__2500 (
            .O(N__13659),
            .I(N__13650));
    Odrv4 I__2499 (
            .O(N__13656),
            .I(\c0.data_in_2_Z0Z_0 ));
    LocalMux I__2498 (
            .O(N__13653),
            .I(\c0.data_in_2_Z0Z_0 ));
    LocalMux I__2497 (
            .O(N__13650),
            .I(\c0.data_in_2_Z0Z_0 ));
    InMux I__2496 (
            .O(N__13643),
            .I(N__13639));
    InMux I__2495 (
            .O(N__13642),
            .I(N__13636));
    LocalMux I__2494 (
            .O(N__13639),
            .I(N__13630));
    LocalMux I__2493 (
            .O(N__13636),
            .I(N__13630));
    InMux I__2492 (
            .O(N__13635),
            .I(N__13626));
    Span4Mux_v I__2491 (
            .O(N__13630),
            .I(N__13623));
    InMux I__2490 (
            .O(N__13629),
            .I(N__13620));
    LocalMux I__2489 (
            .O(N__13626),
            .I(\c0.d_4_16 ));
    Odrv4 I__2488 (
            .O(N__13623),
            .I(\c0.d_4_16 ));
    LocalMux I__2487 (
            .O(N__13620),
            .I(\c0.d_4_16 ));
    CascadeMux I__2486 (
            .O(N__13613),
            .I(N__13610));
    InMux I__2485 (
            .O(N__13610),
            .I(N__13604));
    InMux I__2484 (
            .O(N__13609),
            .I(N__13604));
    LocalMux I__2483 (
            .O(N__13604),
            .I(\c0.d_4_0 ));
    InMux I__2482 (
            .O(N__13601),
            .I(N__13598));
    LocalMux I__2481 (
            .O(N__13598),
            .I(N__13595));
    Span4Mux_v I__2480 (
            .O(N__13595),
            .I(N__13592));
    Odrv4 I__2479 (
            .O(N__13592),
            .I(\c0.tx2_data_RNO_3Z0Z_0 ));
    InMux I__2478 (
            .O(N__13589),
            .I(N__13586));
    LocalMux I__2477 (
            .O(N__13586),
            .I(N__13582));
    CascadeMux I__2476 (
            .O(N__13585),
            .I(N__13579));
    Span4Mux_v I__2475 (
            .O(N__13582),
            .I(N__13576));
    InMux I__2474 (
            .O(N__13579),
            .I(N__13573));
    Odrv4 I__2473 (
            .O(N__13576),
            .I(\c0.data_in_0_Z0Z_4 ));
    LocalMux I__2472 (
            .O(N__13573),
            .I(\c0.data_in_0_Z0Z_4 ));
    CascadeMux I__2471 (
            .O(N__13568),
            .I(\c0.wait_for_transmission_RNOZ0Z_10_cascade_ ));
    CascadeMux I__2470 (
            .O(N__13565),
            .I(N__13562));
    InMux I__2469 (
            .O(N__13562),
            .I(N__13559));
    LocalMux I__2468 (
            .O(N__13559),
            .I(N__13556));
    Span4Mux_h I__2467 (
            .O(N__13556),
            .I(N__13553));
    Odrv4 I__2466 (
            .O(N__13553),
            .I(\c0.g0_5_4 ));
    InMux I__2465 (
            .O(N__13550),
            .I(N__13547));
    LocalMux I__2464 (
            .O(N__13547),
            .I(N__13541));
    InMux I__2463 (
            .O(N__13546),
            .I(N__13538));
    InMux I__2462 (
            .O(N__13545),
            .I(N__13535));
    InMux I__2461 (
            .O(N__13544),
            .I(N__13532));
    Span4Mux_h I__2460 (
            .O(N__13541),
            .I(N__13529));
    LocalMux I__2459 (
            .O(N__13538),
            .I(N__13526));
    LocalMux I__2458 (
            .O(N__13535),
            .I(N__13521));
    LocalMux I__2457 (
            .O(N__13532),
            .I(N__13521));
    Odrv4 I__2456 (
            .O(N__13529),
            .I(\c0.d_4_3 ));
    Odrv12 I__2455 (
            .O(N__13526),
            .I(\c0.d_4_3 ));
    Odrv4 I__2454 (
            .O(N__13521),
            .I(\c0.d_4_3 ));
    CascadeMux I__2453 (
            .O(N__13514),
            .I(N__13511));
    InMux I__2452 (
            .O(N__13511),
            .I(N__13507));
    InMux I__2451 (
            .O(N__13510),
            .I(N__13504));
    LocalMux I__2450 (
            .O(N__13507),
            .I(N__13501));
    LocalMux I__2449 (
            .O(N__13504),
            .I(\c0.d_4_45 ));
    Odrv4 I__2448 (
            .O(N__13501),
            .I(\c0.d_4_45 ));
    CascadeMux I__2447 (
            .O(N__13496),
            .I(N__13493));
    InMux I__2446 (
            .O(N__13493),
            .I(N__13490));
    LocalMux I__2445 (
            .O(N__13490),
            .I(N__13487));
    Span4Mux_v I__2444 (
            .O(N__13487),
            .I(N__13484));
    Odrv4 I__2443 (
            .O(N__13484),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_2 ));
    CascadeMux I__2442 (
            .O(N__13481),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_3_cascade_ ));
    InMux I__2441 (
            .O(N__13478),
            .I(N__13475));
    LocalMux I__2440 (
            .O(N__13475),
            .I(\c0.un1_data_in_6__7_0_a2_17_a2_5 ));
    CascadeMux I__2439 (
            .O(N__13472),
            .I(N__13469));
    InMux I__2438 (
            .O(N__13469),
            .I(N__13466));
    LocalMux I__2437 (
            .O(N__13466),
            .I(N__13463));
    Span4Mux_h I__2436 (
            .O(N__13463),
            .I(N__13460));
    Span4Mux_h I__2435 (
            .O(N__13460),
            .I(N__13457));
    Odrv4 I__2434 (
            .O(N__13457),
            .I(\c0.g3_2_1 ));
    InMux I__2433 (
            .O(N__13454),
            .I(N__13451));
    LocalMux I__2432 (
            .O(N__13451),
            .I(\c0.g0_3_0 ));
    CascadeMux I__2431 (
            .O(N__13448),
            .I(\c0.un1_data_in_7__0_0_a2_1_a2_3_cascade_ ));
    CascadeMux I__2430 (
            .O(N__13445),
            .I(\c0.un1_data_in_7__0_0_a2_1_a2_5_0_cascade_ ));
    InMux I__2429 (
            .O(N__13442),
            .I(N__13439));
    LocalMux I__2428 (
            .O(N__13439),
            .I(\c0.tx2_transmit_0_sqmuxa_1 ));
    CascadeMux I__2427 (
            .O(N__13436),
            .I(N__13433));
    InMux I__2426 (
            .O(N__13433),
            .I(N__13429));
    CascadeMux I__2425 (
            .O(N__13432),
            .I(N__13426));
    LocalMux I__2424 (
            .O(N__13429),
            .I(N__13422));
    InMux I__2423 (
            .O(N__13426),
            .I(N__13419));
    CascadeMux I__2422 (
            .O(N__13425),
            .I(N__13415));
    Span4Mux_v I__2421 (
            .O(N__13422),
            .I(N__13410));
    LocalMux I__2420 (
            .O(N__13419),
            .I(N__13410));
    InMux I__2419 (
            .O(N__13418),
            .I(N__13405));
    InMux I__2418 (
            .O(N__13415),
            .I(N__13405));
    Span4Mux_h I__2417 (
            .O(N__13410),
            .I(N__13400));
    LocalMux I__2416 (
            .O(N__13405),
            .I(N__13400));
    Span4Mux_v I__2415 (
            .O(N__13400),
            .I(N__13397));
    Odrv4 I__2414 (
            .O(N__13397),
            .I(\c0.d_2_24 ));
    CascadeMux I__2413 (
            .O(N__13394),
            .I(N__13383));
    InMux I__2412 (
            .O(N__13393),
            .I(N__13370));
    InMux I__2411 (
            .O(N__13392),
            .I(N__13370));
    InMux I__2410 (
            .O(N__13391),
            .I(N__13370));
    InMux I__2409 (
            .O(N__13390),
            .I(N__13370));
    InMux I__2408 (
            .O(N__13389),
            .I(N__13370));
    InMux I__2407 (
            .O(N__13388),
            .I(N__13370));
    CascadeMux I__2406 (
            .O(N__13387),
            .I(N__13367));
    CascadeMux I__2405 (
            .O(N__13386),
            .I(N__13364));
    InMux I__2404 (
            .O(N__13383),
            .I(N__13345));
    LocalMux I__2403 (
            .O(N__13370),
            .I(N__13342));
    InMux I__2402 (
            .O(N__13367),
            .I(N__13331));
    InMux I__2401 (
            .O(N__13364),
            .I(N__13331));
    InMux I__2400 (
            .O(N__13363),
            .I(N__13331));
    InMux I__2399 (
            .O(N__13362),
            .I(N__13331));
    InMux I__2398 (
            .O(N__13361),
            .I(N__13331));
    InMux I__2397 (
            .O(N__13360),
            .I(N__13327));
    InMux I__2396 (
            .O(N__13359),
            .I(N__13320));
    InMux I__2395 (
            .O(N__13358),
            .I(N__13320));
    InMux I__2394 (
            .O(N__13357),
            .I(N__13320));
    InMux I__2393 (
            .O(N__13356),
            .I(N__13315));
    InMux I__2392 (
            .O(N__13355),
            .I(N__13315));
    InMux I__2391 (
            .O(N__13354),
            .I(N__13304));
    InMux I__2390 (
            .O(N__13353),
            .I(N__13304));
    InMux I__2389 (
            .O(N__13352),
            .I(N__13304));
    InMux I__2388 (
            .O(N__13351),
            .I(N__13304));
    InMux I__2387 (
            .O(N__13350),
            .I(N__13304));
    InMux I__2386 (
            .O(N__13349),
            .I(N__13295));
    InMux I__2385 (
            .O(N__13348),
            .I(N__13292));
    LocalMux I__2384 (
            .O(N__13345),
            .I(N__13289));
    Span4Mux_v I__2383 (
            .O(N__13342),
            .I(N__13284));
    LocalMux I__2382 (
            .O(N__13331),
            .I(N__13284));
    InMux I__2381 (
            .O(N__13330),
            .I(N__13281));
    LocalMux I__2380 (
            .O(N__13327),
            .I(N__13278));
    LocalMux I__2379 (
            .O(N__13320),
            .I(N__13271));
    LocalMux I__2378 (
            .O(N__13315),
            .I(N__13271));
    LocalMux I__2377 (
            .O(N__13304),
            .I(N__13271));
    CascadeMux I__2376 (
            .O(N__13303),
            .I(N__13268));
    CascadeMux I__2375 (
            .O(N__13302),
            .I(N__13265));
    CascadeMux I__2374 (
            .O(N__13301),
            .I(N__13262));
    InMux I__2373 (
            .O(N__13300),
            .I(N__13255));
    InMux I__2372 (
            .O(N__13299),
            .I(N__13255));
    InMux I__2371 (
            .O(N__13298),
            .I(N__13252));
    LocalMux I__2370 (
            .O(N__13295),
            .I(N__13246));
    LocalMux I__2369 (
            .O(N__13292),
            .I(N__13243));
    Span4Mux_h I__2368 (
            .O(N__13289),
            .I(N__13236));
    Span4Mux_h I__2367 (
            .O(N__13284),
            .I(N__13236));
    LocalMux I__2366 (
            .O(N__13281),
            .I(N__13236));
    Span4Mux_h I__2365 (
            .O(N__13278),
            .I(N__13231));
    Span4Mux_v I__2364 (
            .O(N__13271),
            .I(N__13231));
    InMux I__2363 (
            .O(N__13268),
            .I(N__13228));
    InMux I__2362 (
            .O(N__13265),
            .I(N__13219));
    InMux I__2361 (
            .O(N__13262),
            .I(N__13219));
    InMux I__2360 (
            .O(N__13261),
            .I(N__13219));
    InMux I__2359 (
            .O(N__13260),
            .I(N__13219));
    LocalMux I__2358 (
            .O(N__13255),
            .I(N__13214));
    LocalMux I__2357 (
            .O(N__13252),
            .I(N__13214));
    InMux I__2356 (
            .O(N__13251),
            .I(N__13207));
    InMux I__2355 (
            .O(N__13250),
            .I(N__13207));
    InMux I__2354 (
            .O(N__13249),
            .I(N__13207));
    Odrv12 I__2353 (
            .O(N__13246),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2352 (
            .O(N__13243),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2351 (
            .O(N__13236),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2350 (
            .O(N__13231),
            .I(CONSTANT_ONE_NET));
    LocalMux I__2349 (
            .O(N__13228),
            .I(CONSTANT_ONE_NET));
    LocalMux I__2348 (
            .O(N__13219),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2347 (
            .O(N__13214),
            .I(CONSTANT_ONE_NET));
    LocalMux I__2346 (
            .O(N__13207),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__2345 (
            .O(N__13190),
            .I(N__13187));
    InMux I__2344 (
            .O(N__13187),
            .I(N__13183));
    InMux I__2343 (
            .O(N__13186),
            .I(N__13180));
    LocalMux I__2342 (
            .O(N__13183),
            .I(N__13176));
    LocalMux I__2341 (
            .O(N__13180),
            .I(N__13173));
    InMux I__2340 (
            .O(N__13179),
            .I(N__13170));
    Odrv4 I__2339 (
            .O(N__13176),
            .I(\c0.N_105 ));
    Odrv4 I__2338 (
            .O(N__13173),
            .I(\c0.N_105 ));
    LocalMux I__2337 (
            .O(N__13170),
            .I(\c0.N_105 ));
    InMux I__2336 (
            .O(N__13163),
            .I(N__13160));
    LocalMux I__2335 (
            .O(N__13160),
            .I(N__13156));
    InMux I__2334 (
            .O(N__13159),
            .I(N__13153));
    Odrv4 I__2333 (
            .O(N__13156),
            .I(\c0.nextCRC16_3_2_1 ));
    LocalMux I__2332 (
            .O(N__13153),
            .I(\c0.nextCRC16_3_2_1 ));
    InMux I__2331 (
            .O(N__13148),
            .I(N__13144));
    InMux I__2330 (
            .O(N__13147),
            .I(N__13140));
    LocalMux I__2329 (
            .O(N__13144),
            .I(N__13137));
    InMux I__2328 (
            .O(N__13143),
            .I(N__13134));
    LocalMux I__2327 (
            .O(N__13140),
            .I(\c0.N_106 ));
    Odrv4 I__2326 (
            .O(N__13137),
            .I(\c0.N_106 ));
    LocalMux I__2325 (
            .O(N__13134),
            .I(\c0.N_106 ));
    CascadeMux I__2324 (
            .O(N__13127),
            .I(N__13124));
    InMux I__2323 (
            .O(N__13124),
            .I(N__13121));
    LocalMux I__2322 (
            .O(N__13121),
            .I(N__13118));
    Span4Mux_h I__2321 (
            .O(N__13118),
            .I(N__13115));
    Odrv4 I__2320 (
            .O(N__13115),
            .I(\c0.data_out_7_Z0Z_1 ));
    CascadeMux I__2319 (
            .O(N__13112),
            .I(N__13109));
    InMux I__2318 (
            .O(N__13109),
            .I(N__13106));
    LocalMux I__2317 (
            .O(N__13106),
            .I(\c0.data_in_frame_7_Z0Z_5 ));
    CascadeMux I__2316 (
            .O(N__13103),
            .I(N__13100));
    InMux I__2315 (
            .O(N__13100),
            .I(N__13097));
    LocalMux I__2314 (
            .O(N__13097),
            .I(\c0.data_in_frame_7_Z0Z_7 ));
    InMux I__2313 (
            .O(N__13094),
            .I(N__13087));
    InMux I__2312 (
            .O(N__13093),
            .I(N__13087));
    InMux I__2311 (
            .O(N__13092),
            .I(N__13084));
    LocalMux I__2310 (
            .O(N__13087),
            .I(N__13081));
    LocalMux I__2309 (
            .O(N__13084),
            .I(N__13078));
    Span4Mux_v I__2308 (
            .O(N__13081),
            .I(N__13075));
    Odrv4 I__2307 (
            .O(N__13078),
            .I(\c0.d_2_28 ));
    Odrv4 I__2306 (
            .O(N__13075),
            .I(\c0.d_2_28 ));
    InMux I__2305 (
            .O(N__13070),
            .I(N__13067));
    LocalMux I__2304 (
            .O(N__13067),
            .I(\c0.nextCRC16_3_0_a2_1_2 ));
    CascadeMux I__2303 (
            .O(N__13064),
            .I(N__13061));
    InMux I__2302 (
            .O(N__13061),
            .I(N__13056));
    InMux I__2301 (
            .O(N__13060),
            .I(N__13051));
    InMux I__2300 (
            .O(N__13059),
            .I(N__13051));
    LocalMux I__2299 (
            .O(N__13056),
            .I(\c0.d_2_0 ));
    LocalMux I__2298 (
            .O(N__13051),
            .I(\c0.d_2_0 ));
    InMux I__2297 (
            .O(N__13046),
            .I(N__13043));
    LocalMux I__2296 (
            .O(N__13043),
            .I(N__13040));
    Odrv4 I__2295 (
            .O(N__13040),
            .I(\c0.nextCRC16_3_4_0 ));
    CascadeMux I__2294 (
            .O(N__13037),
            .I(N__13034));
    InMux I__2293 (
            .O(N__13034),
            .I(N__13031));
    LocalMux I__2292 (
            .O(N__13031),
            .I(N__13026));
    InMux I__2291 (
            .O(N__13030),
            .I(N__13021));
    InMux I__2290 (
            .O(N__13029),
            .I(N__13021));
    Odrv4 I__2289 (
            .O(N__13026),
            .I(\c0.d_2_13 ));
    LocalMux I__2288 (
            .O(N__13021),
            .I(\c0.d_2_13 ));
    InMux I__2287 (
            .O(N__13016),
            .I(N__13013));
    LocalMux I__2286 (
            .O(N__13013),
            .I(N__13008));
    InMux I__2285 (
            .O(N__13012),
            .I(N__13005));
    CascadeMux I__2284 (
            .O(N__13011),
            .I(N__13000));
    Span4Mux_v I__2283 (
            .O(N__13008),
            .I(N__12995));
    LocalMux I__2282 (
            .O(N__13005),
            .I(N__12995));
    InMux I__2281 (
            .O(N__13004),
            .I(N__12992));
    InMux I__2280 (
            .O(N__13003),
            .I(N__12989));
    InMux I__2279 (
            .O(N__13000),
            .I(N__12986));
    Sp12to4 I__2278 (
            .O(N__12995),
            .I(N__12981));
    LocalMux I__2277 (
            .O(N__12992),
            .I(N__12981));
    LocalMux I__2276 (
            .O(N__12989),
            .I(\c0.d_2_26 ));
    LocalMux I__2275 (
            .O(N__12986),
            .I(\c0.d_2_26 ));
    Odrv12 I__2274 (
            .O(N__12981),
            .I(\c0.d_2_26 ));
    CascadeMux I__2273 (
            .O(N__12974),
            .I(\c0.nextCRC16_3_4_0_cascade_ ));
    InMux I__2272 (
            .O(N__12971),
            .I(N__12968));
    LocalMux I__2271 (
            .O(N__12968),
            .I(N__12964));
    InMux I__2270 (
            .O(N__12967),
            .I(N__12961));
    Span12Mux_s7_v I__2269 (
            .O(N__12964),
            .I(N__12957));
    LocalMux I__2268 (
            .O(N__12961),
            .I(N__12954));
    InMux I__2267 (
            .O(N__12960),
            .I(N__12951));
    Odrv12 I__2266 (
            .O(N__12957),
            .I(\c0.N_99 ));
    Odrv4 I__2265 (
            .O(N__12954),
            .I(\c0.N_99 ));
    LocalMux I__2264 (
            .O(N__12951),
            .I(\c0.N_99 ));
    InMux I__2263 (
            .O(N__12944),
            .I(N__12941));
    LocalMux I__2262 (
            .O(N__12941),
            .I(\c0.nextCRC16_3_0_a2_3_0 ));
    CascadeMux I__2261 (
            .O(N__12938),
            .I(N__12935));
    InMux I__2260 (
            .O(N__12935),
            .I(N__12929));
    InMux I__2259 (
            .O(N__12934),
            .I(N__12926));
    InMux I__2258 (
            .O(N__12933),
            .I(N__12923));
    InMux I__2257 (
            .O(N__12932),
            .I(N__12920));
    LocalMux I__2256 (
            .O(N__12929),
            .I(N__12916));
    LocalMux I__2255 (
            .O(N__12926),
            .I(N__12913));
    LocalMux I__2254 (
            .O(N__12923),
            .I(N__12910));
    LocalMux I__2253 (
            .O(N__12920),
            .I(N__12907));
    InMux I__2252 (
            .O(N__12919),
            .I(N__12904));
    Span4Mux_h I__2251 (
            .O(N__12916),
            .I(N__12901));
    Span4Mux_h I__2250 (
            .O(N__12913),
            .I(N__12896));
    Span4Mux_h I__2249 (
            .O(N__12910),
            .I(N__12896));
    Odrv12 I__2248 (
            .O(N__12907),
            .I(\c0.d_2_39 ));
    LocalMux I__2247 (
            .O(N__12904),
            .I(\c0.d_2_39 ));
    Odrv4 I__2246 (
            .O(N__12901),
            .I(\c0.d_2_39 ));
    Odrv4 I__2245 (
            .O(N__12896),
            .I(\c0.d_2_39 ));
    CascadeMux I__2244 (
            .O(N__12887),
            .I(N__12884));
    InMux I__2243 (
            .O(N__12884),
            .I(N__12881));
    LocalMux I__2242 (
            .O(N__12881),
            .I(N__12878));
    Span4Mux_h I__2241 (
            .O(N__12878),
            .I(N__12875));
    Odrv4 I__2240 (
            .O(N__12875),
            .I(\c0.data_out_6_Z0Z_5 ));
    InMux I__2239 (
            .O(N__12872),
            .I(N__12869));
    LocalMux I__2238 (
            .O(N__12869),
            .I(\c0.nextCRC16_3_0_a2_4_15 ));
    CascadeMux I__2237 (
            .O(N__12866),
            .I(N__12863));
    InMux I__2236 (
            .O(N__12863),
            .I(N__12860));
    LocalMux I__2235 (
            .O(N__12860),
            .I(N__12857));
    Span4Mux_h I__2234 (
            .O(N__12857),
            .I(N__12854));
    Odrv4 I__2233 (
            .O(N__12854),
            .I(\c0.nextCRC16_3_0_a2_3_15 ));
    InMux I__2232 (
            .O(N__12851),
            .I(N__12848));
    LocalMux I__2231 (
            .O(N__12848),
            .I(N__12845));
    Span4Mux_h I__2230 (
            .O(N__12845),
            .I(N__12842));
    Odrv4 I__2229 (
            .O(N__12842),
            .I(\c0.data_out_6_Z0Z_7 ));
    InMux I__2228 (
            .O(N__12839),
            .I(N__12835));
    InMux I__2227 (
            .O(N__12838),
            .I(N__12832));
    LocalMux I__2226 (
            .O(N__12835),
            .I(N__12829));
    LocalMux I__2225 (
            .O(N__12832),
            .I(N__12825));
    Span4Mux_h I__2224 (
            .O(N__12829),
            .I(N__12822));
    InMux I__2223 (
            .O(N__12828),
            .I(N__12817));
    Span4Mux_v I__2222 (
            .O(N__12825),
            .I(N__12814));
    Span4Mux_h I__2221 (
            .O(N__12822),
            .I(N__12811));
    InMux I__2220 (
            .O(N__12821),
            .I(N__12806));
    InMux I__2219 (
            .O(N__12820),
            .I(N__12806));
    LocalMux I__2218 (
            .O(N__12817),
            .I(N__12803));
    Odrv4 I__2217 (
            .O(N__12814),
            .I(\c0.d_2_16 ));
    Odrv4 I__2216 (
            .O(N__12811),
            .I(\c0.d_2_16 ));
    LocalMux I__2215 (
            .O(N__12806),
            .I(\c0.d_2_16 ));
    Odrv4 I__2214 (
            .O(N__12803),
            .I(\c0.d_2_16 ));
    InMux I__2213 (
            .O(N__12794),
            .I(N__12791));
    LocalMux I__2212 (
            .O(N__12791),
            .I(N__12787));
    InMux I__2211 (
            .O(N__12790),
            .I(N__12783));
    Span4Mux_h I__2210 (
            .O(N__12787),
            .I(N__12780));
    InMux I__2209 (
            .O(N__12786),
            .I(N__12777));
    LocalMux I__2208 (
            .O(N__12783),
            .I(\c0.d_2_9 ));
    Odrv4 I__2207 (
            .O(N__12780),
            .I(\c0.d_2_9 ));
    LocalMux I__2206 (
            .O(N__12777),
            .I(\c0.d_2_9 ));
    InMux I__2205 (
            .O(N__12770),
            .I(N__12766));
    InMux I__2204 (
            .O(N__12769),
            .I(N__12763));
    LocalMux I__2203 (
            .O(N__12766),
            .I(N__12760));
    LocalMux I__2202 (
            .O(N__12763),
            .I(N__12757));
    Span4Mux_h I__2201 (
            .O(N__12760),
            .I(N__12754));
    Span4Mux_h I__2200 (
            .O(N__12757),
            .I(N__12751));
    Odrv4 I__2199 (
            .O(N__12754),
            .I(\c0.N_94 ));
    Odrv4 I__2198 (
            .O(N__12751),
            .I(\c0.N_94 ));
    InMux I__2197 (
            .O(N__12746),
            .I(N__12743));
    LocalMux I__2196 (
            .O(N__12743),
            .I(N__12740));
    Span4Mux_h I__2195 (
            .O(N__12740),
            .I(N__12737));
    Span4Mux_h I__2194 (
            .O(N__12737),
            .I(N__12734));
    Odrv4 I__2193 (
            .O(N__12734),
            .I(\c0.tx_data_RNO_4Z0Z_5 ));
    InMux I__2192 (
            .O(N__12731),
            .I(N__12727));
    InMux I__2191 (
            .O(N__12730),
            .I(N__12724));
    LocalMux I__2190 (
            .O(N__12727),
            .I(N__12721));
    LocalMux I__2189 (
            .O(N__12724),
            .I(N__12718));
    Span4Mux_h I__2188 (
            .O(N__12721),
            .I(N__12715));
    Span4Mux_h I__2187 (
            .O(N__12718),
            .I(N__12712));
    Odrv4 I__2186 (
            .O(N__12715),
            .I(\c0.d_2_45 ));
    Odrv4 I__2185 (
            .O(N__12712),
            .I(\c0.d_2_45 ));
    InMux I__2184 (
            .O(N__12707),
            .I(N__12704));
    LocalMux I__2183 (
            .O(N__12704),
            .I(\c0.nextCRC16_3_0_a2_0_0 ));
    InMux I__2182 (
            .O(N__12701),
            .I(N__12698));
    LocalMux I__2181 (
            .O(N__12698),
            .I(\c0.nextCRC16_3_0_a2_4_0 ));
    InMux I__2180 (
            .O(N__12695),
            .I(N__12692));
    LocalMux I__2179 (
            .O(N__12692),
            .I(N__12689));
    Span4Mux_h I__2178 (
            .O(N__12689),
            .I(N__12686));
    Odrv4 I__2177 (
            .O(N__12686),
            .I(\c0.tx2.r_Tx_DataZ0Z_3 ));
    CascadeMux I__2176 (
            .O(N__12683),
            .I(\c0.tx2.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_ ));
    InMux I__2175 (
            .O(N__12680),
            .I(N__12677));
    LocalMux I__2174 (
            .O(N__12677),
            .I(\c0.tx2.N_349 ));
    CascadeMux I__2173 (
            .O(N__12674),
            .I(\c0.tx2.N_346_cascade_ ));
    CascadeMux I__2172 (
            .O(N__12671),
            .I(\c0.tx2.N_279_cascade_ ));
    IoInMux I__2171 (
            .O(N__12668),
            .I(N__12665));
    LocalMux I__2170 (
            .O(N__12665),
            .I(N__12661));
    InMux I__2169 (
            .O(N__12664),
            .I(N__12658));
    Span12Mux_s11_h I__2168 (
            .O(N__12661),
            .I(N__12655));
    LocalMux I__2167 (
            .O(N__12658),
            .I(N__12652));
    Odrv12 I__2166 (
            .O(N__12655),
            .I(PIN_3_c));
    Odrv4 I__2165 (
            .O(N__12652),
            .I(PIN_3_c));
    InMux I__2164 (
            .O(N__12647),
            .I(N__12644));
    LocalMux I__2163 (
            .O(N__12644),
            .I(N__12641));
    Span12Mux_v I__2162 (
            .O(N__12641),
            .I(N__12638));
    Odrv12 I__2161 (
            .O(N__12638),
            .I(\c0.tx2.r_Tx_Active_1_sqmuxa ));
    InMux I__2160 (
            .O(N__12635),
            .I(N__12632));
    LocalMux I__2159 (
            .O(N__12632),
            .I(N__12629));
    Odrv4 I__2158 (
            .O(N__12629),
            .I(\c0.tx_data_RNO_3Z0Z_1 ));
    CascadeMux I__2157 (
            .O(N__12626),
            .I(\c0.tx2.m5_0_0_cascade_ ));
    InMux I__2156 (
            .O(N__12623),
            .I(N__12620));
    LocalMux I__2155 (
            .O(N__12620),
            .I(N__12617));
    Span4Mux_v I__2154 (
            .O(N__12617),
            .I(N__12614));
    Odrv4 I__2153 (
            .O(N__12614),
            .I(\c0.tx2_data_RNO_0Z0Z_0 ));
    CascadeMux I__2152 (
            .O(N__12611),
            .I(\c0.tx2_data_1_0_i_ns_1_0_cascade_ ));
    CascadeMux I__2151 (
            .O(N__12608),
            .I(N__12605));
    InMux I__2150 (
            .O(N__12605),
            .I(N__12602));
    LocalMux I__2149 (
            .O(N__12602),
            .I(N__12595));
    InMux I__2148 (
            .O(N__12601),
            .I(N__12592));
    InMux I__2147 (
            .O(N__12600),
            .I(N__12587));
    InMux I__2146 (
            .O(N__12599),
            .I(N__12587));
    InMux I__2145 (
            .O(N__12598),
            .I(N__12584));
    Odrv12 I__2144 (
            .O(N__12595),
            .I(\c0.d_4_1 ));
    LocalMux I__2143 (
            .O(N__12592),
            .I(\c0.d_4_1 ));
    LocalMux I__2142 (
            .O(N__12587),
            .I(\c0.d_4_1 ));
    LocalMux I__2141 (
            .O(N__12584),
            .I(\c0.d_4_1 ));
    CascadeMux I__2140 (
            .O(N__12575),
            .I(\c0.tx2_data_RNO_3Z0Z_1_cascade_ ));
    InMux I__2139 (
            .O(N__12572),
            .I(N__12569));
    LocalMux I__2138 (
            .O(N__12569),
            .I(N__12566));
    Span4Mux_v I__2137 (
            .O(N__12566),
            .I(N__12563));
    Odrv4 I__2136 (
            .O(N__12563),
            .I(\c0.tx2_data_RNO_1Z0Z_1 ));
    CascadeMux I__2135 (
            .O(N__12560),
            .I(\c0.tx2_data_1_0_i_ns_1_1_cascade_ ));
    InMux I__2134 (
            .O(N__12557),
            .I(N__12554));
    LocalMux I__2133 (
            .O(N__12554),
            .I(N__12551));
    Span4Mux_v I__2132 (
            .O(N__12551),
            .I(N__12548));
    Odrv4 I__2131 (
            .O(N__12548),
            .I(\c0.tx2_data_RNO_0Z0Z_1 ));
    InMux I__2130 (
            .O(N__12545),
            .I(N__12542));
    LocalMux I__2129 (
            .O(N__12542),
            .I(\c0.tx2_data_RNO_4Z0Z_1 ));
    InMux I__2128 (
            .O(N__12539),
            .I(N__12536));
    LocalMux I__2127 (
            .O(N__12536),
            .I(\c0.tx2_data_RNO_1Z0Z_0 ));
    InMux I__2126 (
            .O(N__12533),
            .I(N__12530));
    LocalMux I__2125 (
            .O(N__12530),
            .I(N__12527));
    Span4Mux_v I__2124 (
            .O(N__12527),
            .I(N__12524));
    Odrv4 I__2123 (
            .O(N__12524),
            .I(\c0.tx2.r_Tx_DataZ0Z_2 ));
    InMux I__2122 (
            .O(N__12521),
            .I(N__12518));
    LocalMux I__2121 (
            .O(N__12518),
            .I(\c0.tx2.r_Tx_DataZ0Z_0 ));
    InMux I__2120 (
            .O(N__12515),
            .I(N__12512));
    LocalMux I__2119 (
            .O(N__12512),
            .I(\c0.tx2.r_Tx_Data_pmux_3_i_m2_ns_1 ));
    InMux I__2118 (
            .O(N__12509),
            .I(N__12506));
    LocalMux I__2117 (
            .O(N__12506),
            .I(\c0.tx2.r_Tx_DataZ0Z_1 ));
    CascadeMux I__2116 (
            .O(N__12503),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_2_cascade_ ));
    InMux I__2115 (
            .O(N__12500),
            .I(N__12497));
    LocalMux I__2114 (
            .O(N__12497),
            .I(N__12493));
    CascadeMux I__2113 (
            .O(N__12496),
            .I(N__12488));
    Span4Mux_h I__2112 (
            .O(N__12493),
            .I(N__12484));
    InMux I__2111 (
            .O(N__12492),
            .I(N__12481));
    InMux I__2110 (
            .O(N__12491),
            .I(N__12474));
    InMux I__2109 (
            .O(N__12488),
            .I(N__12474));
    InMux I__2108 (
            .O(N__12487),
            .I(N__12474));
    Odrv4 I__2107 (
            .O(N__12484),
            .I(\c0.d_4_2 ));
    LocalMux I__2106 (
            .O(N__12481),
            .I(\c0.d_4_2 ));
    LocalMux I__2105 (
            .O(N__12474),
            .I(\c0.d_4_2 ));
    InMux I__2104 (
            .O(N__12467),
            .I(N__12464));
    LocalMux I__2103 (
            .O(N__12464),
            .I(N__12460));
    InMux I__2102 (
            .O(N__12463),
            .I(N__12457));
    Odrv4 I__2101 (
            .O(N__12460),
            .I(\c0.N_103 ));
    LocalMux I__2100 (
            .O(N__12457),
            .I(\c0.N_103 ));
    InMux I__2099 (
            .O(N__12452),
            .I(N__12449));
    LocalMux I__2098 (
            .O(N__12449),
            .I(\c0.wait_for_transmission4_13_1_1 ));
    CascadeMux I__2097 (
            .O(N__12446),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_6_cascade_ ));
    CascadeMux I__2096 (
            .O(N__12443),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_1_cascade_ ));
    InMux I__2095 (
            .O(N__12440),
            .I(N__12437));
    LocalMux I__2094 (
            .O(N__12437),
            .I(\c0.un1_data_in_7__1_0_a2_24_a2_5 ));
    InMux I__2093 (
            .O(N__12434),
            .I(N__12431));
    LocalMux I__2092 (
            .O(N__12431),
            .I(N__12428));
    Odrv4 I__2091 (
            .O(N__12428),
            .I(\c0.d_4_RNITCRCZ0Z_29 ));
    CascadeMux I__2090 (
            .O(N__12425),
            .I(\c0.tx2_data_RNO_4Z0Z_0_cascade_ ));
    InMux I__2089 (
            .O(N__12422),
            .I(N__12419));
    LocalMux I__2088 (
            .O(N__12419),
            .I(N__12416));
    Odrv4 I__2087 (
            .O(N__12416),
            .I(\c0.un1_data_in_7__4_0_a2_0_a2_4 ));
    InMux I__2086 (
            .O(N__12413),
            .I(N__12410));
    LocalMux I__2085 (
            .O(N__12410),
            .I(N__12406));
    CascadeMux I__2084 (
            .O(N__12409),
            .I(N__12403));
    Span4Mux_h I__2083 (
            .O(N__12406),
            .I(N__12400));
    InMux I__2082 (
            .O(N__12403),
            .I(N__12397));
    Odrv4 I__2081 (
            .O(N__12400),
            .I(\c0.data_in_0_Z0Z_2 ));
    LocalMux I__2080 (
            .O(N__12397),
            .I(\c0.data_in_0_Z0Z_2 ));
    InMux I__2079 (
            .O(N__12392),
            .I(N__12389));
    LocalMux I__2078 (
            .O(N__12389),
            .I(\c0.d_4_RNID6K21_0Z0Z_15 ));
    InMux I__2077 (
            .O(N__12386),
            .I(N__12383));
    LocalMux I__2076 (
            .O(N__12383),
            .I(\c0.d_4_RNID6K21Z0Z_15 ));
    InMux I__2075 (
            .O(N__12380),
            .I(N__12377));
    LocalMux I__2074 (
            .O(N__12377),
            .I(N__12374));
    Span4Mux_v I__2073 (
            .O(N__12374),
            .I(N__12370));
    InMux I__2072 (
            .O(N__12373),
            .I(N__12367));
    Odrv4 I__2071 (
            .O(N__12370),
            .I(\c0.data_in_0_Z0Z_1 ));
    LocalMux I__2070 (
            .O(N__12367),
            .I(\c0.data_in_0_Z0Z_1 ));
    InMux I__2069 (
            .O(N__12362),
            .I(N__12357));
    CascadeMux I__2068 (
            .O(N__12361),
            .I(N__12354));
    InMux I__2067 (
            .O(N__12360),
            .I(N__12351));
    LocalMux I__2066 (
            .O(N__12357),
            .I(N__12348));
    InMux I__2065 (
            .O(N__12354),
            .I(N__12345));
    LocalMux I__2064 (
            .O(N__12351),
            .I(N__12340));
    Span4Mux_h I__2063 (
            .O(N__12348),
            .I(N__12340));
    LocalMux I__2062 (
            .O(N__12345),
            .I(N__12337));
    Odrv4 I__2061 (
            .O(N__12340),
            .I(\c0.data_in_1_Z0Z_7 ));
    Odrv4 I__2060 (
            .O(N__12337),
            .I(\c0.data_in_1_Z0Z_7 ));
    InMux I__2059 (
            .O(N__12332),
            .I(N__12328));
    InMux I__2058 (
            .O(N__12331),
            .I(N__12325));
    LocalMux I__2057 (
            .O(N__12328),
            .I(N__12321));
    LocalMux I__2056 (
            .O(N__12325),
            .I(N__12318));
    InMux I__2055 (
            .O(N__12324),
            .I(N__12315));
    Odrv4 I__2054 (
            .O(N__12321),
            .I(\c0.data_in_3_Z0Z_7 ));
    Odrv4 I__2053 (
            .O(N__12318),
            .I(\c0.data_in_3_Z0Z_7 ));
    LocalMux I__2052 (
            .O(N__12315),
            .I(\c0.data_in_3_Z0Z_7 ));
    CascadeMux I__2051 (
            .O(N__12308),
            .I(\c0.un1_data_in_6__0_0_a2_5_a2_2_cascade_ ));
    CascadeMux I__2050 (
            .O(N__12305),
            .I(\c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_ ));
    CascadeMux I__2049 (
            .O(N__12302),
            .I(\c0.un1_data_in_7__4_i_cascade_ ));
    InMux I__2048 (
            .O(N__12299),
            .I(N__12296));
    LocalMux I__2047 (
            .O(N__12296),
            .I(\c0.un1_data_in_6__0 ));
    CascadeMux I__2046 (
            .O(N__12293),
            .I(\c0.d_4_RNIF73E2Z0Z_14_cascade_ ));
    CascadeMux I__2045 (
            .O(N__12290),
            .I(\c0.d_4_RNIMKFE3Z0Z_14_cascade_ ));
    CascadeMux I__2044 (
            .O(N__12287),
            .I(\c0.un1_data_in_6__7_cascade_ ));
    InMux I__2043 (
            .O(N__12284),
            .I(N__12281));
    LocalMux I__2042 (
            .O(N__12281),
            .I(\c0.wait_for_transmission4_12 ));
    IoInMux I__2041 (
            .O(N__12278),
            .I(N__12275));
    LocalMux I__2040 (
            .O(N__12275),
            .I(N__12272));
    IoSpan4Mux I__2039 (
            .O(N__12272),
            .I(N__12269));
    Span4Mux_s2_h I__2038 (
            .O(N__12269),
            .I(N__12266));
    Sp12to4 I__2037 (
            .O(N__12266),
            .I(N__12262));
    InMux I__2036 (
            .O(N__12265),
            .I(N__12259));
    Span12Mux_s10_h I__2035 (
            .O(N__12262),
            .I(N__12256));
    LocalMux I__2034 (
            .O(N__12259),
            .I(\c0.data_in_frame_0__0_sqmuxa ));
    Odrv12 I__2033 (
            .O(N__12256),
            .I(\c0.data_in_frame_0__0_sqmuxa ));
    CascadeMux I__2032 (
            .O(N__12251),
            .I(\c0.wait_for_transmission4_12_cascade_ ));
    InMux I__2031 (
            .O(N__12248),
            .I(N__12245));
    LocalMux I__2030 (
            .O(N__12245),
            .I(N__12241));
    InMux I__2029 (
            .O(N__12244),
            .I(N__12238));
    Odrv4 I__2028 (
            .O(N__12241),
            .I(\c0.dataZ0Z_15 ));
    LocalMux I__2027 (
            .O(N__12238),
            .I(\c0.dataZ0Z_15 ));
    InMux I__2026 (
            .O(N__12233),
            .I(N__12226));
    InMux I__2025 (
            .O(N__12232),
            .I(N__12226));
    InMux I__2024 (
            .O(N__12231),
            .I(N__12223));
    LocalMux I__2023 (
            .O(N__12226),
            .I(N__12220));
    LocalMux I__2022 (
            .O(N__12223),
            .I(\c0.tx2_active ));
    Odrv4 I__2021 (
            .O(N__12220),
            .I(\c0.tx2_active ));
    InMux I__2020 (
            .O(N__12215),
            .I(N__12212));
    LocalMux I__2019 (
            .O(N__12212),
            .I(\c0.tx2_data_1_iv_5_1_0_7 ));
    CascadeMux I__2018 (
            .O(N__12209),
            .I(\c0.tx2_data_1_iv_5_1_7_cascade_ ));
    InMux I__2017 (
            .O(N__12206),
            .I(N__12203));
    LocalMux I__2016 (
            .O(N__12203),
            .I(\c0.data_in_frame_6_Z0Z_7 ));
    InMux I__2015 (
            .O(N__12200),
            .I(N__12197));
    LocalMux I__2014 (
            .O(N__12197),
            .I(N__12194));
    Span4Mux_h I__2013 (
            .O(N__12194),
            .I(N__12191));
    Odrv4 I__2012 (
            .O(N__12191),
            .I(\c0.tx2_data_1_iv_3_1_3 ));
    CascadeMux I__2011 (
            .O(N__12188),
            .I(N__12185));
    InMux I__2010 (
            .O(N__12185),
            .I(N__12182));
    LocalMux I__2009 (
            .O(N__12182),
            .I(N__12179));
    Span4Mux_v I__2008 (
            .O(N__12179),
            .I(N__12176));
    Odrv4 I__2007 (
            .O(N__12176),
            .I(\c0.tx2_data_1_iv_3_3 ));
    InMux I__2006 (
            .O(N__12173),
            .I(N__12170));
    LocalMux I__2005 (
            .O(N__12170),
            .I(N__12167));
    Span4Mux_h I__2004 (
            .O(N__12167),
            .I(N__12163));
    InMux I__2003 (
            .O(N__12166),
            .I(N__12160));
    Odrv4 I__2002 (
            .O(N__12163),
            .I(\c0.data_in_0_Z0Z_3 ));
    LocalMux I__2001 (
            .O(N__12160),
            .I(\c0.data_in_0_Z0Z_3 ));
    InMux I__2000 (
            .O(N__12155),
            .I(N__12152));
    LocalMux I__1999 (
            .O(N__12152),
            .I(\c0.N_247_0 ));
    InMux I__1998 (
            .O(N__12149),
            .I(N__12145));
    CascadeMux I__1997 (
            .O(N__12148),
            .I(N__12141));
    LocalMux I__1996 (
            .O(N__12145),
            .I(N__12138));
    InMux I__1995 (
            .O(N__12144),
            .I(N__12133));
    InMux I__1994 (
            .O(N__12141),
            .I(N__12133));
    Span4Mux_h I__1993 (
            .O(N__12138),
            .I(N__12130));
    LocalMux I__1992 (
            .O(N__12133),
            .I(\c0.d_2_41 ));
    Odrv4 I__1991 (
            .O(N__12130),
            .I(\c0.d_2_41 ));
    InMux I__1990 (
            .O(N__12125),
            .I(N__12118));
    InMux I__1989 (
            .O(N__12124),
            .I(N__12118));
    InMux I__1988 (
            .O(N__12123),
            .I(N__12115));
    LocalMux I__1987 (
            .O(N__12118),
            .I(\c0.d_2_12 ));
    LocalMux I__1986 (
            .O(N__12115),
            .I(\c0.d_2_12 ));
    InMux I__1985 (
            .O(N__12110),
            .I(N__12107));
    LocalMux I__1984 (
            .O(N__12107),
            .I(N__12102));
    InMux I__1983 (
            .O(N__12106),
            .I(N__12099));
    CascadeMux I__1982 (
            .O(N__12105),
            .I(N__12094));
    Span4Mux_v I__1981 (
            .O(N__12102),
            .I(N__12089));
    LocalMux I__1980 (
            .O(N__12099),
            .I(N__12089));
    InMux I__1979 (
            .O(N__12098),
            .I(N__12086));
    InMux I__1978 (
            .O(N__12097),
            .I(N__12083));
    InMux I__1977 (
            .O(N__12094),
            .I(N__12080));
    Odrv4 I__1976 (
            .O(N__12089),
            .I(\c0.d_2_40 ));
    LocalMux I__1975 (
            .O(N__12086),
            .I(\c0.d_2_40 ));
    LocalMux I__1974 (
            .O(N__12083),
            .I(\c0.d_2_40 ));
    LocalMux I__1973 (
            .O(N__12080),
            .I(\c0.d_2_40 ));
    InMux I__1972 (
            .O(N__12071),
            .I(N__12068));
    LocalMux I__1971 (
            .O(N__12068),
            .I(\c0.nextCRC16_3_0_a2_2_2 ));
    InMux I__1970 (
            .O(N__12065),
            .I(N__12061));
    InMux I__1969 (
            .O(N__12064),
            .I(N__12058));
    LocalMux I__1968 (
            .O(N__12061),
            .I(N__12055));
    LocalMux I__1967 (
            .O(N__12058),
            .I(N__12052));
    Span4Mux_h I__1966 (
            .O(N__12055),
            .I(N__12049));
    Span4Mux_v I__1965 (
            .O(N__12052),
            .I(N__12046));
    Span4Mux_h I__1964 (
            .O(N__12049),
            .I(N__12043));
    Odrv4 I__1963 (
            .O(N__12046),
            .I(\c0.d_2_3 ));
    Odrv4 I__1962 (
            .O(N__12043),
            .I(\c0.d_2_3 ));
    InMux I__1961 (
            .O(N__12038),
            .I(N__12035));
    LocalMux I__1960 (
            .O(N__12035),
            .I(N__12031));
    InMux I__1959 (
            .O(N__12034),
            .I(N__12028));
    Odrv12 I__1958 (
            .O(N__12031),
            .I(\c0.N_75 ));
    LocalMux I__1957 (
            .O(N__12028),
            .I(\c0.N_75 ));
    CascadeMux I__1956 (
            .O(N__12023),
            .I(\c0.N_75_cascade_ ));
    CascadeMux I__1955 (
            .O(N__12020),
            .I(N__12017));
    InMux I__1954 (
            .O(N__12017),
            .I(N__12014));
    LocalMux I__1953 (
            .O(N__12014),
            .I(N__12010));
    InMux I__1952 (
            .O(N__12013),
            .I(N__12007));
    Odrv4 I__1951 (
            .O(N__12010),
            .I(\c0.d_2_44 ));
    LocalMux I__1950 (
            .O(N__12007),
            .I(\c0.d_2_44 ));
    InMux I__1949 (
            .O(N__12002),
            .I(N__11999));
    LocalMux I__1948 (
            .O(N__11999),
            .I(\c0.N_95 ));
    CascadeMux I__1947 (
            .O(N__11996),
            .I(N__11992));
    CascadeMux I__1946 (
            .O(N__11995),
            .I(N__11988));
    InMux I__1945 (
            .O(N__11992),
            .I(N__11985));
    InMux I__1944 (
            .O(N__11991),
            .I(N__11982));
    InMux I__1943 (
            .O(N__11988),
            .I(N__11979));
    LocalMux I__1942 (
            .O(N__11985),
            .I(N__11974));
    LocalMux I__1941 (
            .O(N__11982),
            .I(N__11974));
    LocalMux I__1940 (
            .O(N__11979),
            .I(N__11971));
    Span4Mux_h I__1939 (
            .O(N__11974),
            .I(N__11968));
    Span4Mux_v I__1938 (
            .O(N__11971),
            .I(N__11965));
    Odrv4 I__1937 (
            .O(N__11968),
            .I(\c0.d_2_14 ));
    Odrv4 I__1936 (
            .O(N__11965),
            .I(\c0.d_2_14 ));
    CascadeMux I__1935 (
            .O(N__11960),
            .I(\c0.N_95_cascade_ ));
    InMux I__1934 (
            .O(N__11957),
            .I(N__11951));
    InMux I__1933 (
            .O(N__11956),
            .I(N__11948));
    InMux I__1932 (
            .O(N__11955),
            .I(N__11945));
    InMux I__1931 (
            .O(N__11954),
            .I(N__11942));
    LocalMux I__1930 (
            .O(N__11951),
            .I(N__11939));
    LocalMux I__1929 (
            .O(N__11948),
            .I(N__11936));
    LocalMux I__1928 (
            .O(N__11945),
            .I(N__11933));
    LocalMux I__1927 (
            .O(N__11942),
            .I(N__11930));
    Span4Mux_h I__1926 (
            .O(N__11939),
            .I(N__11927));
    Span4Mux_v I__1925 (
            .O(N__11936),
            .I(N__11924));
    Span4Mux_v I__1924 (
            .O(N__11933),
            .I(N__11919));
    Span4Mux_h I__1923 (
            .O(N__11930),
            .I(N__11919));
    Odrv4 I__1922 (
            .O(N__11927),
            .I(\c0.d_2_25 ));
    Odrv4 I__1921 (
            .O(N__11924),
            .I(\c0.d_2_25 ));
    Odrv4 I__1920 (
            .O(N__11919),
            .I(\c0.d_2_25 ));
    InMux I__1919 (
            .O(N__11912),
            .I(N__11908));
    InMux I__1918 (
            .O(N__11911),
            .I(N__11904));
    LocalMux I__1917 (
            .O(N__11908),
            .I(N__11900));
    InMux I__1916 (
            .O(N__11907),
            .I(N__11897));
    LocalMux I__1915 (
            .O(N__11904),
            .I(N__11894));
    CascadeMux I__1914 (
            .O(N__11903),
            .I(N__11891));
    Span4Mux_v I__1913 (
            .O(N__11900),
            .I(N__11888));
    LocalMux I__1912 (
            .O(N__11897),
            .I(N__11883));
    Span12Mux_s6_v I__1911 (
            .O(N__11894),
            .I(N__11883));
    InMux I__1910 (
            .O(N__11891),
            .I(N__11880));
    Odrv4 I__1909 (
            .O(N__11888),
            .I(\c0.d_2_11 ));
    Odrv12 I__1908 (
            .O(N__11883),
            .I(\c0.d_2_11 ));
    LocalMux I__1907 (
            .O(N__11880),
            .I(\c0.d_2_11 ));
    InMux I__1906 (
            .O(N__11873),
            .I(N__11870));
    LocalMux I__1905 (
            .O(N__11870),
            .I(N__11866));
    InMux I__1904 (
            .O(N__11869),
            .I(N__11863));
    Odrv4 I__1903 (
            .O(N__11866),
            .I(\c0.dataZ0Z_8 ));
    LocalMux I__1902 (
            .O(N__11863),
            .I(\c0.dataZ0Z_8 ));
    CascadeMux I__1901 (
            .O(N__11858),
            .I(N__11855));
    InMux I__1900 (
            .O(N__11855),
            .I(N__11852));
    LocalMux I__1899 (
            .O(N__11852),
            .I(\c0.nextCRC16_3_0_a2_1_8 ));
    InMux I__1898 (
            .O(N__11849),
            .I(N__11845));
    InMux I__1897 (
            .O(N__11848),
            .I(N__11842));
    LocalMux I__1896 (
            .O(N__11845),
            .I(N__11837));
    LocalMux I__1895 (
            .O(N__11842),
            .I(N__11837));
    Span4Mux_h I__1894 (
            .O(N__11837),
            .I(N__11834));
    Span4Mux_h I__1893 (
            .O(N__11834),
            .I(N__11830));
    InMux I__1892 (
            .O(N__11833),
            .I(N__11827));
    Odrv4 I__1891 (
            .O(N__11830),
            .I(\c0.N_77 ));
    LocalMux I__1890 (
            .O(N__11827),
            .I(\c0.N_77 ));
    InMux I__1889 (
            .O(N__11822),
            .I(N__11819));
    LocalMux I__1888 (
            .O(N__11819),
            .I(\c0.data_out_6_Z0Z_0 ));
    InMux I__1887 (
            .O(N__11816),
            .I(N__11813));
    LocalMux I__1886 (
            .O(N__11813),
            .I(N__11810));
    Span4Mux_h I__1885 (
            .O(N__11810),
            .I(N__11806));
    InMux I__1884 (
            .O(N__11809),
            .I(N__11803));
    Odrv4 I__1883 (
            .O(N__11806),
            .I(\c0.dataZ0Z_0 ));
    LocalMux I__1882 (
            .O(N__11803),
            .I(\c0.dataZ0Z_0 ));
    InMux I__1881 (
            .O(N__11798),
            .I(N__11795));
    LocalMux I__1880 (
            .O(N__11795),
            .I(\c0.data_out_7_Z0Z_0 ));
    InMux I__1879 (
            .O(N__11792),
            .I(N__11789));
    LocalMux I__1878 (
            .O(N__11789),
            .I(N__11785));
    InMux I__1877 (
            .O(N__11788),
            .I(N__11782));
    Odrv4 I__1876 (
            .O(N__11785),
            .I(\c0.d_2_8 ));
    LocalMux I__1875 (
            .O(N__11782),
            .I(\c0.d_2_8 ));
    InMux I__1874 (
            .O(N__11777),
            .I(N__11774));
    LocalMux I__1873 (
            .O(N__11774),
            .I(N__11771));
    Odrv12 I__1872 (
            .O(N__11771),
            .I(\c0.tx_data_RNO_0Z0Z_0 ));
    InMux I__1871 (
            .O(N__11768),
            .I(N__11765));
    LocalMux I__1870 (
            .O(N__11765),
            .I(\c0.N_93 ));
    CascadeMux I__1869 (
            .O(N__11762),
            .I(N__11759));
    InMux I__1868 (
            .O(N__11759),
            .I(N__11756));
    LocalMux I__1867 (
            .O(N__11756),
            .I(N__11753));
    Odrv4 I__1866 (
            .O(N__11753),
            .I(\c0.nextCRC16_3_0_a2_0_10 ));
    InMux I__1865 (
            .O(N__11750),
            .I(N__11743));
    InMux I__1864 (
            .O(N__11749),
            .I(N__11743));
    CascadeMux I__1863 (
            .O(N__11748),
            .I(N__11740));
    LocalMux I__1862 (
            .O(N__11743),
            .I(N__11736));
    InMux I__1861 (
            .O(N__11740),
            .I(N__11731));
    InMux I__1860 (
            .O(N__11739),
            .I(N__11731));
    Span4Mux_h I__1859 (
            .O(N__11736),
            .I(N__11728));
    LocalMux I__1858 (
            .O(N__11731),
            .I(\c0.d_2_22 ));
    Odrv4 I__1857 (
            .O(N__11728),
            .I(\c0.d_2_22 ));
    InMux I__1856 (
            .O(N__11723),
            .I(N__11720));
    LocalMux I__1855 (
            .O(N__11720),
            .I(N__11717));
    Span4Mux_v I__1854 (
            .O(N__11717),
            .I(N__11713));
    InMux I__1853 (
            .O(N__11716),
            .I(N__11710));
    Span4Mux_h I__1852 (
            .O(N__11713),
            .I(N__11704));
    LocalMux I__1851 (
            .O(N__11710),
            .I(N__11704));
    InMux I__1850 (
            .O(N__11709),
            .I(N__11700));
    Span4Mux_v I__1849 (
            .O(N__11704),
            .I(N__11697));
    InMux I__1848 (
            .O(N__11703),
            .I(N__11694));
    LocalMux I__1847 (
            .O(N__11700),
            .I(\c0.d_2_6 ));
    Odrv4 I__1846 (
            .O(N__11697),
            .I(\c0.d_2_6 ));
    LocalMux I__1845 (
            .O(N__11694),
            .I(\c0.d_2_6 ));
    InMux I__1844 (
            .O(N__11687),
            .I(N__11684));
    LocalMux I__1843 (
            .O(N__11684),
            .I(N__11681));
    Odrv12 I__1842 (
            .O(N__11681),
            .I(\c0.nextCRC16_3_9 ));
    CascadeMux I__1841 (
            .O(N__11678),
            .I(\c0.nextCRC16_3_0_a2_6_0_15_cascade_ ));
    InMux I__1840 (
            .O(N__11675),
            .I(N__11672));
    LocalMux I__1839 (
            .O(N__11672),
            .I(N__11668));
    InMux I__1838 (
            .O(N__11671),
            .I(N__11665));
    Span4Mux_v I__1837 (
            .O(N__11668),
            .I(N__11660));
    LocalMux I__1836 (
            .O(N__11665),
            .I(N__11660));
    Odrv4 I__1835 (
            .O(N__11660),
            .I(\c0.N_92 ));
    InMux I__1834 (
            .O(N__11657),
            .I(\c0.tx2.r_Clock_Count12 ));
    InMux I__1833 (
            .O(N__11654),
            .I(N__11650));
    CascadeMux I__1832 (
            .O(N__11653),
            .I(N__11646));
    LocalMux I__1831 (
            .O(N__11650),
            .I(N__11643));
    InMux I__1830 (
            .O(N__11649),
            .I(N__11640));
    InMux I__1829 (
            .O(N__11646),
            .I(N__11637));
    Span4Mux_h I__1828 (
            .O(N__11643),
            .I(N__11634));
    LocalMux I__1827 (
            .O(N__11640),
            .I(N__11631));
    LocalMux I__1826 (
            .O(N__11637),
            .I(\c0.N_76 ));
    Odrv4 I__1825 (
            .O(N__11634),
            .I(\c0.N_76 ));
    Odrv12 I__1824 (
            .O(N__11631),
            .I(\c0.N_76 ));
    CascadeMux I__1823 (
            .O(N__11624),
            .I(N__11621));
    InMux I__1822 (
            .O(N__11621),
            .I(N__11618));
    LocalMux I__1821 (
            .O(N__11618),
            .I(\c0.data_out_6_Z0Z_2 ));
    InMux I__1820 (
            .O(N__11615),
            .I(N__11612));
    LocalMux I__1819 (
            .O(N__11612),
            .I(\c0.tx_data_RNO_0Z0Z_2 ));
    InMux I__1818 (
            .O(N__11609),
            .I(N__11606));
    LocalMux I__1817 (
            .O(N__11606),
            .I(N__11601));
    InMux I__1816 (
            .O(N__11605),
            .I(N__11598));
    InMux I__1815 (
            .O(N__11604),
            .I(N__11595));
    Span4Mux_v I__1814 (
            .O(N__11601),
            .I(N__11588));
    LocalMux I__1813 (
            .O(N__11598),
            .I(N__11588));
    LocalMux I__1812 (
            .O(N__11595),
            .I(N__11588));
    Span4Mux_h I__1811 (
            .O(N__11588),
            .I(N__11584));
    InMux I__1810 (
            .O(N__11587),
            .I(N__11581));
    Odrv4 I__1809 (
            .O(N__11584),
            .I(\c0.d_2_21 ));
    LocalMux I__1808 (
            .O(N__11581),
            .I(\c0.d_2_21 ));
    CascadeMux I__1807 (
            .O(N__11576),
            .I(\c0.tx_data_1_iv_i_m2_0_ns_1_0_cascade_ ));
    CascadeMux I__1806 (
            .O(N__11573),
            .I(\c0.N_304_cascade_ ));
    InMux I__1805 (
            .O(N__11570),
            .I(N__11567));
    LocalMux I__1804 (
            .O(N__11567),
            .I(N__11564));
    Span4Mux_h I__1803 (
            .O(N__11564),
            .I(N__11561));
    Odrv4 I__1802 (
            .O(N__11561),
            .I(\c0.tx_data_1_iv_i_1_0 ));
    InMux I__1801 (
            .O(N__11558),
            .I(\c0.tx2.un1_r_Clock_Count_cry_2 ));
    InMux I__1800 (
            .O(N__11555),
            .I(N__11552));
    LocalMux I__1799 (
            .O(N__11552),
            .I(\c0.tx2.r_Clock_Count_RNO_0_0_3 ));
    CascadeMux I__1798 (
            .O(N__11549),
            .I(N__11545));
    InMux I__1797 (
            .O(N__11548),
            .I(N__11542));
    InMux I__1796 (
            .O(N__11545),
            .I(N__11539));
    LocalMux I__1795 (
            .O(N__11542),
            .I(\c0.tx2.r_Clock_Count_0_sqmuxa ));
    LocalMux I__1794 (
            .O(N__11539),
            .I(\c0.tx2.r_Clock_Count_0_sqmuxa ));
    InMux I__1793 (
            .O(N__11534),
            .I(N__11531));
    LocalMux I__1792 (
            .O(N__11531),
            .I(\c0.tx2.r_Clock_Count_RNO_0_0_0 ));
    InMux I__1791 (
            .O(N__11528),
            .I(N__11524));
    InMux I__1790 (
            .O(N__11527),
            .I(N__11521));
    LocalMux I__1789 (
            .O(N__11524),
            .I(\c0.tx2.r_Clock_CountZ0Z_0 ));
    LocalMux I__1788 (
            .O(N__11521),
            .I(\c0.tx2.r_Clock_CountZ0Z_0 ));
    InMux I__1787 (
            .O(N__11516),
            .I(N__11513));
    LocalMux I__1786 (
            .O(N__11513),
            .I(\c0.tx2.r_Clock_Count_RNO_0_0_1 ));
    InMux I__1785 (
            .O(N__11510),
            .I(N__11506));
    InMux I__1784 (
            .O(N__11509),
            .I(N__11503));
    LocalMux I__1783 (
            .O(N__11506),
            .I(\c0.tx2.r_Clock_Count_i_0 ));
    LocalMux I__1782 (
            .O(N__11503),
            .I(\c0.tx2.r_Clock_Count_i_0 ));
    InMux I__1781 (
            .O(N__11498),
            .I(N__11494));
    InMux I__1780 (
            .O(N__11497),
            .I(N__11491));
    LocalMux I__1779 (
            .O(N__11494),
            .I(\c0.tx2.r_Clock_CountZ0Z_1 ));
    LocalMux I__1778 (
            .O(N__11491),
            .I(\c0.tx2.r_Clock_CountZ0Z_1 ));
    InMux I__1777 (
            .O(N__11486),
            .I(N__11483));
    LocalMux I__1776 (
            .O(N__11483),
            .I(\c0.tx2.r_Clock_Count_i_1 ));
    InMux I__1775 (
            .O(N__11480),
            .I(N__11476));
    InMux I__1774 (
            .O(N__11479),
            .I(N__11473));
    LocalMux I__1773 (
            .O(N__11476),
            .I(\c0.tx2.r_Clock_CountZ0Z_2 ));
    LocalMux I__1772 (
            .O(N__11473),
            .I(\c0.tx2.r_Clock_CountZ0Z_2 ));
    InMux I__1771 (
            .O(N__11468),
            .I(N__11465));
    LocalMux I__1770 (
            .O(N__11465),
            .I(\c0.tx2.r_Clock_Count_i_2 ));
    InMux I__1769 (
            .O(N__11462),
            .I(N__11458));
    InMux I__1768 (
            .O(N__11461),
            .I(N__11455));
    LocalMux I__1767 (
            .O(N__11458),
            .I(\c0.tx2.r_Clock_CountZ0Z_3 ));
    LocalMux I__1766 (
            .O(N__11455),
            .I(\c0.tx2.r_Clock_CountZ0Z_3 ));
    InMux I__1765 (
            .O(N__11450),
            .I(N__11447));
    LocalMux I__1764 (
            .O(N__11447),
            .I(\c0.tx2.r_Clock_Count_i_3 ));
    InMux I__1763 (
            .O(N__11444),
            .I(N__11440));
    InMux I__1762 (
            .O(N__11443),
            .I(N__11437));
    LocalMux I__1761 (
            .O(N__11440),
            .I(N__11433));
    LocalMux I__1760 (
            .O(N__11437),
            .I(N__11430));
    InMux I__1759 (
            .O(N__11436),
            .I(N__11427));
    Odrv12 I__1758 (
            .O(N__11433),
            .I(\c0.data_in_3_Z0Z_4 ));
    Odrv4 I__1757 (
            .O(N__11430),
            .I(\c0.data_in_3_Z0Z_4 ));
    LocalMux I__1756 (
            .O(N__11427),
            .I(\c0.data_in_3_Z0Z_4 ));
    InMux I__1755 (
            .O(N__11420),
            .I(N__11415));
    InMux I__1754 (
            .O(N__11419),
            .I(N__11412));
    InMux I__1753 (
            .O(N__11418),
            .I(N__11409));
    LocalMux I__1752 (
            .O(N__11415),
            .I(N__11406));
    LocalMux I__1751 (
            .O(N__11412),
            .I(N__11403));
    LocalMux I__1750 (
            .O(N__11409),
            .I(\c0.data_in_1_Z0Z_6 ));
    Odrv12 I__1749 (
            .O(N__11406),
            .I(\c0.data_in_1_Z0Z_6 ));
    Odrv4 I__1748 (
            .O(N__11403),
            .I(\c0.data_in_1_Z0Z_6 ));
    InMux I__1747 (
            .O(N__11396),
            .I(N__11392));
    InMux I__1746 (
            .O(N__11395),
            .I(N__11389));
    LocalMux I__1745 (
            .O(N__11392),
            .I(N__11385));
    LocalMux I__1744 (
            .O(N__11389),
            .I(N__11382));
    InMux I__1743 (
            .O(N__11388),
            .I(N__11379));
    Odrv4 I__1742 (
            .O(N__11385),
            .I(\c0.data_in_3_Z0Z_5 ));
    Odrv12 I__1741 (
            .O(N__11382),
            .I(\c0.data_in_3_Z0Z_5 ));
    LocalMux I__1740 (
            .O(N__11379),
            .I(\c0.data_in_3_Z0Z_5 ));
    InMux I__1739 (
            .O(N__11372),
            .I(N__11368));
    InMux I__1738 (
            .O(N__11371),
            .I(N__11365));
    LocalMux I__1737 (
            .O(N__11368),
            .I(\c0.data_in_5_Z0Z_2 ));
    LocalMux I__1736 (
            .O(N__11365),
            .I(\c0.data_in_5_Z0Z_2 ));
    InMux I__1735 (
            .O(N__11360),
            .I(\c0.tx2.un1_r_Clock_Count_cry_0 ));
    InMux I__1734 (
            .O(N__11357),
            .I(N__11354));
    LocalMux I__1733 (
            .O(N__11354),
            .I(\c0.tx2.r_Clock_Count_RNO_0_0_2 ));
    InMux I__1732 (
            .O(N__11351),
            .I(\c0.tx2.un1_r_Clock_Count_cry_1 ));
    CascadeMux I__1731 (
            .O(N__11348),
            .I(\c0.g3_2_0_cascade_ ));
    InMux I__1730 (
            .O(N__11345),
            .I(N__11342));
    LocalMux I__1729 (
            .O(N__11342),
            .I(\c0.g0_2 ));
    InMux I__1728 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1727 (
            .O(N__11336),
            .I(N__11333));
    Span4Mux_h I__1726 (
            .O(N__11333),
            .I(N__11329));
    InMux I__1725 (
            .O(N__11332),
            .I(N__11326));
    Odrv4 I__1724 (
            .O(N__11329),
            .I(\c0.rx_data_1 ));
    LocalMux I__1723 (
            .O(N__11326),
            .I(\c0.rx_data_1 ));
    InMux I__1722 (
            .O(N__11321),
            .I(N__11317));
    InMux I__1721 (
            .O(N__11320),
            .I(N__11314));
    LocalMux I__1720 (
            .O(N__11317),
            .I(\c0.data_in_4_Z0Z_0 ));
    LocalMux I__1719 (
            .O(N__11314),
            .I(\c0.data_in_4_Z0Z_0 ));
    CascadeMux I__1718 (
            .O(N__11309),
            .I(\c0.g1_cascade_ ));
    InMux I__1717 (
            .O(N__11306),
            .I(N__11303));
    LocalMux I__1716 (
            .O(N__11303),
            .I(\c0.g0_3 ));
    InMux I__1715 (
            .O(N__11300),
            .I(N__11297));
    LocalMux I__1714 (
            .O(N__11297),
            .I(\c0.byte_transmit_counter2_0_sqmuxa_0 ));
    CascadeMux I__1713 (
            .O(N__11294),
            .I(\c0.g1_1_cascade_ ));
    InMux I__1712 (
            .O(N__11291),
            .I(N__11288));
    LocalMux I__1711 (
            .O(N__11288),
            .I(\c0.N_72_mux ));
    CascadeMux I__1710 (
            .O(N__11285),
            .I(\c0.N_249_cascade_ ));
    InMux I__1709 (
            .O(N__11282),
            .I(N__11278));
    InMux I__1708 (
            .O(N__11281),
            .I(N__11275));
    LocalMux I__1707 (
            .O(N__11278),
            .I(\c0.dataZ0Z_5 ));
    LocalMux I__1706 (
            .O(N__11275),
            .I(\c0.dataZ0Z_5 ));
    InMux I__1705 (
            .O(N__11270),
            .I(N__11266));
    InMux I__1704 (
            .O(N__11269),
            .I(N__11263));
    LocalMux I__1703 (
            .O(N__11266),
            .I(\c0.dataZ0Z_13 ));
    LocalMux I__1702 (
            .O(N__11263),
            .I(\c0.dataZ0Z_13 ));
    InMux I__1701 (
            .O(N__11258),
            .I(N__11253));
    InMux I__1700 (
            .O(N__11257),
            .I(N__11250));
    InMux I__1699 (
            .O(N__11256),
            .I(N__11246));
    LocalMux I__1698 (
            .O(N__11253),
            .I(N__11241));
    LocalMux I__1697 (
            .O(N__11250),
            .I(N__11241));
    InMux I__1696 (
            .O(N__11249),
            .I(N__11238));
    LocalMux I__1695 (
            .O(N__11246),
            .I(N__11235));
    Span4Mux_h I__1694 (
            .O(N__11241),
            .I(N__11232));
    LocalMux I__1693 (
            .O(N__11238),
            .I(N__11229));
    Odrv12 I__1692 (
            .O(N__11235),
            .I(\c0.d_2_37 ));
    Odrv4 I__1691 (
            .O(N__11232),
            .I(\c0.d_2_37 ));
    Odrv4 I__1690 (
            .O(N__11229),
            .I(\c0.d_2_37 ));
    InMux I__1689 (
            .O(N__11222),
            .I(N__11218));
    InMux I__1688 (
            .O(N__11221),
            .I(N__11215));
    LocalMux I__1687 (
            .O(N__11218),
            .I(\c0.dataZ0Z_4 ));
    LocalMux I__1686 (
            .O(N__11215),
            .I(\c0.dataZ0Z_4 ));
    InMux I__1685 (
            .O(N__11210),
            .I(N__11206));
    InMux I__1684 (
            .O(N__11209),
            .I(N__11203));
    LocalMux I__1683 (
            .O(N__11206),
            .I(\c0.dataZ0Z_9 ));
    LocalMux I__1682 (
            .O(N__11203),
            .I(\c0.dataZ0Z_9 ));
    CascadeMux I__1681 (
            .O(N__11198),
            .I(N__11195));
    InMux I__1680 (
            .O(N__11195),
            .I(N__11192));
    LocalMux I__1679 (
            .O(N__11192),
            .I(\c0.i12_7_and ));
    CascadeMux I__1678 (
            .O(N__11189),
            .I(\c0.tx_data_RNO_3Z0Z_4_cascade_ ));
    InMux I__1677 (
            .O(N__11186),
            .I(N__11183));
    LocalMux I__1676 (
            .O(N__11183),
            .I(N__11180));
    Odrv4 I__1675 (
            .O(N__11180),
            .I(\c0.tx_data_1_0_i_ns_1_4 ));
    InMux I__1674 (
            .O(N__11177),
            .I(N__11174));
    LocalMux I__1673 (
            .O(N__11174),
            .I(\c0.tx_data_RNO_4Z0Z_4 ));
    InMux I__1672 (
            .O(N__11171),
            .I(N__11168));
    LocalMux I__1671 (
            .O(N__11168),
            .I(N__11165));
    Odrv4 I__1670 (
            .O(N__11165),
            .I(\c0.data_out_7_Z0Z_4 ));
    InMux I__1669 (
            .O(N__11162),
            .I(N__11158));
    InMux I__1668 (
            .O(N__11161),
            .I(N__11155));
    LocalMux I__1667 (
            .O(N__11158),
            .I(\c0.dataZ0Z_7 ));
    LocalMux I__1666 (
            .O(N__11155),
            .I(\c0.dataZ0Z_7 ));
    InMux I__1665 (
            .O(N__11150),
            .I(N__11146));
    InMux I__1664 (
            .O(N__11149),
            .I(N__11143));
    LocalMux I__1663 (
            .O(N__11146),
            .I(\c0.dataZ0Z_3 ));
    LocalMux I__1662 (
            .O(N__11143),
            .I(\c0.dataZ0Z_3 ));
    InMux I__1661 (
            .O(N__11138),
            .I(N__11134));
    InMux I__1660 (
            .O(N__11137),
            .I(N__11131));
    LocalMux I__1659 (
            .O(N__11134),
            .I(\c0.dataZ0Z_10 ));
    LocalMux I__1658 (
            .O(N__11131),
            .I(\c0.dataZ0Z_10 ));
    InMux I__1657 (
            .O(N__11126),
            .I(N__11122));
    InMux I__1656 (
            .O(N__11125),
            .I(N__11119));
    LocalMux I__1655 (
            .O(N__11122),
            .I(\c0.dataZ0Z_6 ));
    LocalMux I__1654 (
            .O(N__11119),
            .I(\c0.dataZ0Z_6 ));
    InMux I__1653 (
            .O(N__11114),
            .I(N__11110));
    InMux I__1652 (
            .O(N__11113),
            .I(N__11107));
    LocalMux I__1651 (
            .O(N__11110),
            .I(\c0.dataZ0Z_2 ));
    LocalMux I__1650 (
            .O(N__11107),
            .I(\c0.dataZ0Z_2 ));
    InMux I__1649 (
            .O(N__11102),
            .I(N__11099));
    LocalMux I__1648 (
            .O(N__11099),
            .I(N__11096));
    Span4Mux_v I__1647 (
            .O(N__11096),
            .I(N__11093));
    Odrv4 I__1646 (
            .O(N__11093),
            .I(\c0.data_out_7_Z0Z_2 ));
    InMux I__1645 (
            .O(N__11090),
            .I(N__11087));
    LocalMux I__1644 (
            .O(N__11087),
            .I(N__11084));
    Span4Mux_h I__1643 (
            .O(N__11084),
            .I(N__11081));
    Odrv4 I__1642 (
            .O(N__11081),
            .I(\c0.tx_data_RNO_0Z0Z_5 ));
    InMux I__1641 (
            .O(N__11078),
            .I(N__11071));
    InMux I__1640 (
            .O(N__11077),
            .I(N__11071));
    InMux I__1639 (
            .O(N__11076),
            .I(N__11068));
    LocalMux I__1638 (
            .O(N__11071),
            .I(N__11065));
    LocalMux I__1637 (
            .O(N__11068),
            .I(N__11059));
    Span4Mux_h I__1636 (
            .O(N__11065),
            .I(N__11059));
    CascadeMux I__1635 (
            .O(N__11064),
            .I(N__11056));
    Span4Mux_h I__1634 (
            .O(N__11059),
            .I(N__11053));
    InMux I__1633 (
            .O(N__11056),
            .I(N__11050));
    Odrv4 I__1632 (
            .O(N__11053),
            .I(\c0.d_2_23 ));
    LocalMux I__1631 (
            .O(N__11050),
            .I(\c0.d_2_23 ));
    InMux I__1630 (
            .O(N__11045),
            .I(N__11042));
    LocalMux I__1629 (
            .O(N__11042),
            .I(\c0.tx_data_RNO_0Z0Z_7 ));
    CascadeMux I__1628 (
            .O(N__11039),
            .I(N__11036));
    InMux I__1627 (
            .O(N__11036),
            .I(N__11033));
    LocalMux I__1626 (
            .O(N__11033),
            .I(N__11030));
    Span4Mux_h I__1625 (
            .O(N__11030),
            .I(N__11027));
    Span4Mux_h I__1624 (
            .O(N__11027),
            .I(N__11024));
    Odrv4 I__1623 (
            .O(N__11024),
            .I(\c0.tx_data_RNO_1Z0Z_1 ));
    CascadeMux I__1622 (
            .O(N__11021),
            .I(N__11018));
    InMux I__1621 (
            .O(N__11018),
            .I(N__11015));
    LocalMux I__1620 (
            .O(N__11015),
            .I(\c0.tx_data_RNO_1Z0Z_2 ));
    CascadeMux I__1619 (
            .O(N__11012),
            .I(\c0.nextCRC16_3_0_a2_1_15_cascade_ ));
    InMux I__1618 (
            .O(N__11009),
            .I(N__11006));
    LocalMux I__1617 (
            .O(N__11006),
            .I(N__11003));
    Odrv4 I__1616 (
            .O(N__11003),
            .I(\c0.m115_amcf1 ));
    CascadeMux I__1615 (
            .O(N__11000),
            .I(\c0.N_293_cascade_ ));
    InMux I__1614 (
            .O(N__10997),
            .I(N__10994));
    LocalMux I__1613 (
            .O(N__10994),
            .I(N__10991));
    Odrv4 I__1612 (
            .O(N__10991),
            .I(\c0.tx_data_1_0_i_1_6 ));
    CascadeMux I__1611 (
            .O(N__10988),
            .I(\c0.tx_data_RNO_1Z0Z_6_cascade_ ));
    InMux I__1610 (
            .O(N__10985),
            .I(N__10982));
    LocalMux I__1609 (
            .O(N__10982),
            .I(N__10979));
    Span4Mux_h I__1608 (
            .O(N__10979),
            .I(N__10976));
    Odrv4 I__1607 (
            .O(N__10976),
            .I(\c0.tx.r_Tx_DataZ0Z_6 ));
    InMux I__1606 (
            .O(N__10973),
            .I(N__10970));
    LocalMux I__1605 (
            .O(N__10970),
            .I(N__10967));
    Span4Mux_h I__1604 (
            .O(N__10967),
            .I(N__10964));
    Odrv4 I__1603 (
            .O(N__10964),
            .I(\c0.tx.r_Tx_DataZ0Z_2 ));
    InMux I__1602 (
            .O(N__10961),
            .I(N__10958));
    LocalMux I__1601 (
            .O(N__10958),
            .I(\c0.tx_data_1_0_i_ns_1_7 ));
    InMux I__1600 (
            .O(N__10955),
            .I(N__10952));
    LocalMux I__1599 (
            .O(N__10952),
            .I(N__10949));
    Span4Mux_h I__1598 (
            .O(N__10949),
            .I(N__10946));
    Odrv4 I__1597 (
            .O(N__10946),
            .I(\c0.tx.r_Tx_DataZ0Z_7 ));
    CEMux I__1596 (
            .O(N__10943),
            .I(N__10937));
    CEMux I__1595 (
            .O(N__10942),
            .I(N__10934));
    CEMux I__1594 (
            .O(N__10941),
            .I(N__10931));
    CascadeMux I__1593 (
            .O(N__10940),
            .I(N__10928));
    LocalMux I__1592 (
            .O(N__10937),
            .I(N__10925));
    LocalMux I__1591 (
            .O(N__10934),
            .I(N__10922));
    LocalMux I__1590 (
            .O(N__10931),
            .I(N__10918));
    InMux I__1589 (
            .O(N__10928),
            .I(N__10915));
    Span4Mux_h I__1588 (
            .O(N__10925),
            .I(N__10912));
    Span4Mux_h I__1587 (
            .O(N__10922),
            .I(N__10909));
    InMux I__1586 (
            .O(N__10921),
            .I(N__10906));
    Span4Mux_v I__1585 (
            .O(N__10918),
            .I(N__10901));
    LocalMux I__1584 (
            .O(N__10915),
            .I(N__10901));
    Span4Mux_h I__1583 (
            .O(N__10912),
            .I(N__10898));
    Span4Mux_h I__1582 (
            .O(N__10909),
            .I(N__10895));
    LocalMux I__1581 (
            .O(N__10906),
            .I(N__10892));
    Span4Mux_h I__1580 (
            .O(N__10901),
            .I(N__10889));
    Odrv4 I__1579 (
            .O(N__10898),
            .I(\c0.tx.r_Tx_Data_0_sqmuxa ));
    Odrv4 I__1578 (
            .O(N__10895),
            .I(\c0.tx.r_Tx_Data_0_sqmuxa ));
    Odrv12 I__1577 (
            .O(N__10892),
            .I(\c0.tx.r_Tx_Data_0_sqmuxa ));
    Odrv4 I__1576 (
            .O(N__10889),
            .I(\c0.tx.r_Tx_Data_0_sqmuxa ));
    CascadeMux I__1575 (
            .O(N__10880),
            .I(N__10877));
    InMux I__1574 (
            .O(N__10877),
            .I(N__10874));
    LocalMux I__1573 (
            .O(N__10874),
            .I(N__10871));
    Span4Mux_h I__1572 (
            .O(N__10871),
            .I(N__10868));
    Odrv4 I__1571 (
            .O(N__10868),
            .I(\c0.tx_data_RNO_1Z0Z_4 ));
    CascadeMux I__1570 (
            .O(N__10865),
            .I(N__10862));
    InMux I__1569 (
            .O(N__10862),
            .I(N__10859));
    LocalMux I__1568 (
            .O(N__10859),
            .I(N__10856));
    Span4Mux_v I__1567 (
            .O(N__10856),
            .I(N__10853));
    Odrv4 I__1566 (
            .O(N__10853),
            .I(\c0.data_out_6_Z0Z_1 ));
    CascadeMux I__1565 (
            .O(N__10850),
            .I(N__10846));
    InMux I__1564 (
            .O(N__10849),
            .I(N__10843));
    InMux I__1563 (
            .O(N__10846),
            .I(N__10840));
    LocalMux I__1562 (
            .O(N__10843),
            .I(N__10837));
    LocalMux I__1561 (
            .O(N__10840),
            .I(N__10834));
    Odrv12 I__1560 (
            .O(N__10837),
            .I(\c0.rx.un1_r_Rx_Byte_7 ));
    Odrv4 I__1559 (
            .O(N__10834),
            .I(\c0.rx.un1_r_Rx_Byte_7 ));
    CascadeMux I__1558 (
            .O(N__10829),
            .I(\c0.tx2.o_Tx_Serial12_cascade_ ));
    InMux I__1557 (
            .O(N__10826),
            .I(N__10823));
    LocalMux I__1556 (
            .O(N__10823),
            .I(N__10820));
    Span4Mux_h I__1555 (
            .O(N__10820),
            .I(N__10817));
    Odrv4 I__1554 (
            .O(N__10817),
            .I(\c0.tx_data_RNO_3Z0Z_3 ));
    InMux I__1553 (
            .O(N__10814),
            .I(N__10808));
    InMux I__1552 (
            .O(N__10813),
            .I(N__10805));
    InMux I__1551 (
            .O(N__10812),
            .I(N__10802));
    InMux I__1550 (
            .O(N__10811),
            .I(N__10799));
    LocalMux I__1549 (
            .O(N__10808),
            .I(N__10796));
    LocalMux I__1548 (
            .O(N__10805),
            .I(\c0.d_2_38 ));
    LocalMux I__1547 (
            .O(N__10802),
            .I(\c0.d_2_38 ));
    LocalMux I__1546 (
            .O(N__10799),
            .I(\c0.d_2_38 ));
    Odrv4 I__1545 (
            .O(N__10796),
            .I(\c0.d_2_38 ));
    InMux I__1544 (
            .O(N__10787),
            .I(N__10784));
    LocalMux I__1543 (
            .O(N__10784),
            .I(N__10780));
    InMux I__1542 (
            .O(N__10783),
            .I(N__10777));
    Odrv12 I__1541 (
            .O(N__10780),
            .I(\c0.rx_data_5 ));
    LocalMux I__1540 (
            .O(N__10777),
            .I(\c0.rx_data_5 ));
    InMux I__1539 (
            .O(N__10772),
            .I(N__10769));
    LocalMux I__1538 (
            .O(N__10769),
            .I(\c0.tx2_data_RNO_4Z0Z_2 ));
    InMux I__1537 (
            .O(N__10766),
            .I(N__10763));
    LocalMux I__1536 (
            .O(N__10763),
            .I(\c0.tx2_data_RNO_1Z0Z_2 ));
    CascadeMux I__1535 (
            .O(N__10760),
            .I(\c0.tx2_data_RNO_0Z0Z_2_cascade_ ));
    InMux I__1534 (
            .O(N__10757),
            .I(N__10754));
    LocalMux I__1533 (
            .O(N__10754),
            .I(\c0.tx2_data_1_0_i_ns_1_2 ));
    InMux I__1532 (
            .O(N__10751),
            .I(N__10748));
    LocalMux I__1531 (
            .O(N__10748),
            .I(N__10745));
    Odrv4 I__1530 (
            .O(N__10745),
            .I(\c0.tx2_data_1_iv_4_3 ));
    CascadeMux I__1529 (
            .O(N__10742),
            .I(N__10739));
    InMux I__1528 (
            .O(N__10739),
            .I(N__10736));
    LocalMux I__1527 (
            .O(N__10736),
            .I(\c0.i12_4_and ));
    CascadeMux I__1526 (
            .O(N__10733),
            .I(N__10730));
    InMux I__1525 (
            .O(N__10730),
            .I(N__10727));
    LocalMux I__1524 (
            .O(N__10727),
            .I(N__10724));
    Odrv4 I__1523 (
            .O(N__10724),
            .I(\c0.i12_6_and ));
    CascadeMux I__1522 (
            .O(N__10721),
            .I(N__10718));
    InMux I__1521 (
            .O(N__10718),
            .I(N__10715));
    LocalMux I__1520 (
            .O(N__10715),
            .I(\c0.i12_5_and ));
    InMux I__1519 (
            .O(N__10712),
            .I(bfn_10_18_0_));
    CascadeMux I__1518 (
            .O(N__10709),
            .I(N__10706));
    InMux I__1517 (
            .O(N__10706),
            .I(N__10703));
    LocalMux I__1516 (
            .O(N__10703),
            .I(\c0.i12_1_and ));
    CascadeMux I__1515 (
            .O(N__10700),
            .I(N__10697));
    InMux I__1514 (
            .O(N__10697),
            .I(N__10694));
    LocalMux I__1513 (
            .O(N__10694),
            .I(\c0.i12_3_and ));
    InMux I__1512 (
            .O(N__10691),
            .I(\c0.data_cry_13 ));
    InMux I__1511 (
            .O(N__10688),
            .I(\c0.data_cry_14 ));
    CascadeMux I__1510 (
            .O(N__10685),
            .I(N__10682));
    InMux I__1509 (
            .O(N__10682),
            .I(N__10679));
    LocalMux I__1508 (
            .O(N__10679),
            .I(\c0.i12_0_and ));
    CascadeMux I__1507 (
            .O(N__10676),
            .I(N__10673));
    InMux I__1506 (
            .O(N__10673),
            .I(N__10670));
    LocalMux I__1505 (
            .O(N__10670),
            .I(\c0.i12_2_and ));
    InMux I__1504 (
            .O(N__10667),
            .I(\c0.data_cry_5 ));
    InMux I__1503 (
            .O(N__10664),
            .I(\c0.data_cry_6 ));
    InMux I__1502 (
            .O(N__10661),
            .I(bfn_9_28_0_));
    InMux I__1501 (
            .O(N__10658),
            .I(\c0.data_cry_8 ));
    InMux I__1500 (
            .O(N__10655),
            .I(\c0.data_cry_9 ));
    InMux I__1499 (
            .O(N__10652),
            .I(N__10649));
    LocalMux I__1498 (
            .O(N__10649),
            .I(N__10646));
    Span4Mux_h I__1497 (
            .O(N__10646),
            .I(N__10642));
    InMux I__1496 (
            .O(N__10645),
            .I(N__10639));
    Odrv4 I__1495 (
            .O(N__10642),
            .I(\c0.dataZ0Z_11 ));
    LocalMux I__1494 (
            .O(N__10639),
            .I(\c0.dataZ0Z_11 ));
    InMux I__1493 (
            .O(N__10634),
            .I(\c0.data_cry_10 ));
    InMux I__1492 (
            .O(N__10631),
            .I(N__10628));
    LocalMux I__1491 (
            .O(N__10628),
            .I(N__10624));
    InMux I__1490 (
            .O(N__10627),
            .I(N__10621));
    Odrv4 I__1489 (
            .O(N__10624),
            .I(\c0.dataZ0Z_12 ));
    LocalMux I__1488 (
            .O(N__10621),
            .I(\c0.dataZ0Z_12 ));
    InMux I__1487 (
            .O(N__10616),
            .I(\c0.data_cry_11 ));
    InMux I__1486 (
            .O(N__10613),
            .I(\c0.data_cry_12 ));
    InMux I__1485 (
            .O(N__10610),
            .I(N__10607));
    LocalMux I__1484 (
            .O(N__10607),
            .I(N__10603));
    InMux I__1483 (
            .O(N__10606),
            .I(N__10600));
    Odrv12 I__1482 (
            .O(N__10603),
            .I(\c0.dataZ0Z_14 ));
    LocalMux I__1481 (
            .O(N__10600),
            .I(\c0.dataZ0Z_14 ));
    CascadeMux I__1480 (
            .O(N__10595),
            .I(\c0.N_74_cascade_ ));
    InMux I__1479 (
            .O(N__10592),
            .I(N__10588));
    InMux I__1478 (
            .O(N__10591),
            .I(N__10585));
    LocalMux I__1477 (
            .O(N__10588),
            .I(\c0.d_2_19 ));
    LocalMux I__1476 (
            .O(N__10585),
            .I(\c0.d_2_19 ));
    InMux I__1475 (
            .O(N__10580),
            .I(bfn_9_27_0_));
    InMux I__1474 (
            .O(N__10577),
            .I(N__10574));
    LocalMux I__1473 (
            .O(N__10574),
            .I(N__10570));
    InMux I__1472 (
            .O(N__10573),
            .I(N__10567));
    Odrv4 I__1471 (
            .O(N__10570),
            .I(\c0.dataZ0Z_1 ));
    LocalMux I__1470 (
            .O(N__10567),
            .I(\c0.dataZ0Z_1 ));
    InMux I__1469 (
            .O(N__10562),
            .I(\c0.data_cry_0 ));
    InMux I__1468 (
            .O(N__10559),
            .I(\c0.data_cry_1 ));
    InMux I__1467 (
            .O(N__10556),
            .I(\c0.data_cry_2 ));
    InMux I__1466 (
            .O(N__10553),
            .I(\c0.data_cry_3 ));
    InMux I__1465 (
            .O(N__10550),
            .I(\c0.data_cry_4 ));
    CascadeMux I__1464 (
            .O(N__10547),
            .I(\c0.tx_data_RNO_4Z0Z_1_cascade_ ));
    InMux I__1463 (
            .O(N__10544),
            .I(N__10541));
    LocalMux I__1462 (
            .O(N__10541),
            .I(N__10538));
    Odrv4 I__1461 (
            .O(N__10538),
            .I(\c0.tx_data_1_0_i_ns_1_1 ));
    InMux I__1460 (
            .O(N__10535),
            .I(N__10532));
    LocalMux I__1459 (
            .O(N__10532),
            .I(N__10529));
    Span4Mux_v I__1458 (
            .O(N__10529),
            .I(N__10526));
    Odrv4 I__1457 (
            .O(N__10526),
            .I(\c0.tx_data_RNO_0Z0Z_3 ));
    CascadeMux I__1456 (
            .O(N__10523),
            .I(\c0.nextCRC16_3_0_a2_1_11_cascade_ ));
    CascadeMux I__1455 (
            .O(N__10520),
            .I(N__10517));
    InMux I__1454 (
            .O(N__10517),
            .I(N__10514));
    LocalMux I__1453 (
            .O(N__10514),
            .I(\c0.data_out_6_Z0Z_3 ));
    InMux I__1452 (
            .O(N__10511),
            .I(N__10507));
    InMux I__1451 (
            .O(N__10510),
            .I(N__10504));
    LocalMux I__1450 (
            .O(N__10507),
            .I(N__10501));
    LocalMux I__1449 (
            .O(N__10504),
            .I(N__10498));
    Odrv12 I__1448 (
            .O(N__10501),
            .I(\c0.d_2_7 ));
    Odrv4 I__1447 (
            .O(N__10498),
            .I(\c0.d_2_7 ));
    CascadeMux I__1446 (
            .O(N__10493),
            .I(\c0.tx_data_RNO_3Z0Z_7_cascade_ ));
    InMux I__1445 (
            .O(N__10490),
            .I(N__10487));
    LocalMux I__1444 (
            .O(N__10487),
            .I(\c0.tx_data_RNO_4Z0Z_7 ));
    InMux I__1443 (
            .O(N__10484),
            .I(N__10481));
    LocalMux I__1442 (
            .O(N__10481),
            .I(N__10478));
    Span4Mux_h I__1441 (
            .O(N__10478),
            .I(N__10475));
    Odrv4 I__1440 (
            .O(N__10475),
            .I(\c0.N_74 ));
    InMux I__1439 (
            .O(N__10472),
            .I(N__10465));
    InMux I__1438 (
            .O(N__10471),
            .I(N__10462));
    InMux I__1437 (
            .O(N__10470),
            .I(N__10459));
    InMux I__1436 (
            .O(N__10469),
            .I(N__10454));
    InMux I__1435 (
            .O(N__10468),
            .I(N__10454));
    LocalMux I__1434 (
            .O(N__10465),
            .I(N__10450));
    LocalMux I__1433 (
            .O(N__10462),
            .I(N__10445));
    LocalMux I__1432 (
            .O(N__10459),
            .I(N__10445));
    LocalMux I__1431 (
            .O(N__10454),
            .I(N__10442));
    InMux I__1430 (
            .O(N__10453),
            .I(N__10436));
    Span4Mux_v I__1429 (
            .O(N__10450),
            .I(N__10431));
    Span4Mux_v I__1428 (
            .O(N__10445),
            .I(N__10431));
    Span4Mux_v I__1427 (
            .O(N__10442),
            .I(N__10428));
    InMux I__1426 (
            .O(N__10441),
            .I(N__10423));
    InMux I__1425 (
            .O(N__10440),
            .I(N__10423));
    InMux I__1424 (
            .O(N__10439),
            .I(N__10420));
    LocalMux I__1423 (
            .O(N__10436),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    Odrv4 I__1422 (
            .O(N__10431),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    Odrv4 I__1421 (
            .O(N__10428),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    LocalMux I__1420 (
            .O(N__10423),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    LocalMux I__1419 (
            .O(N__10420),
            .I(\c0.tx.r_SM_MainZ0Z_0 ));
    CascadeMux I__1418 (
            .O(N__10409),
            .I(N__10404));
    CascadeMux I__1417 (
            .O(N__10408),
            .I(N__10399));
    InMux I__1416 (
            .O(N__10407),
            .I(N__10394));
    InMux I__1415 (
            .O(N__10404),
            .I(N__10391));
    InMux I__1414 (
            .O(N__10403),
            .I(N__10388));
    InMux I__1413 (
            .O(N__10402),
            .I(N__10385));
    InMux I__1412 (
            .O(N__10399),
            .I(N__10382));
    InMux I__1411 (
            .O(N__10398),
            .I(N__10379));
    InMux I__1410 (
            .O(N__10397),
            .I(N__10375));
    LocalMux I__1409 (
            .O(N__10394),
            .I(N__10370));
    LocalMux I__1408 (
            .O(N__10391),
            .I(N__10370));
    LocalMux I__1407 (
            .O(N__10388),
            .I(N__10363));
    LocalMux I__1406 (
            .O(N__10385),
            .I(N__10363));
    LocalMux I__1405 (
            .O(N__10382),
            .I(N__10358));
    LocalMux I__1404 (
            .O(N__10379),
            .I(N__10358));
    InMux I__1403 (
            .O(N__10378),
            .I(N__10355));
    LocalMux I__1402 (
            .O(N__10375),
            .I(N__10350));
    Span4Mux_v I__1401 (
            .O(N__10370),
            .I(N__10350));
    InMux I__1400 (
            .O(N__10369),
            .I(N__10345));
    InMux I__1399 (
            .O(N__10368),
            .I(N__10345));
    Span4Mux_h I__1398 (
            .O(N__10363),
            .I(N__10342));
    Span4Mux_h I__1397 (
            .O(N__10358),
            .I(N__10339));
    LocalMux I__1396 (
            .O(N__10355),
            .I(\c0.tx.r_SM_MainZ0Z_1 ));
    Odrv4 I__1395 (
            .O(N__10350),
            .I(\c0.tx.r_SM_MainZ0Z_1 ));
    LocalMux I__1394 (
            .O(N__10345),
            .I(\c0.tx.r_SM_MainZ0Z_1 ));
    Odrv4 I__1393 (
            .O(N__10342),
            .I(\c0.tx.r_SM_MainZ0Z_1 ));
    Odrv4 I__1392 (
            .O(N__10339),
            .I(\c0.tx.r_SM_MainZ0Z_1 ));
    InMux I__1391 (
            .O(N__10328),
            .I(N__10324));
    InMux I__1390 (
            .O(N__10327),
            .I(N__10321));
    LocalMux I__1389 (
            .O(N__10324),
            .I(N__10313));
    LocalMux I__1388 (
            .O(N__10321),
            .I(N__10313));
    InMux I__1387 (
            .O(N__10320),
            .I(N__10310));
    InMux I__1386 (
            .O(N__10319),
            .I(N__10307));
    InMux I__1385 (
            .O(N__10318),
            .I(N__10297));
    Span4Mux_h I__1384 (
            .O(N__10313),
            .I(N__10294));
    LocalMux I__1383 (
            .O(N__10310),
            .I(N__10289));
    LocalMux I__1382 (
            .O(N__10307),
            .I(N__10289));
    InMux I__1381 (
            .O(N__10306),
            .I(N__10282));
    InMux I__1380 (
            .O(N__10305),
            .I(N__10282));
    InMux I__1379 (
            .O(N__10304),
            .I(N__10282));
    InMux I__1378 (
            .O(N__10303),
            .I(N__10273));
    InMux I__1377 (
            .O(N__10302),
            .I(N__10273));
    InMux I__1376 (
            .O(N__10301),
            .I(N__10273));
    InMux I__1375 (
            .O(N__10300),
            .I(N__10273));
    LocalMux I__1374 (
            .O(N__10297),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    Odrv4 I__1373 (
            .O(N__10294),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    Odrv4 I__1372 (
            .O(N__10289),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    LocalMux I__1371 (
            .O(N__10282),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    LocalMux I__1370 (
            .O(N__10273),
            .I(\c0.tx.r_Clock_Count12_THRU_CO ));
    CascadeMux I__1369 (
            .O(N__10262),
            .I(N__10256));
    InMux I__1368 (
            .O(N__10261),
            .I(N__10250));
    InMux I__1367 (
            .O(N__10260),
            .I(N__10247));
    CascadeMux I__1366 (
            .O(N__10259),
            .I(N__10241));
    InMux I__1365 (
            .O(N__10256),
            .I(N__10236));
    CascadeMux I__1364 (
            .O(N__10255),
            .I(N__10233));
    InMux I__1363 (
            .O(N__10254),
            .I(N__10228));
    InMux I__1362 (
            .O(N__10253),
            .I(N__10228));
    LocalMux I__1361 (
            .O(N__10250),
            .I(N__10225));
    LocalMux I__1360 (
            .O(N__10247),
            .I(N__10222));
    InMux I__1359 (
            .O(N__10246),
            .I(N__10213));
    InMux I__1358 (
            .O(N__10245),
            .I(N__10213));
    InMux I__1357 (
            .O(N__10244),
            .I(N__10213));
    InMux I__1356 (
            .O(N__10241),
            .I(N__10213));
    InMux I__1355 (
            .O(N__10240),
            .I(N__10210));
    CascadeMux I__1354 (
            .O(N__10239),
            .I(N__10206));
    LocalMux I__1353 (
            .O(N__10236),
            .I(N__10203));
    InMux I__1352 (
            .O(N__10233),
            .I(N__10200));
    LocalMux I__1351 (
            .O(N__10228),
            .I(N__10197));
    Span4Mux_h I__1350 (
            .O(N__10225),
            .I(N__10190));
    Span4Mux_v I__1349 (
            .O(N__10222),
            .I(N__10190));
    LocalMux I__1348 (
            .O(N__10213),
            .I(N__10190));
    LocalMux I__1347 (
            .O(N__10210),
            .I(N__10187));
    InMux I__1346 (
            .O(N__10209),
            .I(N__10182));
    InMux I__1345 (
            .O(N__10206),
            .I(N__10182));
    Span4Mux_v I__1344 (
            .O(N__10203),
            .I(N__10175));
    LocalMux I__1343 (
            .O(N__10200),
            .I(N__10175));
    Span4Mux_v I__1342 (
            .O(N__10197),
            .I(N__10175));
    Span4Mux_h I__1341 (
            .O(N__10190),
            .I(N__10172));
    Odrv4 I__1340 (
            .O(N__10187),
            .I(\c0.tx.r_SM_MainZ0Z_2 ));
    LocalMux I__1339 (
            .O(N__10182),
            .I(\c0.tx.r_SM_MainZ0Z_2 ));
    Odrv4 I__1338 (
            .O(N__10175),
            .I(\c0.tx.r_SM_MainZ0Z_2 ));
    Odrv4 I__1337 (
            .O(N__10172),
            .I(\c0.tx.r_SM_MainZ0Z_2 ));
    CascadeMux I__1336 (
            .O(N__10163),
            .I(\c0.nextCRC16_3_3_12_cascade_ ));
    InMux I__1335 (
            .O(N__10160),
            .I(N__10157));
    LocalMux I__1334 (
            .O(N__10157),
            .I(\c0.nextCRC16_3_4_12 ));
    InMux I__1333 (
            .O(N__10154),
            .I(N__10151));
    LocalMux I__1332 (
            .O(N__10151),
            .I(N__10148));
    Odrv4 I__1331 (
            .O(N__10148),
            .I(\c0.data_out_6_Z0Z_4 ));
    InMux I__1330 (
            .O(N__10145),
            .I(N__10142));
    LocalMux I__1329 (
            .O(N__10142),
            .I(N__10139));
    Span4Mux_v I__1328 (
            .O(N__10139),
            .I(N__10136));
    Odrv4 I__1327 (
            .O(N__10136),
            .I(\c0.tx_data_RNO_0Z0Z_4 ));
    CascadeMux I__1326 (
            .O(N__10133),
            .I(\c0.rx.r_Rx_Bytece_0_3_cascade_ ));
    InMux I__1325 (
            .O(N__10130),
            .I(N__10126));
    InMux I__1324 (
            .O(N__10129),
            .I(N__10123));
    LocalMux I__1323 (
            .O(N__10126),
            .I(\c0.rx_data_3 ));
    LocalMux I__1322 (
            .O(N__10123),
            .I(\c0.rx_data_3 ));
    CascadeMux I__1321 (
            .O(N__10118),
            .I(\c0.tx2_data_RNO_3Z0Z_2_cascade_ ));
    CascadeMux I__1320 (
            .O(N__10115),
            .I(\c0.tx_data_RNO_1Z0Z_0_cascade_ ));
    InMux I__1319 (
            .O(N__10112),
            .I(N__10109));
    LocalMux I__1318 (
            .O(N__10109),
            .I(N__10106));
    Odrv4 I__1317 (
            .O(N__10106),
            .I(\c0.tx.r_Tx_DataZ0Z_0 ));
    CascadeMux I__1316 (
            .O(N__10103),
            .I(N__10100));
    InMux I__1315 (
            .O(N__10100),
            .I(N__10097));
    LocalMux I__1314 (
            .O(N__10097),
            .I(\c0.tx.r_Tx_DataZ0Z_4 ));
    CascadeMux I__1313 (
            .O(N__10094),
            .I(N__10091));
    InMux I__1312 (
            .O(N__10091),
            .I(N__10088));
    LocalMux I__1311 (
            .O(N__10088),
            .I(N__10085));
    Span4Mux_h I__1310 (
            .O(N__10085),
            .I(N__10082));
    Odrv4 I__1309 (
            .O(N__10082),
            .I(\c0.data_out_7_Z0Z_5 ));
    CascadeMux I__1308 (
            .O(N__10079),
            .I(\c0.tx_data_1_0_i_ns_1_3_cascade_ ));
    InMux I__1307 (
            .O(N__10076),
            .I(N__10073));
    LocalMux I__1306 (
            .O(N__10073),
            .I(\c0.tx.r_Tx_DataZ0Z_3 ));
    CascadeMux I__1305 (
            .O(N__10070),
            .I(N__10067));
    InMux I__1304 (
            .O(N__10067),
            .I(N__10064));
    LocalMux I__1303 (
            .O(N__10064),
            .I(\c0.tx_data_RNO_1Z0Z_5 ));
    CascadeMux I__1302 (
            .O(N__10061),
            .I(N__10058));
    InMux I__1301 (
            .O(N__10058),
            .I(N__10055));
    LocalMux I__1300 (
            .O(N__10055),
            .I(\c0.tx.r_Tx_DataZ0Z_5 ));
    InMux I__1299 (
            .O(N__10052),
            .I(N__10049));
    LocalMux I__1298 (
            .O(N__10049),
            .I(\c0.tx_data_RNO_4Z0Z_3 ));
    InMux I__1297 (
            .O(N__10046),
            .I(N__10040));
    InMux I__1296 (
            .O(N__10045),
            .I(N__10037));
    InMux I__1295 (
            .O(N__10044),
            .I(N__10034));
    InMux I__1294 (
            .O(N__10043),
            .I(N__10031));
    LocalMux I__1293 (
            .O(N__10040),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__1292 (
            .O(N__10037),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__1291 (
            .O(N__10034),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    LocalMux I__1290 (
            .O(N__10031),
            .I(\c0.tx.r_Bit_IndexZ0Z_2 ));
    InMux I__1289 (
            .O(N__10022),
            .I(N__10012));
    InMux I__1288 (
            .O(N__10021),
            .I(N__10012));
    InMux I__1287 (
            .O(N__10020),
            .I(N__10007));
    InMux I__1286 (
            .O(N__10019),
            .I(N__10007));
    InMux I__1285 (
            .O(N__10018),
            .I(N__10002));
    InMux I__1284 (
            .O(N__10017),
            .I(N__10002));
    LocalMux I__1283 (
            .O(N__10012),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__1282 (
            .O(N__10007),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    LocalMux I__1281 (
            .O(N__10002),
            .I(\c0.tx.r_Bit_IndexZ0Z_1 ));
    CascadeMux I__1280 (
            .O(N__9995),
            .I(\c0.tx.r_Tx_Data_pmux_3_i_m2_ns_1_cascade_ ));
    InMux I__1279 (
            .O(N__9992),
            .I(N__9989));
    LocalMux I__1278 (
            .O(N__9989),
            .I(\c0.tx.N_354 ));
    CascadeMux I__1277 (
            .O(N__9986),
            .I(N__9982));
    InMux I__1276 (
            .O(N__9985),
            .I(N__9977));
    InMux I__1275 (
            .O(N__9982),
            .I(N__9974));
    InMux I__1274 (
            .O(N__9981),
            .I(N__9969));
    InMux I__1273 (
            .O(N__9980),
            .I(N__9969));
    LocalMux I__1272 (
            .O(N__9977),
            .I(N__9966));
    LocalMux I__1271 (
            .O(N__9974),
            .I(\c0.tx.r_Bit_IndexZ0Z_0 ));
    LocalMux I__1270 (
            .O(N__9969),
            .I(\c0.tx.r_Bit_IndexZ0Z_0 ));
    Odrv4 I__1269 (
            .O(N__9966),
            .I(\c0.tx.r_Bit_IndexZ0Z_0 ));
    CascadeMux I__1268 (
            .O(N__9959),
            .I(\c0.tx.N_357_cascade_ ));
    InMux I__1267 (
            .O(N__9956),
            .I(N__9953));
    LocalMux I__1266 (
            .O(N__9953),
            .I(N__9950));
    Odrv12 I__1265 (
            .O(N__9950),
            .I(\c0.tx.N_320 ));
    CascadeMux I__1264 (
            .O(N__9947),
            .I(\c0.tx_data_RNO_3Z0Z_5_cascade_ ));
    InMux I__1263 (
            .O(N__9944),
            .I(N__9941));
    LocalMux I__1262 (
            .O(N__9941),
            .I(\c0.tx_data_1_0_i_ns_1_5 ));
    InMux I__1261 (
            .O(N__9938),
            .I(N__9934));
    InMux I__1260 (
            .O(N__9937),
            .I(N__9931));
    LocalMux I__1259 (
            .O(N__9934),
            .I(N__9928));
    LocalMux I__1258 (
            .O(N__9931),
            .I(N__9925));
    Span4Mux_h I__1257 (
            .O(N__9928),
            .I(N__9919));
    Span4Mux_v I__1256 (
            .O(N__9925),
            .I(N__9919));
    InMux I__1255 (
            .O(N__9924),
            .I(N__9916));
    Odrv4 I__1254 (
            .O(N__9919),
            .I(\c0.rx.r_Rx_DV6 ));
    LocalMux I__1253 (
            .O(N__9916),
            .I(\c0.rx.r_Rx_DV6 ));
    CascadeMux I__1252 (
            .O(N__9911),
            .I(\c0.tx.r_Tx_Active_1_sqmuxa_cascade_ ));
    InMux I__1251 (
            .O(N__9908),
            .I(N__9905));
    LocalMux I__1250 (
            .O(N__9905),
            .I(\c0.tx_data_RNO_0Z0Z_1 ));
    InMux I__1249 (
            .O(N__9902),
            .I(N__9899));
    LocalMux I__1248 (
            .O(N__9899),
            .I(\c0.tx.r_Tx_DataZ0Z_1 ));
    CascadeMux I__1247 (
            .O(N__9896),
            .I(\c0.tx.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_ ));
    CascadeMux I__1246 (
            .O(N__9893),
            .I(\c0.rx.r_Rx_Bytece_1_1_cascade_ ));
    InMux I__1245 (
            .O(N__9890),
            .I(N__9887));
    LocalMux I__1244 (
            .O(N__9887),
            .I(\c0.rx.r_Rx_Bytece_1_5 ));
    InMux I__1243 (
            .O(N__9884),
            .I(N__9880));
    InMux I__1242 (
            .O(N__9883),
            .I(N__9877));
    LocalMux I__1241 (
            .O(N__9880),
            .I(\c0.tx.r_Clock_Count_i_0 ));
    LocalMux I__1240 (
            .O(N__9877),
            .I(\c0.tx.r_Clock_Count_i_0 ));
    InMux I__1239 (
            .O(N__9872),
            .I(N__9868));
    InMux I__1238 (
            .O(N__9871),
            .I(N__9865));
    LocalMux I__1237 (
            .O(N__9868),
            .I(\c0.tx.r_Clock_CountZ0Z_1 ));
    LocalMux I__1236 (
            .O(N__9865),
            .I(\c0.tx.r_Clock_CountZ0Z_1 ));
    InMux I__1235 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1234 (
            .O(N__9857),
            .I(\c0.tx.r_Clock_Count_i_1 ));
    InMux I__1233 (
            .O(N__9854),
            .I(N__9850));
    InMux I__1232 (
            .O(N__9853),
            .I(N__9847));
    LocalMux I__1231 (
            .O(N__9850),
            .I(\c0.tx.r_Clock_CountZ0Z_2 ));
    LocalMux I__1230 (
            .O(N__9847),
            .I(\c0.tx.r_Clock_CountZ0Z_2 ));
    InMux I__1229 (
            .O(N__9842),
            .I(N__9839));
    LocalMux I__1228 (
            .O(N__9839),
            .I(\c0.tx.r_Clock_Count_i_2 ));
    InMux I__1227 (
            .O(N__9836),
            .I(N__9832));
    InMux I__1226 (
            .O(N__9835),
            .I(N__9829));
    LocalMux I__1225 (
            .O(N__9832),
            .I(\c0.tx.r_Clock_CountZ0Z_3 ));
    LocalMux I__1224 (
            .O(N__9829),
            .I(\c0.tx.r_Clock_CountZ0Z_3 ));
    InMux I__1223 (
            .O(N__9824),
            .I(N__9821));
    LocalMux I__1222 (
            .O(N__9821),
            .I(\c0.tx.r_Clock_Count_i_3 ));
    InMux I__1221 (
            .O(N__9818),
            .I(\c0.tx.r_Clock_Count12 ));
    InMux I__1220 (
            .O(N__9815),
            .I(blink_counter_cry_24));
    InMux I__1219 (
            .O(N__9812),
            .I(N__9808));
    InMux I__1218 (
            .O(N__9811),
            .I(N__9805));
    LocalMux I__1217 (
            .O(N__9808),
            .I(N__9800));
    LocalMux I__1216 (
            .O(N__9805),
            .I(N__9800));
    Span4Mux_v I__1215 (
            .O(N__9800),
            .I(N__9796));
    InMux I__1214 (
            .O(N__9799),
            .I(N__9793));
    Odrv4 I__1213 (
            .O(N__9796),
            .I(blink_counterZ0Z_25));
    LocalMux I__1212 (
            .O(N__9793),
            .I(blink_counterZ0Z_25));
    CascadeMux I__1211 (
            .O(N__9788),
            .I(\c0.tx.N_287_cascade_ ));
    InMux I__1210 (
            .O(N__9785),
            .I(N__9782));
    LocalMux I__1209 (
            .O(N__9782),
            .I(\c0.tx.N_294 ));
    SRMux I__1208 (
            .O(N__9779),
            .I(N__9774));
    CascadeMux I__1207 (
            .O(N__9778),
            .I(N__9770));
    CascadeMux I__1206 (
            .O(N__9777),
            .I(N__9767));
    LocalMux I__1205 (
            .O(N__9774),
            .I(N__9763));
    InMux I__1204 (
            .O(N__9773),
            .I(N__9756));
    InMux I__1203 (
            .O(N__9770),
            .I(N__9756));
    InMux I__1202 (
            .O(N__9767),
            .I(N__9756));
    CascadeMux I__1201 (
            .O(N__9766),
            .I(N__9753));
    Span4Mux_v I__1200 (
            .O(N__9763),
            .I(N__9749));
    LocalMux I__1199 (
            .O(N__9756),
            .I(N__9746));
    InMux I__1198 (
            .O(N__9753),
            .I(N__9743));
    InMux I__1197 (
            .O(N__9752),
            .I(N__9740));
    Odrv4 I__1196 (
            .O(N__9749),
            .I(\c0.tx.o_Tx_Serial12 ));
    Odrv4 I__1195 (
            .O(N__9746),
            .I(\c0.tx.o_Tx_Serial12 ));
    LocalMux I__1194 (
            .O(N__9743),
            .I(\c0.tx.o_Tx_Serial12 ));
    LocalMux I__1193 (
            .O(N__9740),
            .I(\c0.tx.o_Tx_Serial12 ));
    CascadeMux I__1192 (
            .O(N__9731),
            .I(\c0.tx.N_294_cascade_ ));
    InMux I__1191 (
            .O(N__9728),
            .I(N__9725));
    LocalMux I__1190 (
            .O(N__9725),
            .I(\c0.tx.m5_0_0 ));
    InMux I__1189 (
            .O(N__9722),
            .I(N__9718));
    InMux I__1188 (
            .O(N__9721),
            .I(N__9715));
    LocalMux I__1187 (
            .O(N__9718),
            .I(\c0.tx.N_287 ));
    LocalMux I__1186 (
            .O(N__9715),
            .I(\c0.tx.N_287 ));
    CascadeMux I__1185 (
            .O(N__9710),
            .I(\c0.tx.N_288_cascade_ ));
    InMux I__1184 (
            .O(N__9707),
            .I(N__9704));
    LocalMux I__1183 (
            .O(N__9704),
            .I(blink_counterZ0Z_17));
    InMux I__1182 (
            .O(N__9701),
            .I(blink_counter_cry_16));
    InMux I__1181 (
            .O(N__9698),
            .I(N__9695));
    LocalMux I__1180 (
            .O(N__9695),
            .I(blink_counterZ0Z_18));
    InMux I__1179 (
            .O(N__9692),
            .I(blink_counter_cry_17));
    InMux I__1178 (
            .O(N__9689),
            .I(N__9686));
    LocalMux I__1177 (
            .O(N__9686),
            .I(blink_counterZ0Z_19));
    InMux I__1176 (
            .O(N__9683),
            .I(blink_counter_cry_18));
    InMux I__1175 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__1174 (
            .O(N__9677),
            .I(blink_counterZ0Z_20));
    InMux I__1173 (
            .O(N__9674),
            .I(blink_counter_cry_19));
    InMux I__1172 (
            .O(N__9671),
            .I(N__9668));
    LocalMux I__1171 (
            .O(N__9668),
            .I(N__9665));
    Span4Mux_h I__1170 (
            .O(N__9665),
            .I(N__9661));
    InMux I__1169 (
            .O(N__9664),
            .I(N__9658));
    Odrv4 I__1168 (
            .O(N__9661),
            .I(blink_counterZ0Z_21));
    LocalMux I__1167 (
            .O(N__9658),
            .I(blink_counterZ0Z_21));
    InMux I__1166 (
            .O(N__9653),
            .I(blink_counter_cry_20));
    InMux I__1165 (
            .O(N__9650),
            .I(N__9644));
    InMux I__1164 (
            .O(N__9649),
            .I(N__9644));
    LocalMux I__1163 (
            .O(N__9644),
            .I(N__9641));
    Span4Mux_v I__1162 (
            .O(N__9641),
            .I(N__9637));
    InMux I__1161 (
            .O(N__9640),
            .I(N__9634));
    Odrv4 I__1160 (
            .O(N__9637),
            .I(blink_counterZ0Z_22));
    LocalMux I__1159 (
            .O(N__9634),
            .I(blink_counterZ0Z_22));
    InMux I__1158 (
            .O(N__9629),
            .I(blink_counter_cry_21));
    CascadeMux I__1157 (
            .O(N__9626),
            .I(N__9623));
    InMux I__1156 (
            .O(N__9623),
            .I(N__9620));
    LocalMux I__1155 (
            .O(N__9620),
            .I(N__9617));
    Span4Mux_v I__1154 (
            .O(N__9617),
            .I(N__9613));
    InMux I__1153 (
            .O(N__9616),
            .I(N__9610));
    Odrv4 I__1152 (
            .O(N__9613),
            .I(blink_counterZ0Z_23));
    LocalMux I__1151 (
            .O(N__9610),
            .I(blink_counterZ0Z_23));
    InMux I__1150 (
            .O(N__9605),
            .I(blink_counter_cry_22));
    CascadeMux I__1149 (
            .O(N__9602),
            .I(N__9599));
    InMux I__1148 (
            .O(N__9599),
            .I(N__9593));
    InMux I__1147 (
            .O(N__9598),
            .I(N__9593));
    LocalMux I__1146 (
            .O(N__9593),
            .I(N__9590));
    Span4Mux_v I__1145 (
            .O(N__9590),
            .I(N__9586));
    InMux I__1144 (
            .O(N__9589),
            .I(N__9583));
    Odrv4 I__1143 (
            .O(N__9586),
            .I(blink_counterZ0Z_24));
    LocalMux I__1142 (
            .O(N__9583),
            .I(blink_counterZ0Z_24));
    InMux I__1141 (
            .O(N__9578),
            .I(bfn_6_23_0_));
    InMux I__1140 (
            .O(N__9575),
            .I(N__9572));
    LocalMux I__1139 (
            .O(N__9572),
            .I(blink_counterZ0Z_9));
    InMux I__1138 (
            .O(N__9569),
            .I(blink_counter_cry_8));
    InMux I__1137 (
            .O(N__9566),
            .I(N__9563));
    LocalMux I__1136 (
            .O(N__9563),
            .I(blink_counterZ0Z_10));
    InMux I__1135 (
            .O(N__9560),
            .I(blink_counter_cry_9));
    InMux I__1134 (
            .O(N__9557),
            .I(N__9554));
    LocalMux I__1133 (
            .O(N__9554),
            .I(blink_counterZ0Z_11));
    InMux I__1132 (
            .O(N__9551),
            .I(blink_counter_cry_10));
    InMux I__1131 (
            .O(N__9548),
            .I(N__9545));
    LocalMux I__1130 (
            .O(N__9545),
            .I(blink_counterZ0Z_12));
    InMux I__1129 (
            .O(N__9542),
            .I(blink_counter_cry_11));
    InMux I__1128 (
            .O(N__9539),
            .I(N__9536));
    LocalMux I__1127 (
            .O(N__9536),
            .I(blink_counterZ0Z_13));
    InMux I__1126 (
            .O(N__9533),
            .I(blink_counter_cry_12));
    InMux I__1125 (
            .O(N__9530),
            .I(N__9527));
    LocalMux I__1124 (
            .O(N__9527),
            .I(blink_counterZ0Z_14));
    InMux I__1123 (
            .O(N__9524),
            .I(blink_counter_cry_13));
    InMux I__1122 (
            .O(N__9521),
            .I(N__9518));
    LocalMux I__1121 (
            .O(N__9518),
            .I(blink_counterZ0Z_15));
    InMux I__1120 (
            .O(N__9515),
            .I(blink_counter_cry_14));
    InMux I__1119 (
            .O(N__9512),
            .I(N__9509));
    LocalMux I__1118 (
            .O(N__9509),
            .I(blink_counterZ0Z_16));
    InMux I__1117 (
            .O(N__9506),
            .I(bfn_6_22_0_));
    InMux I__1116 (
            .O(N__9503),
            .I(N__9500));
    LocalMux I__1115 (
            .O(N__9500),
            .I(blink_counterZ0Z_0));
    InMux I__1114 (
            .O(N__9497),
            .I(bfn_6_20_0_));
    InMux I__1113 (
            .O(N__9494),
            .I(N__9491));
    LocalMux I__1112 (
            .O(N__9491),
            .I(blink_counterZ0Z_1));
    InMux I__1111 (
            .O(N__9488),
            .I(blink_counter_cry_0));
    InMux I__1110 (
            .O(N__9485),
            .I(N__9482));
    LocalMux I__1109 (
            .O(N__9482),
            .I(blink_counterZ0Z_2));
    InMux I__1108 (
            .O(N__9479),
            .I(blink_counter_cry_1));
    InMux I__1107 (
            .O(N__9476),
            .I(N__9473));
    LocalMux I__1106 (
            .O(N__9473),
            .I(blink_counterZ0Z_3));
    InMux I__1105 (
            .O(N__9470),
            .I(blink_counter_cry_2));
    InMux I__1104 (
            .O(N__9467),
            .I(N__9464));
    LocalMux I__1103 (
            .O(N__9464),
            .I(blink_counterZ0Z_4));
    InMux I__1102 (
            .O(N__9461),
            .I(blink_counter_cry_3));
    InMux I__1101 (
            .O(N__9458),
            .I(N__9455));
    LocalMux I__1100 (
            .O(N__9455),
            .I(blink_counterZ0Z_5));
    InMux I__1099 (
            .O(N__9452),
            .I(blink_counter_cry_4));
    InMux I__1098 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1097 (
            .O(N__9446),
            .I(blink_counterZ0Z_6));
    InMux I__1096 (
            .O(N__9443),
            .I(blink_counter_cry_5));
    InMux I__1095 (
            .O(N__9440),
            .I(N__9437));
    LocalMux I__1094 (
            .O(N__9437),
            .I(blink_counterZ0Z_7));
    InMux I__1093 (
            .O(N__9434),
            .I(blink_counter_cry_6));
    InMux I__1092 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__1091 (
            .O(N__9428),
            .I(blink_counterZ0Z_8));
    InMux I__1090 (
            .O(N__9425),
            .I(bfn_6_21_0_));
    InMux I__1089 (
            .O(N__9422),
            .I(\c0.tx.un1_r_Clock_Count_cry_0 ));
    InMux I__1088 (
            .O(N__9419),
            .I(N__9416));
    LocalMux I__1087 (
            .O(N__9416),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_2 ));
    InMux I__1086 (
            .O(N__9413),
            .I(\c0.tx.un1_r_Clock_Count_cry_1 ));
    InMux I__1085 (
            .O(N__9410),
            .I(\c0.tx.un1_r_Clock_Count_cry_2 ));
    CascadeMux I__1084 (
            .O(N__9407),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_3_cascade_ ));
    InMux I__1083 (
            .O(N__9404),
            .I(N__9401));
    LocalMux I__1082 (
            .O(N__9401),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_0 ));
    InMux I__1081 (
            .O(N__9398),
            .I(N__9394));
    InMux I__1080 (
            .O(N__9397),
            .I(N__9391));
    LocalMux I__1079 (
            .O(N__9394),
            .I(\c0.tx.r_Clock_CountZ0Z_0 ));
    LocalMux I__1078 (
            .O(N__9391),
            .I(\c0.tx.r_Clock_CountZ0Z_0 ));
    CascadeMux I__1077 (
            .O(N__9386),
            .I(N__9382));
    InMux I__1076 (
            .O(N__9385),
            .I(N__9379));
    InMux I__1075 (
            .O(N__9382),
            .I(N__9376));
    LocalMux I__1074 (
            .O(N__9379),
            .I(\c0.tx.r_Clock_Count_0_sqmuxa ));
    LocalMux I__1073 (
            .O(N__9376),
            .I(\c0.tx.r_Clock_Count_0_sqmuxa ));
    InMux I__1072 (
            .O(N__9371),
            .I(N__9368));
    LocalMux I__1071 (
            .O(N__9368),
            .I(\c0.tx.r_Clock_Count_RNO_0Z0Z_1 ));
    CascadeMux I__1070 (
            .O(N__9365),
            .I(\c0.rx.g0_i_a4_0_3_cascade_ ));
    InMux I__1069 (
            .O(N__9362),
            .I(N__9356));
    InMux I__1068 (
            .O(N__9361),
            .I(N__9353));
    InMux I__1067 (
            .O(N__9360),
            .I(N__9348));
    InMux I__1066 (
            .O(N__9359),
            .I(N__9348));
    LocalMux I__1065 (
            .O(N__9356),
            .I(\c0.rx.r_Clock_Count14_3 ));
    LocalMux I__1064 (
            .O(N__9353),
            .I(\c0.rx.r_Clock_Count14_3 ));
    LocalMux I__1063 (
            .O(N__9348),
            .I(\c0.rx.r_Clock_Count14_3 ));
    InMux I__1062 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__1061 (
            .O(N__9338),
            .I(\c0.rx.N_13 ));
    InMux I__1060 (
            .O(N__9335),
            .I(N__9331));
    InMux I__1059 (
            .O(N__9334),
            .I(N__9328));
    LocalMux I__1058 (
            .O(N__9331),
            .I(N__9322));
    LocalMux I__1057 (
            .O(N__9328),
            .I(N__9322));
    CascadeMux I__1056 (
            .O(N__9327),
            .I(N__9316));
    Span4Mux_h I__1055 (
            .O(N__9322),
            .I(N__9309));
    InMux I__1054 (
            .O(N__9321),
            .I(N__9306));
    InMux I__1053 (
            .O(N__9320),
            .I(N__9297));
    InMux I__1052 (
            .O(N__9319),
            .I(N__9297));
    InMux I__1051 (
            .O(N__9316),
            .I(N__9297));
    InMux I__1050 (
            .O(N__9315),
            .I(N__9297));
    InMux I__1049 (
            .O(N__9314),
            .I(N__9292));
    InMux I__1048 (
            .O(N__9313),
            .I(N__9292));
    InMux I__1047 (
            .O(N__9312),
            .I(N__9289));
    Odrv4 I__1046 (
            .O(N__9309),
            .I(\c0.rx.r_Clock_Count26 ));
    LocalMux I__1045 (
            .O(N__9306),
            .I(\c0.rx.r_Clock_Count26 ));
    LocalMux I__1044 (
            .O(N__9297),
            .I(\c0.rx.r_Clock_Count26 ));
    LocalMux I__1043 (
            .O(N__9292),
            .I(\c0.rx.r_Clock_Count26 ));
    LocalMux I__1042 (
            .O(N__9289),
            .I(\c0.rx.r_Clock_Count26 ));
    CascadeMux I__1041 (
            .O(N__9278),
            .I(N__9272));
    CascadeMux I__1040 (
            .O(N__9277),
            .I(N__9269));
    CascadeMux I__1039 (
            .O(N__9276),
            .I(N__9266));
    CascadeMux I__1038 (
            .O(N__9275),
            .I(N__9259));
    InMux I__1037 (
            .O(N__9272),
            .I(N__9255));
    InMux I__1036 (
            .O(N__9269),
            .I(N__9252));
    InMux I__1035 (
            .O(N__9266),
            .I(N__9249));
    CascadeMux I__1034 (
            .O(N__9265),
            .I(N__9244));
    CascadeMux I__1033 (
            .O(N__9264),
            .I(N__9236));
    CascadeMux I__1032 (
            .O(N__9263),
            .I(N__9229));
    CascadeMux I__1031 (
            .O(N__9262),
            .I(N__9226));
    InMux I__1030 (
            .O(N__9259),
            .I(N__9220));
    InMux I__1029 (
            .O(N__9258),
            .I(N__9220));
    LocalMux I__1028 (
            .O(N__9255),
            .I(N__9217));
    LocalMux I__1027 (
            .O(N__9252),
            .I(N__9214));
    LocalMux I__1026 (
            .O(N__9249),
            .I(N__9211));
    InMux I__1025 (
            .O(N__9248),
            .I(N__9204));
    InMux I__1024 (
            .O(N__9247),
            .I(N__9204));
    InMux I__1023 (
            .O(N__9244),
            .I(N__9204));
    CascadeMux I__1022 (
            .O(N__9243),
            .I(N__9201));
    CascadeMux I__1021 (
            .O(N__9242),
            .I(N__9197));
    CascadeMux I__1020 (
            .O(N__9241),
            .I(N__9192));
    CascadeMux I__1019 (
            .O(N__9240),
            .I(N__9188));
    InMux I__1018 (
            .O(N__9239),
            .I(N__9185));
    InMux I__1017 (
            .O(N__9236),
            .I(N__9180));
    InMux I__1016 (
            .O(N__9235),
            .I(N__9180));
    InMux I__1015 (
            .O(N__9234),
            .I(N__9175));
    InMux I__1014 (
            .O(N__9233),
            .I(N__9175));
    InMux I__1013 (
            .O(N__9232),
            .I(N__9166));
    InMux I__1012 (
            .O(N__9229),
            .I(N__9166));
    InMux I__1011 (
            .O(N__9226),
            .I(N__9166));
    InMux I__1010 (
            .O(N__9225),
            .I(N__9166));
    LocalMux I__1009 (
            .O(N__9220),
            .I(N__9161));
    Span4Mux_h I__1008 (
            .O(N__9217),
            .I(N__9161));
    Span4Mux_h I__1007 (
            .O(N__9214),
            .I(N__9156));
    Span4Mux_h I__1006 (
            .O(N__9211),
            .I(N__9156));
    LocalMux I__1005 (
            .O(N__9204),
            .I(N__9153));
    InMux I__1004 (
            .O(N__9201),
            .I(N__9144));
    InMux I__1003 (
            .O(N__9200),
            .I(N__9144));
    InMux I__1002 (
            .O(N__9197),
            .I(N__9144));
    InMux I__1001 (
            .O(N__9196),
            .I(N__9144));
    InMux I__1000 (
            .O(N__9195),
            .I(N__9135));
    InMux I__999 (
            .O(N__9192),
            .I(N__9135));
    InMux I__998 (
            .O(N__9191),
            .I(N__9135));
    InMux I__997 (
            .O(N__9188),
            .I(N__9135));
    LocalMux I__996 (
            .O(N__9185),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    LocalMux I__995 (
            .O(N__9180),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    LocalMux I__994 (
            .O(N__9175),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    LocalMux I__993 (
            .O(N__9166),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    Odrv4 I__992 (
            .O(N__9161),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    Odrv4 I__991 (
            .O(N__9156),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    Odrv4 I__990 (
            .O(N__9153),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    LocalMux I__989 (
            .O(N__9144),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    LocalMux I__988 (
            .O(N__9135),
            .I(\c0.rx.r_SM_MainZ0Z_2 ));
    CascadeMux I__987 (
            .O(N__9116),
            .I(\c0.rx.r_Rx_DV_1_sqmuxa_cascade_ ));
    CascadeMux I__986 (
            .O(N__9113),
            .I(N__9110));
    InMux I__985 (
            .O(N__9110),
            .I(N__9104));
    InMux I__984 (
            .O(N__9109),
            .I(N__9101));
    InMux I__983 (
            .O(N__9108),
            .I(N__9098));
    CascadeMux I__982 (
            .O(N__9107),
            .I(N__9089));
    LocalMux I__981 (
            .O(N__9104),
            .I(N__9085));
    LocalMux I__980 (
            .O(N__9101),
            .I(N__9079));
    LocalMux I__979 (
            .O(N__9098),
            .I(N__9079));
    InMux I__978 (
            .O(N__9097),
            .I(N__9065));
    InMux I__977 (
            .O(N__9096),
            .I(N__9065));
    InMux I__976 (
            .O(N__9095),
            .I(N__9062));
    InMux I__975 (
            .O(N__9094),
            .I(N__9051));
    InMux I__974 (
            .O(N__9093),
            .I(N__9051));
    InMux I__973 (
            .O(N__9092),
            .I(N__9051));
    InMux I__972 (
            .O(N__9089),
            .I(N__9051));
    InMux I__971 (
            .O(N__9088),
            .I(N__9051));
    Span4Mux_h I__970 (
            .O(N__9085),
            .I(N__9048));
    InMux I__969 (
            .O(N__9084),
            .I(N__9045));
    Span4Mux_h I__968 (
            .O(N__9079),
            .I(N__9042));
    InMux I__967 (
            .O(N__9078),
            .I(N__9031));
    InMux I__966 (
            .O(N__9077),
            .I(N__9031));
    InMux I__965 (
            .O(N__9076),
            .I(N__9031));
    InMux I__964 (
            .O(N__9075),
            .I(N__9031));
    InMux I__963 (
            .O(N__9074),
            .I(N__9031));
    InMux I__962 (
            .O(N__9073),
            .I(N__9022));
    InMux I__961 (
            .O(N__9072),
            .I(N__9022));
    InMux I__960 (
            .O(N__9071),
            .I(N__9022));
    InMux I__959 (
            .O(N__9070),
            .I(N__9022));
    LocalMux I__958 (
            .O(N__9065),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    LocalMux I__957 (
            .O(N__9062),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    LocalMux I__956 (
            .O(N__9051),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    Odrv4 I__955 (
            .O(N__9048),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    LocalMux I__954 (
            .O(N__9045),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    Odrv4 I__953 (
            .O(N__9042),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    LocalMux I__952 (
            .O(N__9031),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    LocalMux I__951 (
            .O(N__9022),
            .I(\c0.rx.r_SM_MainZ0Z_1 ));
    InMux I__950 (
            .O(N__9005),
            .I(N__9000));
    InMux I__949 (
            .O(N__9004),
            .I(N__8997));
    InMux I__948 (
            .O(N__9003),
            .I(N__8982));
    LocalMux I__947 (
            .O(N__9000),
            .I(N__8977));
    LocalMux I__946 (
            .O(N__8997),
            .I(N__8977));
    InMux I__945 (
            .O(N__8996),
            .I(N__8974));
    InMux I__944 (
            .O(N__8995),
            .I(N__8969));
    InMux I__943 (
            .O(N__8994),
            .I(N__8969));
    InMux I__942 (
            .O(N__8993),
            .I(N__8966));
    InMux I__941 (
            .O(N__8992),
            .I(N__8957));
    InMux I__940 (
            .O(N__8991),
            .I(N__8957));
    InMux I__939 (
            .O(N__8990),
            .I(N__8957));
    InMux I__938 (
            .O(N__8989),
            .I(N__8957));
    InMux I__937 (
            .O(N__8988),
            .I(N__8948));
    InMux I__936 (
            .O(N__8987),
            .I(N__8948));
    InMux I__935 (
            .O(N__8986),
            .I(N__8948));
    InMux I__934 (
            .O(N__8985),
            .I(N__8948));
    LocalMux I__933 (
            .O(N__8982),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    Odrv4 I__932 (
            .O(N__8977),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__931 (
            .O(N__8974),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__930 (
            .O(N__8969),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__929 (
            .O(N__8966),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__928 (
            .O(N__8957),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    LocalMux I__927 (
            .O(N__8948),
            .I(\c0.rx.r_SM_MainZ0Z_0 ));
    InMux I__926 (
            .O(N__8933),
            .I(N__8925));
    InMux I__925 (
            .O(N__8932),
            .I(N__8925));
    InMux I__924 (
            .O(N__8931),
            .I(N__8922));
    InMux I__923 (
            .O(N__8930),
            .I(N__8919));
    LocalMux I__922 (
            .O(N__8925),
            .I(\c0.rx.r_Clock_Count14 ));
    LocalMux I__921 (
            .O(N__8922),
            .I(\c0.rx.r_Clock_Count14 ));
    LocalMux I__920 (
            .O(N__8919),
            .I(\c0.rx.r_Clock_Count14 ));
    InMux I__919 (
            .O(N__8912),
            .I(N__8909));
    LocalMux I__918 (
            .O(N__8909),
            .I(\c0.rx.N_9 ));
    InMux I__917 (
            .O(N__8906),
            .I(N__8902));
    InMux I__916 (
            .O(N__8905),
            .I(N__8896));
    LocalMux I__915 (
            .O(N__8902),
            .I(N__8890));
    InMux I__914 (
            .O(N__8901),
            .I(N__8883));
    InMux I__913 (
            .O(N__8900),
            .I(N__8883));
    InMux I__912 (
            .O(N__8899),
            .I(N__8883));
    LocalMux I__911 (
            .O(N__8896),
            .I(N__8880));
    InMux I__910 (
            .O(N__8895),
            .I(N__8873));
    InMux I__909 (
            .O(N__8894),
            .I(N__8870));
    InMux I__908 (
            .O(N__8893),
            .I(N__8867));
    Span4Mux_s3_h I__907 (
            .O(N__8890),
            .I(N__8860));
    LocalMux I__906 (
            .O(N__8883),
            .I(N__8860));
    Span4Mux_h I__905 (
            .O(N__8880),
            .I(N__8860));
    InMux I__904 (
            .O(N__8879),
            .I(N__8855));
    InMux I__903 (
            .O(N__8878),
            .I(N__8855));
    InMux I__902 (
            .O(N__8877),
            .I(N__8852));
    InMux I__901 (
            .O(N__8876),
            .I(N__8849));
    LocalMux I__900 (
            .O(N__8873),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    LocalMux I__899 (
            .O(N__8870),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    LocalMux I__898 (
            .O(N__8867),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    Odrv4 I__897 (
            .O(N__8860),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    LocalMux I__896 (
            .O(N__8855),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    LocalMux I__895 (
            .O(N__8852),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    LocalMux I__894 (
            .O(N__8849),
            .I(\c0.rx.r_Clock_CountZ0Z_0 ));
    CascadeMux I__893 (
            .O(N__8834),
            .I(N__8828));
    InMux I__892 (
            .O(N__8833),
            .I(N__8822));
    InMux I__891 (
            .O(N__8832),
            .I(N__8818));
    InMux I__890 (
            .O(N__8831),
            .I(N__8813));
    InMux I__889 (
            .O(N__8828),
            .I(N__8813));
    InMux I__888 (
            .O(N__8827),
            .I(N__8808));
    InMux I__887 (
            .O(N__8826),
            .I(N__8808));
    InMux I__886 (
            .O(N__8825),
            .I(N__8802));
    LocalMux I__885 (
            .O(N__8822),
            .I(N__8799));
    InMux I__884 (
            .O(N__8821),
            .I(N__8796));
    LocalMux I__883 (
            .O(N__8818),
            .I(N__8789));
    LocalMux I__882 (
            .O(N__8813),
            .I(N__8789));
    LocalMux I__881 (
            .O(N__8808),
            .I(N__8789));
    InMux I__880 (
            .O(N__8807),
            .I(N__8784));
    InMux I__879 (
            .O(N__8806),
            .I(N__8784));
    InMux I__878 (
            .O(N__8805),
            .I(N__8781));
    LocalMux I__877 (
            .O(N__8802),
            .I(\c0.rx.r_Clock_CountZ0Z_1 ));
    Odrv4 I__876 (
            .O(N__8799),
            .I(\c0.rx.r_Clock_CountZ0Z_1 ));
    LocalMux I__875 (
            .O(N__8796),
            .I(\c0.rx.r_Clock_CountZ0Z_1 ));
    Odrv4 I__874 (
            .O(N__8789),
            .I(\c0.rx.r_Clock_CountZ0Z_1 ));
    LocalMux I__873 (
            .O(N__8784),
            .I(\c0.rx.r_Clock_CountZ0Z_1 ));
    LocalMux I__872 (
            .O(N__8781),
            .I(\c0.rx.r_Clock_CountZ0Z_1 ));
    InMux I__871 (
            .O(N__8768),
            .I(N__8765));
    LocalMux I__870 (
            .O(N__8765),
            .I(\c0.rx.r_Clock_Count14_1 ));
    CascadeMux I__869 (
            .O(N__8762),
            .I(N__8759));
    InMux I__868 (
            .O(N__8759),
            .I(N__8756));
    LocalMux I__867 (
            .O(N__8756),
            .I(\c0.rx.N_12_0 ));
    CascadeMux I__866 (
            .O(N__8753),
            .I(\c0.rx.N_9_0_cascade_ ));
    InMux I__865 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__864 (
            .O(N__8747),
            .I(N__8744));
    Odrv4 I__863 (
            .O(N__8744),
            .I(\c0.rx.N_11_i ));
    InMux I__862 (
            .O(N__8741),
            .I(N__8737));
    InMux I__861 (
            .O(N__8740),
            .I(N__8733));
    LocalMux I__860 (
            .O(N__8737),
            .I(N__8730));
    InMux I__859 (
            .O(N__8736),
            .I(N__8727));
    LocalMux I__858 (
            .O(N__8733),
            .I(\c0.rx.r_Clock_CountZ0Z_6 ));
    Odrv4 I__857 (
            .O(N__8730),
            .I(\c0.rx.r_Clock_CountZ0Z_6 ));
    LocalMux I__856 (
            .O(N__8727),
            .I(\c0.rx.r_Clock_CountZ0Z_6 ));
    InMux I__855 (
            .O(N__8720),
            .I(N__8716));
    InMux I__854 (
            .O(N__8719),
            .I(N__8713));
    LocalMux I__853 (
            .O(N__8716),
            .I(N__8710));
    LocalMux I__852 (
            .O(N__8713),
            .I(N__8705));
    Span4Mux_h I__851 (
            .O(N__8710),
            .I(N__8702));
    InMux I__850 (
            .O(N__8709),
            .I(N__8699));
    InMux I__849 (
            .O(N__8708),
            .I(N__8696));
    Odrv4 I__848 (
            .O(N__8705),
            .I(\c0.rx.r_Clock_CountZ0Z_5 ));
    Odrv4 I__847 (
            .O(N__8702),
            .I(\c0.rx.r_Clock_CountZ0Z_5 ));
    LocalMux I__846 (
            .O(N__8699),
            .I(\c0.rx.r_Clock_CountZ0Z_5 ));
    LocalMux I__845 (
            .O(N__8696),
            .I(\c0.rx.r_Clock_CountZ0Z_5 ));
    CascadeMux I__844 (
            .O(N__8687),
            .I(N__8684));
    InMux I__843 (
            .O(N__8684),
            .I(N__8680));
    InMux I__842 (
            .O(N__8683),
            .I(N__8677));
    LocalMux I__841 (
            .O(N__8680),
            .I(N__8674));
    LocalMux I__840 (
            .O(N__8677),
            .I(\c0.rx.r_Clock_CountZ0Z_7 ));
    Odrv4 I__839 (
            .O(N__8674),
            .I(\c0.rx.r_Clock_CountZ0Z_7 ));
    CascadeMux I__838 (
            .O(N__8669),
            .I(N__8663));
    InMux I__837 (
            .O(N__8668),
            .I(N__8658));
    InMux I__836 (
            .O(N__8667),
            .I(N__8655));
    InMux I__835 (
            .O(N__8666),
            .I(N__8652));
    InMux I__834 (
            .O(N__8663),
            .I(N__8649));
    InMux I__833 (
            .O(N__8662),
            .I(N__8646));
    InMux I__832 (
            .O(N__8661),
            .I(N__8643));
    LocalMux I__831 (
            .O(N__8658),
            .I(\c0.rx.r_Clock_CountZ0Z_4 ));
    LocalMux I__830 (
            .O(N__8655),
            .I(\c0.rx.r_Clock_CountZ0Z_4 ));
    LocalMux I__829 (
            .O(N__8652),
            .I(\c0.rx.r_Clock_CountZ0Z_4 ));
    LocalMux I__828 (
            .O(N__8649),
            .I(\c0.rx.r_Clock_CountZ0Z_4 ));
    LocalMux I__827 (
            .O(N__8646),
            .I(\c0.rx.r_Clock_CountZ0Z_4 ));
    LocalMux I__826 (
            .O(N__8643),
            .I(\c0.rx.r_Clock_CountZ0Z_4 ));
    CascadeMux I__825 (
            .O(N__8630),
            .I(\c0.rx.r_Clock_Count14_3_cascade_ ));
    CascadeMux I__824 (
            .O(N__8627),
            .I(\c0.rx.r_Clock_Count26_cascade_ ));
    CascadeMux I__823 (
            .O(N__8624),
            .I(N__8617));
    InMux I__822 (
            .O(N__8623),
            .I(N__8608));
    InMux I__821 (
            .O(N__8622),
            .I(N__8605));
    InMux I__820 (
            .O(N__8621),
            .I(N__8602));
    InMux I__819 (
            .O(N__8620),
            .I(N__8599));
    InMux I__818 (
            .O(N__8617),
            .I(N__8596));
    InMux I__817 (
            .O(N__8616),
            .I(N__8593));
    InMux I__816 (
            .O(N__8615),
            .I(N__8586));
    InMux I__815 (
            .O(N__8614),
            .I(N__8586));
    InMux I__814 (
            .O(N__8613),
            .I(N__8586));
    InMux I__813 (
            .O(N__8612),
            .I(N__8583));
    InMux I__812 (
            .O(N__8611),
            .I(N__8580));
    LocalMux I__811 (
            .O(N__8608),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__810 (
            .O(N__8605),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__809 (
            .O(N__8602),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__808 (
            .O(N__8599),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__807 (
            .O(N__8596),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__806 (
            .O(N__8593),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__805 (
            .O(N__8586),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__804 (
            .O(N__8583),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    LocalMux I__803 (
            .O(N__8580),
            .I(\c0.rx.r_Clock_CountZ0Z_2 ));
    InMux I__802 (
            .O(N__8561),
            .I(N__8556));
    InMux I__801 (
            .O(N__8560),
            .I(N__8550));
    InMux I__800 (
            .O(N__8559),
            .I(N__8545));
    LocalMux I__799 (
            .O(N__8556),
            .I(N__8542));
    InMux I__798 (
            .O(N__8555),
            .I(N__8535));
    InMux I__797 (
            .O(N__8554),
            .I(N__8535));
    InMux I__796 (
            .O(N__8553),
            .I(N__8535));
    LocalMux I__795 (
            .O(N__8550),
            .I(N__8532));
    InMux I__794 (
            .O(N__8549),
            .I(N__8529));
    InMux I__793 (
            .O(N__8548),
            .I(N__8524));
    LocalMux I__792 (
            .O(N__8545),
            .I(N__8513));
    Span4Mux_v I__791 (
            .O(N__8542),
            .I(N__8513));
    LocalMux I__790 (
            .O(N__8535),
            .I(N__8513));
    Span4Mux_v I__789 (
            .O(N__8532),
            .I(N__8513));
    LocalMux I__788 (
            .O(N__8529),
            .I(N__8513));
    InMux I__787 (
            .O(N__8528),
            .I(N__8508));
    InMux I__786 (
            .O(N__8527),
            .I(N__8508));
    LocalMux I__785 (
            .O(N__8524),
            .I(\c0.rx.r_Clock_CountZ0Z_3 ));
    Odrv4 I__784 (
            .O(N__8513),
            .I(\c0.rx.r_Clock_CountZ0Z_3 ));
    LocalMux I__783 (
            .O(N__8508),
            .I(\c0.rx.r_Clock_CountZ0Z_3 ));
    InMux I__782 (
            .O(N__8501),
            .I(N__8495));
    InMux I__781 (
            .O(N__8500),
            .I(N__8495));
    LocalMux I__780 (
            .O(N__8495),
            .I(\c0.rx.r_Clock_Count_1_sqmuxa_0 ));
    CascadeMux I__779 (
            .O(N__8492),
            .I(\c0.rx.un1_r_Clock_Count_5_m_1_cascade_ ));
    InMux I__778 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__777 (
            .O(N__8486),
            .I(N_12));
    InMux I__776 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__775 (
            .O(N__8480),
            .I(N_8_0));
    IoInMux I__774 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__773 (
            .O(N__8474),
            .I(N__8471));
    Span4Mux_s0_v I__772 (
            .O(N__8471),
            .I(N__8468));
    Span4Mux_v I__771 (
            .O(N__8468),
            .I(N__8465));
    Odrv4 I__770 (
            .O(N__8465),
            .I(LED_c));
    CascadeMux I__769 (
            .O(N__8462),
            .I(\c0.rx.CO1_cascade_ ));
    CascadeMux I__768 (
            .O(N__8459),
            .I(\c0.rx.g0_i_o3_0_4_cascade_ ));
    InMux I__767 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__766 (
            .O(N__8453),
            .I(\c0.rx.N_10 ));
    InMux I__765 (
            .O(N__8450),
            .I(N__8447));
    LocalMux I__764 (
            .O(N__8447),
            .I(\c0.rx.g1_4 ));
    CascadeMux I__763 (
            .O(N__8444),
            .I(\c0.rx.g1_5_cascade_ ));
    InMux I__762 (
            .O(N__8441),
            .I(N__8438));
    LocalMux I__761 (
            .O(N__8438),
            .I(\c0.rx.g1 ));
    CascadeMux I__760 (
            .O(N__8435),
            .I(\c0.rx.g0_0_1_cascade_ ));
    CascadeMux I__759 (
            .O(N__8432),
            .I(\c0.rx.r_Clock_Count14_cascade_ ));
    InMux I__758 (
            .O(N__8429),
            .I(N__8426));
    LocalMux I__757 (
            .O(N__8426),
            .I(\c0.rx.m6_ns_1 ));
    CascadeMux I__756 (
            .O(N__8423),
            .I(\c0.rx.un1_r_Clock_Count_5_m_0_cascade_ ));
    InMux I__755 (
            .O(N__8420),
            .I(N__8415));
    InMux I__754 (
            .O(N__8419),
            .I(N__8410));
    InMux I__753 (
            .O(N__8418),
            .I(N__8410));
    LocalMux I__752 (
            .O(N__8415),
            .I(\c0.rx.un1_r_Clock_Count_2_sqmuxa_0 ));
    LocalMux I__751 (
            .O(N__8410),
            .I(\c0.rx.un1_r_Clock_Count_2_sqmuxa_0 ));
    CascadeMux I__750 (
            .O(N__8405),
            .I(\c0.rx.N_7_cascade_ ));
    SRMux I__749 (
            .O(N__8402),
            .I(N__8399));
    LocalMux I__748 (
            .O(N__8399),
            .I(N__8396));
    Span4Mux_h I__747 (
            .O(N__8396),
            .I(N__8392));
    InMux I__746 (
            .O(N__8395),
            .I(N__8389));
    Odrv4 I__745 (
            .O(N__8392),
            .I(\c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1 ));
    LocalMux I__744 (
            .O(N__8389),
            .I(\c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1 ));
    InMux I__743 (
            .O(N__8384),
            .I(N__8381));
    LocalMux I__742 (
            .O(N__8381),
            .I(\c0.rx.N_10_0 ));
    InMux I__741 (
            .O(N__8378),
            .I(N__8375));
    LocalMux I__740 (
            .O(N__8375),
            .I(\c0.rx.N_13_0 ));
    CascadeMux I__739 (
            .O(N__8372),
            .I(\c0.rx.N_12_1_cascade_ ));
    InMux I__738 (
            .O(N__8369),
            .I(N__8366));
    LocalMux I__737 (
            .O(N__8366),
            .I(\c0.rx.un1_r_Clock_Count_5_c2 ));
    CascadeMux I__736 (
            .O(N__8363),
            .I(\c0.rx.N_6_cascade_ ));
    InMux I__735 (
            .O(N__8360),
            .I(N__8354));
    InMux I__734 (
            .O(N__8359),
            .I(N__8354));
    LocalMux I__733 (
            .O(N__8354),
            .I(\c0.rx.r_Clock_Count_2_sqmuxa_0 ));
    CascadeMux I__732 (
            .O(N__8351),
            .I(\c0.rx.r_Clock_Count_2_sqmuxa_0_cascade_ ));
    CascadeMux I__731 (
            .O(N__8348),
            .I(\c0.rx.g0_i_o4_0_1_cascade_ ));
    CascadeMux I__730 (
            .O(N__8345),
            .I(\c0.rx.g0_i_o2_2_3_cascade_ ));
    InMux I__729 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__728 (
            .O(N__8339),
            .I(\c0.rx.g0_i_a4_1_1 ));
    IoInMux I__727 (
            .O(N__8336),
            .I(N__8333));
    LocalMux I__726 (
            .O(N__8333),
            .I(N__8330));
    Span4Mux_s0_v I__725 (
            .O(N__8330),
            .I(N__8326));
    CascadeMux I__724 (
            .O(N__8329),
            .I(N__8323));
    Span4Mux_v I__723 (
            .O(N__8326),
            .I(N__8320));
    InMux I__722 (
            .O(N__8323),
            .I(N__8317));
    Odrv4 I__721 (
            .O(N__8320),
            .I(PIN_1_c));
    LocalMux I__720 (
            .O(N__8317),
            .I(PIN_1_c));
    CEMux I__719 (
            .O(N__8312),
            .I(N__8309));
    LocalMux I__718 (
            .O(N__8309),
            .I(N__8306));
    Odrv4 I__717 (
            .O(N__8306),
            .I(\c0.rx.un1_r_Rx_DV7_0 ));
    InMux I__716 (
            .O(N__8303),
            .I(N__8300));
    LocalMux I__715 (
            .O(N__8300),
            .I(\c0.rx.g0_i_o2_5 ));
    InMux I__714 (
            .O(N__8297),
            .I(N__8294));
    LocalMux I__713 (
            .O(N__8294),
            .I(\c0.rx.g0_i_o2_4 ));
    CascadeMux I__712 (
            .O(N__8291),
            .I(N__8288));
    InMux I__711 (
            .O(N__8288),
            .I(N__8285));
    LocalMux I__710 (
            .O(N__8285),
            .I(\c0.rx.g0_i_o2_6 ));
    InMux I__709 (
            .O(N__8282),
            .I(N__8279));
    LocalMux I__708 (
            .O(N__8279),
            .I(\c0.rx.g0_i_a4_1_3 ));
    InMux I__707 (
            .O(N__8276),
            .I(N__8273));
    LocalMux I__706 (
            .O(N__8273),
            .I(N__8270));
    Odrv12 I__705 (
            .O(N__8270),
            .I(PIN_2_c));
    InMux I__704 (
            .O(N__8267),
            .I(N__8264));
    LocalMux I__703 (
            .O(N__8264),
            .I(\c0.rx.r_Rx_Data_RZ0 ));
    IoInMux I__702 (
            .O(N__8261),
            .I(N__8258));
    LocalMux I__701 (
            .O(N__8258),
            .I(N__8255));
    IoSpan4Mux I__700 (
            .O(N__8255),
            .I(N__8252));
    Odrv4 I__699 (
            .O(N__8252),
            .I(\c0.rx.rx_data_ready ));
    CascadeMux I__698 (
            .O(N__8249),
            .I(\c0.rx.un1_r_Clock_Count_5_c2_cascade_ ));
    IoInMux I__697 (
            .O(N__8246),
            .I(N__8243));
    LocalMux I__696 (
            .O(N__8243),
            .I(N__8240));
    IoSpan4Mux I__695 (
            .O(N__8240),
            .I(N__8237));
    IoSpan4Mux I__694 (
            .O(N__8237),
            .I(N__8234));
    IoSpan4Mux I__693 (
            .O(N__8234),
            .I(N__8231));
    Odrv4 I__692 (
            .O(N__8231),
            .I(CLK_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_6_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_25_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\c0.i12 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\c0.data_cry_7 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_6_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_20_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(blink_counter_cry_7),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(blink_counter_cry_15),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(blink_counter_cry_23),
            .carryinitout(bfn_6_23_0_));
    ICE_GB CLK_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__8246),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    ICE_GB \c0.rx.r_Rx_DV_e_RNIHVG2  (
            .USERSIGNALTOGLOBALBUFFER(N__8261),
            .GLOBALBUFFEROUTPUT(\c0.rx_data_ready_g ));
    ICE_GB \c0.byte_transmit_counter_RNIA0ET3_0_2  (
            .USERSIGNALTOGLOBALBUFFER(N__16949),
            .GLOBALBUFFEROUTPUT(\c0.data_out_0__1_sqmuxa_g ));
    ICE_GB \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_0  (
            .USERSIGNALTOGLOBALBUFFER(N__12278),
            .GLOBALBUFFEROUTPUT(\c0.data_in_frame_0__0_sqmuxa_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_LC_2_23_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_LC_2_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_LC_2_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8267),
            .lcout(\c0.rx.r_Rx_DataZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21826),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_R_LC_2_24_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_LC_2_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_LC_2_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_R_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8276),
            .lcout(\c0.rx.r_Rx_Data_RZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_e_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_e_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_e_LC_3_19_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.rx.r_Rx_DV_e_LC_3_19_2  (
            .in0(N__9005),
            .in1(N__9109),
            .in2(N__9277),
            .in3(N__9335),
            .lcout(\c0.rx.rx_data_ready ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21824),
            .ce(N__8312),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_1_7_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_1_7_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_1_7_LC_3_21_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_1_7_LC_3_21_0  (
            .in0(N__8906),
            .in1(N__8720),
            .in2(N__9278),
            .in3(N__8667),
            .lcout(\c0.rx.g0_i_o2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_2_7_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_2_7_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_2_7_LC_3_21_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_2_7_LC_3_21_5  (
            .in0(N__8621),
            .in1(N__8741),
            .in2(N__9113),
            .in3(N__8832),
            .lcout(\c0.rx.g0_i_o2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_7_LC_3_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_7_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_7_LC_3_21_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_7_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__8993),
            .in2(_gnd_net_),
            .in3(N__8548),
            .lcout(\c0.rx.g0_i_o2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNIPDG17_1_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNIPDG17_1_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNIPDG17_1_LC_3_22_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.rx.r_Clock_Count_RNIPDG17_1_LC_3_22_0  (
            .in0(N__8831),
            .in1(N__8901),
            .in2(_gnd_net_),
            .in3(N__8420),
            .lcout(\c0.rx.un1_r_Clock_Count_5_c2 ),
            .ltout(\c0.rx.un1_r_Clock_Count_5_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_3_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_3_LC_3_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_3_LC_3_22_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \c0.rx.r_Clock_Count_3_LC_3_22_1  (
            .in0(N__8622),
            .in1(N__8395),
            .in2(N__8249),
            .in3(N__8555),
            .lcout(\c0.rx.r_Clock_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21827),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_3_4_LC_3_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_3_4_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_3_4_LC_3_22_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_3_4_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__9248),
            .in2(_gnd_net_),
            .in3(N__8900),
            .lcout(),
            .ltout(\c0.rx.g0_i_o4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_4_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_4_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_4_LC_3_22_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_4_LC_3_22_3  (
            .in0(N__8827),
            .in1(N__8615),
            .in2(N__8348),
            .in3(N__8554),
            .lcout(\c0.rx.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_4_4_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_4_4_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_4_4_LC_3_22_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_4_4_LC_3_22_5  (
            .in0(N__8826),
            .in1(N__8342),
            .in2(N__9265),
            .in3(N__8613),
            .lcout(\c0.rx.g0_i_a4_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_3_5_LC_3_22_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_3_5_LC_3_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_3_5_LC_3_22_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_3_5_LC_3_22_6  (
            .in0(N__8614),
            .in1(N__8899),
            .in2(N__8834),
            .in3(N__9247),
            .lcout(),
            .ltout(\c0.rx.g0_i_o2_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_1_5_LC_3_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_1_5_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_1_5_LC_3_22_7 .LUT_INIT=16'b0101100101010101;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_1_5_LC_3_22_7  (
            .in0(N__8719),
            .in1(N__8553),
            .in2(N__8345),
            .in3(N__8666),
            .lcout(\c0.rx.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_2_2_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_2_2_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_2_2_LC_3_23_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_2_2_LC_3_23_1  (
            .in0(N__8879),
            .in1(N__8616),
            .in2(N__21193),
            .in3(N__8821),
            .lcout(\c0.rx.g1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_5_4_LC_3_23_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_5_4_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_5_4_LC_3_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_5_4_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__8878),
            .in2(_gnd_net_),
            .in3(N__8662),
            .lcout(\c0.rx.g0_i_a4_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_LC_3_25_3 .SEQ_MODE=4'b1001;
    defparam \c0.tx.o_Tx_Serial_LC_3_25_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \c0.tx.o_Tx_Serial_LC_3_25_3  (
            .in0(N__10261),
            .in1(N__9956),
            .in2(N__8329),
            .in3(N__10403),
            .lcout(PIN_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21842),
            .ce(),
            .sr(N__9779));
    defparam \c0.rx.r_Rx_DV_e_RNO_LC_4_19_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_e_RNO_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_DV_e_RNO_LC_4_19_5 .LUT_INIT=16'b0001000100011001;
    LogicCell40 \c0.rx.r_Rx_DV_e_RNO_LC_4_19_5  (
            .in0(N__9108),
            .in1(N__9004),
            .in2(N__9276),
            .in3(N__9334),
            .lcout(\c0.rx.un1_r_Rx_DV7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_7_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_7_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_7_LC_4_21_2 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \c0.rx.r_Clock_Count_7_LC_4_21_2  (
            .in0(N__8303),
            .in1(N__8297),
            .in2(N__8291),
            .in3(N__8683),
            .lcout(\c0.rx.r_Clock_CountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21828),
            .ce(),
            .sr(N__8402));
    defparam \c0.rx.r_Clock_Count_RNO_2_4_LC_4_22_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_2_4_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_2_4_LC_4_22_0 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_2_4_LC_4_22_0  (
            .in0(N__8282),
            .in1(N__8559),
            .in2(N__9107),
            .in3(N__9361),
            .lcout(\c0.rx.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_8_1_0__m6_ns_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_8_1_0__m6_ns_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_8_1_0__m6_ns_LC_4_22_1 .LUT_INIT=16'b1000110001110111;
    LogicCell40 \c0.rx.r_SM_Main_8_1_0__m6_ns_LC_4_22_1  (
            .in0(N__9320),
            .in1(N__9094),
            .in2(N__10850),
            .in3(N__8429),
            .lcout(),
            .ltout(\c0.rx.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0_LC_4_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0_LC_4_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_0_LC_4_22_2 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \c0.rx.r_SM_Main_0_LC_4_22_2  (
            .in0(N__9232),
            .in1(_gnd_net_),
            .in2(N__8405),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21831),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNICMJF6_0_1_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNICMJF6_0_1_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNICMJF6_0_1_LC_4_22_3 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \c0.rx.r_SM_Main_RNICMJF6_0_1_LC_4_22_3  (
            .in0(N__8359),
            .in1(N__9225),
            .in2(N__9327),
            .in3(N__9088),
            .lcout(\c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_1_4_LC_4_22_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_1_4_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_1_4_LC_4_22_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_1_4_LC_4_22_4  (
            .in0(N__9093),
            .in1(N__8996),
            .in2(N__9263),
            .in3(N__9319),
            .lcout(),
            .ltout(\c0.rx.N_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_4_LC_4_22_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_4_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_4_LC_4_22_5 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \c0.rx.r_Clock_Count_4_LC_4_22_5  (
            .in0(N__8384),
            .in1(N__8378),
            .in2(N__8372),
            .in3(N__8668),
            .lcout(\c0.rx.r_Clock_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21831),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_2_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_2_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_2_LC_4_22_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_2_LC_4_22_6  (
            .in0(N__9092),
            .in1(N__9315),
            .in2(N__9262),
            .in3(N__8360),
            .lcout(),
            .ltout(\c0.rx.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_2_LC_4_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_2_LC_4_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_2_LC_4_22_7 .LUT_INIT=16'b1111111101100000;
    LogicCell40 \c0.rx.r_Clock_Count_2_LC_4_22_7  (
            .in0(N__8623),
            .in1(N__8369),
            .in2(N__8363),
            .in3(N__8441),
            .lcout(\c0.rx.r_Clock_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21831),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNIHR7E3_1_0_LC_4_23_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNIHR7E3_1_0_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNIHR7E3_1_0_LC_4_23_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.rx.r_SM_Main_RNIHR7E3_1_0_LC_4_23_0  (
            .in0(N__9070),
            .in1(N__8985),
            .in2(N__9240),
            .in3(N__8930),
            .lcout(\c0.rx.r_Clock_Count_2_sqmuxa_0 ),
            .ltout(\c0.rx.r_Clock_Count_2_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNICMJF6_1_LC_4_23_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNICMJF6_1_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNICMJF6_1_LC_4_23_1 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \c0.rx.r_SM_Main_RNICMJF6_1_LC_4_23_1  (
            .in0(N__9084),
            .in1(N__9191),
            .in2(N__8351),
            .in3(N__9312),
            .lcout(\c0.rx.un1_r_Clock_Count_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_3_2_LC_4_23_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_3_2_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_3_2_LC_4_23_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_3_2_LC_4_23_2  (
            .in0(N__9072),
            .in1(N__8986),
            .in2(N__9241),
            .in3(N__8528),
            .lcout(),
            .ltout(\c0.rx.g1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_1_2_LC_4_23_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_1_2_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_1_2_LC_4_23_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_1_2_LC_4_23_3  (
            .in0(N__8450),
            .in1(_gnd_net_),
            .in2(N__8444),
            .in3(N__9360),
            .lcout(\c0.rx.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNIGQSH_3_LC_4_23_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNIGQSH_3_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNIGQSH_3_LC_4_23_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNIGQSH_3_LC_4_23_4  (
            .in0(_gnd_net_),
            .in1(N__8527),
            .in2(_gnd_net_),
            .in3(N__8805),
            .lcout(),
            .ltout(\c0.rx.g0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNICMJ72_2_LC_4_23_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_2_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_2_LC_4_23_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNICMJ72_2_LC_4_23_5  (
            .in0(N__8611),
            .in1(N__8877),
            .in2(N__8435),
            .in3(N__9359),
            .lcout(\c0.rx.r_Clock_Count14 ),
            .ltout(\c0.rx.r_Clock_Count14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_8_1_0__m6_ns_1_LC_4_23_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_8_1_0__m6_ns_1_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_8_1_0__m6_ns_1_LC_4_23_6 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \c0.rx.r_SM_Main_8_1_0__m6_ns_1_LC_4_23_6  (
            .in0(N__9071),
            .in1(N__21194),
            .in2(N__8432),
            .in3(N__8987),
            .lcout(\c0.rx.m6_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_RNIIGH91_LC_4_23_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_RNIIGH91_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Data_RNIIGH91_LC_4_23_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \c0.rx.r_Rx_Data_RNIIGH91_LC_4_23_7  (
            .in0(N__8988),
            .in1(N__9195),
            .in2(N__21213),
            .in3(N__9073),
            .lcout(\c0.rx.r_Clock_Count_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_0_LC_4_24_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_0_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_0_LC_4_24_0 .LUT_INIT=16'b1000100000110011;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_0_LC_4_24_0  (
            .in0(N__9258),
            .in1(N__8418),
            .in2(_gnd_net_),
            .in3(N__8894),
            .lcout(),
            .ltout(\c0.rx.un1_r_Clock_Count_5_m_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_0_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_0_LC_4_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_0_LC_4_24_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \c0.rx.r_Clock_Count_0_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__8500),
            .in2(N__8423),
            .in3(N__8932),
            .lcout(\c0.rx.r_Clock_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21843),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_1_LC_4_24_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_1_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_1_LC_4_24_4 .LUT_INIT=16'b1101000100100010;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_1_LC_4_24_4  (
            .in0(N__8895),
            .in1(N__8419),
            .in2(N__9275),
            .in3(N__8825),
            .lcout(),
            .ltout(\c0.rx.un1_r_Clock_Count_5_m_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_1_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_1_LC_4_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_1_LC_4_24_5 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \c0.rx.r_Clock_Count_1_LC_4_24_5  (
            .in0(_gnd_net_),
            .in1(N__8501),
            .in2(N__8492),
            .in3(N__8933),
            .lcout(\c0.rx.r_Clock_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21843),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_obuf_RNO_0_LC_4_25_1.C_ON=1'b0;
    defparam LED_obuf_RNO_0_LC_4_25_1.SEQ_MODE=4'b0000;
    defparam LED_obuf_RNO_0_LC_4_25_1.LUT_INIT=16'b0010001000100010;
    LogicCell40 LED_obuf_RNO_0_LC_4_25_1 (
            .in0(N__9649),
            .in1(N__9598),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_obuf_RNO_1_LC_4_25_6.C_ON=1'b0;
    defparam LED_obuf_RNO_1_LC_4_25_6.SEQ_MODE=4'b0000;
    defparam LED_obuf_RNO_1_LC_4_25_6.LUT_INIT=16'b1110110100000000;
    LogicCell40 LED_obuf_RNO_1_LC_4_25_6 (
            .in0(N__9811),
            .in1(N__9650),
            .in2(N__9602),
            .in3(N__9671),
            .lcout(N_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_obuf_RNO_LC_4_26_0.C_ON=1'b0;
    defparam LED_obuf_RNO_LC_4_26_0.SEQ_MODE=4'b0000;
    defparam LED_obuf_RNO_LC_4_26_0.LUT_INIT=16'b0100010100010101;
    LogicCell40 LED_obuf_RNO_LC_4_26_0 (
            .in0(N__8489),
            .in1(N__8483),
            .in2(N__9626),
            .in3(N__9812),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_RNO_0_2_LC_5_21_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_RNO_0_2_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Bit_Index_RNO_0_2_LC_5_21_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.r_Bit_Index_RNO_0_2_LC_5_21_2  (
            .in0(N__21410),
            .in1(N__21304),
            .in2(_gnd_net_),
            .in3(N__21096),
            .lcout(),
            .ltout(\c0.rx.CO1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_2_LC_5_21_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_2_LC_5_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_2_LC_5_21_3 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \c0.rx.r_Bit_Index_2_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(N__9924),
            .in2(N__8462),
            .in3(N__21452),
            .lcout(\c0.rx.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21832),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_6_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_6_LC_5_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_6_LC_5_21_5 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \c0.rx.r_Clock_Count_6_LC_5_21_5  (
            .in0(N__9234),
            .in1(N__8456),
            .in2(N__8762),
            .in3(N__8740),
            .lcout(\c0.rx.r_Clock_CountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21832),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_2_6_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_2_6_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_2_6_LC_5_21_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_2_6_LC_5_21_6  (
            .in0(N__8905),
            .in1(N__8709),
            .in2(N__8669),
            .in3(N__9233),
            .lcout(),
            .ltout(\c0.rx.g0_i_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_6_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_6_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_6_LC_5_21_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_6_LC_5_21_7  (
            .in0(N__8620),
            .in1(N__8561),
            .in2(N__8459),
            .in3(N__8833),
            .lcout(\c0.rx.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNI55K61_0_LC_5_22_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNI55K61_0_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNI55K61_0_LC_5_22_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \c0.rx.r_SM_Main_RNI55K61_0_LC_5_22_0  (
            .in0(N__8991),
            .in1(_gnd_net_),
            .in2(N__9242),
            .in3(N__9075),
            .lcout(\c0.rx.r_Rx_DV6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_1_6_LC_5_22_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_1_6_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_1_6_LC_5_22_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_1_6_LC_5_22_1  (
            .in0(N__9076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8990),
            .lcout(\c0.rx.N_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2_LC_5_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2_LC_5_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_2_LC_5_22_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.rx.r_SM_Main_2_LC_5_22_2  (
            .in0(N__9314),
            .in1(N__9078),
            .in2(N__9243),
            .in3(N__9003),
            .lcout(\c0.rx.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21836),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_0_5_LC_5_22_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_0_5_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_0_5_LC_5_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_0_5_LC_5_22_3  (
            .in0(N__9077),
            .in1(N__8992),
            .in2(_gnd_net_),
            .in3(N__9313),
            .lcout(),
            .ltout(\c0.rx.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_5_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_5_LC_5_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count_5_LC_5_22_4 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \c0.rx.r_Clock_Count_5_LC_5_22_4  (
            .in0(N__9200),
            .in1(N__9341),
            .in2(N__8753),
            .in3(N__8750),
            .lcout(\c0.rx.r_Clock_CountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21836),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_5_22_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_5_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_5_22_5  (
            .in0(N__8736),
            .in1(N__8708),
            .in2(N__8687),
            .in3(N__8661),
            .lcout(\c0.rx.r_Clock_Count14_3 ),
            .ltout(\c0.rx.r_Clock_Count14_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNICMJ72_3_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_3_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNICMJ72_3_LC_5_22_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \c0.rx.r_Clock_Count_RNICMJ72_3_LC_5_22_6  (
            .in0(N__8612),
            .in1(N__8768),
            .in2(N__8630),
            .in3(N__8549),
            .lcout(\c0.rx.r_Clock_Count26 ),
            .ltout(\c0.rx.r_Clock_Count26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNIHR7E3_0_0_LC_5_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNIHR7E3_0_0_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNIHR7E3_0_0_LC_5_22_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.rx.r_SM_Main_RNIHR7E3_0_0_LC_5_22_7  (
            .in0(N__9074),
            .in1(N__9196),
            .in2(N__8627),
            .in3(N__8989),
            .lcout(\c0.rx.r_Rx_Byte_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_4_5_LC_5_23_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_4_5_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_4_5_LC_5_23_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_4_5_LC_5_23_0  (
            .in0(N__8807),
            .in1(N__8893),
            .in2(N__8624),
            .in3(N__8560),
            .lcout(),
            .ltout(\c0.rx.g0_i_a4_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNO_2_5_LC_5_23_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNO_2_5_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNO_2_5_LC_5_23_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNO_2_5_LC_5_23_1  (
            .in0(N__9235),
            .in1(N__9095),
            .in2(N__9365),
            .in3(N__9362),
            .lcout(\c0.rx.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_RNIHR7E3_0_LC_5_23_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_RNIHR7E3_0_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_RNIHR7E3_0_LC_5_23_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.rx.r_SM_Main_RNIHR7E3_0_LC_5_23_3  (
            .in0(N__9096),
            .in1(N__8994),
            .in2(N__9264),
            .in3(N__9321),
            .lcout(),
            .ltout(\c0.rx.r_Rx_DV_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_1_LC_5_23_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_1_LC_5_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_1_LC_5_23_4 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \c0.rx.r_SM_Main_1_LC_5_23_4  (
            .in0(N__9239),
            .in1(N__9097),
            .in2(N__9116),
            .in3(N__8912),
            .lcout(\c0.rx.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21844),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_8_1_0__m8_LC_5_23_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_8_1_0__m8_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_8_1_0__m8_LC_5_23_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.rx.r_SM_Main_8_1_0__m8_LC_5_23_6  (
            .in0(N__8995),
            .in1(N__21214),
            .in2(_gnd_net_),
            .in3(N__8931),
            .lcout(\c0.rx.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count_RNIDNSH_1_LC_5_23_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count_RNIDNSH_1_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Clock_Count_RNIDNSH_1_LC_5_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.r_Clock_Count_RNIDNSH_1_LC_5_23_7  (
            .in0(_gnd_net_),
            .in1(N__8876),
            .in2(_gnd_net_),
            .in3(N__8806),
            .lcout(\c0.rx.r_Clock_Count14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_0_LC_5_24_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_0_LC_5_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_0_LC_5_24_0 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \c0.tx.r_SM_Main_0_LC_5_24_0  (
            .in0(N__9728),
            .in1(N__10045),
            .in2(N__10409),
            .in3(N__9785),
            .lcout(\c0.tx.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21851),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_2_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_2_LC_5_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_2_LC_5_24_2 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.tx.r_Clock_Count_2_LC_5_24_2  (
            .in0(N__10260),
            .in1(N__9419),
            .in2(N__9766),
            .in3(N__10318),
            .lcout(\c0.tx.r_Clock_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21851),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_24_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_24_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_24_6  (
            .in0(N__13360),
            .in1(N__9397),
            .in2(_gnd_net_),
            .in3(N__9884),
            .lcout(\c0.tx.r_Clock_Count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_0_LC_5_25_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count_RNO_0_0_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_0_LC_5_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_0_LC_5_25_0  (
            .in0(_gnd_net_),
            .in1(N__9398),
            .in2(N__9386),
            .in3(N__9385),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(\c0.tx.un1_r_Clock_Count_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_1_LC_5_25_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count_RNO_0_1_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_1_LC_5_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_1_LC_5_25_1  (
            .in0(_gnd_net_),
            .in1(N__9872),
            .in2(_gnd_net_),
            .in3(N__9422),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\c0.tx.un1_r_Clock_Count_cry_0 ),
            .carryout(\c0.tx.un1_r_Clock_Count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_2_LC_5_25_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count_RNO_0_2_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_2_LC_5_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_2_LC_5_25_2  (
            .in0(_gnd_net_),
            .in1(N__9854),
            .in2(_gnd_net_),
            .in3(N__9413),
            .lcout(\c0.tx.r_Clock_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\c0.tx.un1_r_Clock_Count_cry_1 ),
            .carryout(\c0.tx.un1_r_Clock_Count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_RNO_0_3_LC_5_25_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_RNO_0_3_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count_RNO_0_3_LC_5_25_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.tx.r_Clock_Count_RNO_0_3_LC_5_25_3  (
            .in0(_gnd_net_),
            .in1(N__9836),
            .in2(_gnd_net_),
            .in3(N__9410),
            .lcout(),
            .ltout(\c0.tx.r_Clock_Count_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_3_LC_5_25_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_3_LC_5_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_3_LC_5_25_4 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \c0.tx.r_Clock_Count_3_LC_5_25_4  (
            .in0(N__10246),
            .in1(N__9773),
            .in2(N__9407),
            .in3(N__10303),
            .lcout(\c0.tx.r_Clock_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21858),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_0_LC_5_25_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_0_LC_5_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_0_LC_5_25_5 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.tx.r_Clock_Count_0_LC_5_25_5  (
            .in0(N__10301),
            .in1(N__10244),
            .in2(N__9777),
            .in3(N__9404),
            .lcout(\c0.tx.r_Clock_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21858),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNIFAME1_0_LC_5_25_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNIFAME1_0_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNIFAME1_0_LC_5_25_6 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.tx.r_SM_Main_RNIFAME1_0_LC_5_25_6  (
            .in0(N__10402),
            .in1(N__10439),
            .in2(N__10259),
            .in3(N__10300),
            .lcout(\c0.tx.r_Clock_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count_1_LC_5_25_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count_1_LC_5_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count_1_LC_5_25_7 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.tx.r_Clock_Count_1_LC_5_25_7  (
            .in0(N__10302),
            .in1(N__10245),
            .in2(N__9778),
            .in3(N__9371),
            .lcout(\c0.tx.r_Clock_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21858),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNID5VK2_21_LC_5_26_7 .C_ON=1'b0;
    defparam \c0.d_2_RNID5VK2_21_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNID5VK2_21_LC_5_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNID5VK2_21_LC_5_26_7  (
            .in0(N__11587),
            .in1(N__11833),
            .in2(N__11064),
            .in3(N__11649),
            .lcout(\c0.nextCRC16_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_5_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_5_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_5_LC_6_19_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_5_LC_6_19_0  (
            .in0(N__21395),
            .in1(N__21461),
            .in2(_gnd_net_),
            .in3(N__21295),
            .lcout(\c0.rx.r_Rx_Bytece_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_0_LC_6_20_0.C_ON=1'b1;
    defparam blink_counter_0_LC_6_20_0.SEQ_MODE=4'b1000;
    defparam blink_counter_0_LC_6_20_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_0_LC_6_20_0 (
            .in0(_gnd_net_),
            .in1(N__9503),
            .in2(_gnd_net_),
            .in3(N__9497),
            .lcout(blink_counterZ0Z_0),
            .ltout(),
            .carryin(bfn_6_20_0_),
            .carryout(blink_counter_cry_0),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_1_LC_6_20_1.C_ON=1'b1;
    defparam blink_counter_1_LC_6_20_1.SEQ_MODE=4'b1000;
    defparam blink_counter_1_LC_6_20_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_1_LC_6_20_1 (
            .in0(_gnd_net_),
            .in1(N__9494),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(blink_counterZ0Z_1),
            .ltout(),
            .carryin(blink_counter_cry_0),
            .carryout(blink_counter_cry_1),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2_LC_6_20_2.C_ON=1'b1;
    defparam blink_counter_2_LC_6_20_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2_LC_6_20_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_2_LC_6_20_2 (
            .in0(_gnd_net_),
            .in1(N__9485),
            .in2(_gnd_net_),
            .in3(N__9479),
            .lcout(blink_counterZ0Z_2),
            .ltout(),
            .carryin(blink_counter_cry_1),
            .carryout(blink_counter_cry_2),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_3_LC_6_20_3.C_ON=1'b1;
    defparam blink_counter_3_LC_6_20_3.SEQ_MODE=4'b1000;
    defparam blink_counter_3_LC_6_20_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_3_LC_6_20_3 (
            .in0(_gnd_net_),
            .in1(N__9476),
            .in2(_gnd_net_),
            .in3(N__9470),
            .lcout(blink_counterZ0Z_3),
            .ltout(),
            .carryin(blink_counter_cry_2),
            .carryout(blink_counter_cry_3),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_4_LC_6_20_4.C_ON=1'b1;
    defparam blink_counter_4_LC_6_20_4.SEQ_MODE=4'b1000;
    defparam blink_counter_4_LC_6_20_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_4_LC_6_20_4 (
            .in0(_gnd_net_),
            .in1(N__9467),
            .in2(_gnd_net_),
            .in3(N__9461),
            .lcout(blink_counterZ0Z_4),
            .ltout(),
            .carryin(blink_counter_cry_3),
            .carryout(blink_counter_cry_4),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_5_LC_6_20_5.C_ON=1'b1;
    defparam blink_counter_5_LC_6_20_5.SEQ_MODE=4'b1000;
    defparam blink_counter_5_LC_6_20_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_5_LC_6_20_5 (
            .in0(_gnd_net_),
            .in1(N__9458),
            .in2(_gnd_net_),
            .in3(N__9452),
            .lcout(blink_counterZ0Z_5),
            .ltout(),
            .carryin(blink_counter_cry_4),
            .carryout(blink_counter_cry_5),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_6_LC_6_20_6.C_ON=1'b1;
    defparam blink_counter_6_LC_6_20_6.SEQ_MODE=4'b1000;
    defparam blink_counter_6_LC_6_20_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_6_LC_6_20_6 (
            .in0(_gnd_net_),
            .in1(N__9449),
            .in2(_gnd_net_),
            .in3(N__9443),
            .lcout(blink_counterZ0Z_6),
            .ltout(),
            .carryin(blink_counter_cry_5),
            .carryout(blink_counter_cry_6),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_7_LC_6_20_7.C_ON=1'b1;
    defparam blink_counter_7_LC_6_20_7.SEQ_MODE=4'b1000;
    defparam blink_counter_7_LC_6_20_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_7_LC_6_20_7 (
            .in0(_gnd_net_),
            .in1(N__9440),
            .in2(_gnd_net_),
            .in3(N__9434),
            .lcout(blink_counterZ0Z_7),
            .ltout(),
            .carryin(blink_counter_cry_6),
            .carryout(blink_counter_cry_7),
            .clk(N__21833),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_8_LC_6_21_0.C_ON=1'b1;
    defparam blink_counter_8_LC_6_21_0.SEQ_MODE=4'b1000;
    defparam blink_counter_8_LC_6_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_8_LC_6_21_0 (
            .in0(_gnd_net_),
            .in1(N__9431),
            .in2(_gnd_net_),
            .in3(N__9425),
            .lcout(blink_counterZ0Z_8),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(blink_counter_cry_8),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_9_LC_6_21_1.C_ON=1'b1;
    defparam blink_counter_9_LC_6_21_1.SEQ_MODE=4'b1000;
    defparam blink_counter_9_LC_6_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_9_LC_6_21_1 (
            .in0(_gnd_net_),
            .in1(N__9575),
            .in2(_gnd_net_),
            .in3(N__9569),
            .lcout(blink_counterZ0Z_9),
            .ltout(),
            .carryin(blink_counter_cry_8),
            .carryout(blink_counter_cry_9),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_10_LC_6_21_2.C_ON=1'b1;
    defparam blink_counter_10_LC_6_21_2.SEQ_MODE=4'b1000;
    defparam blink_counter_10_LC_6_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_10_LC_6_21_2 (
            .in0(_gnd_net_),
            .in1(N__9566),
            .in2(_gnd_net_),
            .in3(N__9560),
            .lcout(blink_counterZ0Z_10),
            .ltout(),
            .carryin(blink_counter_cry_9),
            .carryout(blink_counter_cry_10),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_11_LC_6_21_3.C_ON=1'b1;
    defparam blink_counter_11_LC_6_21_3.SEQ_MODE=4'b1000;
    defparam blink_counter_11_LC_6_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_11_LC_6_21_3 (
            .in0(_gnd_net_),
            .in1(N__9557),
            .in2(_gnd_net_),
            .in3(N__9551),
            .lcout(blink_counterZ0Z_11),
            .ltout(),
            .carryin(blink_counter_cry_10),
            .carryout(blink_counter_cry_11),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_12_LC_6_21_4.C_ON=1'b1;
    defparam blink_counter_12_LC_6_21_4.SEQ_MODE=4'b1000;
    defparam blink_counter_12_LC_6_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_12_LC_6_21_4 (
            .in0(_gnd_net_),
            .in1(N__9548),
            .in2(_gnd_net_),
            .in3(N__9542),
            .lcout(blink_counterZ0Z_12),
            .ltout(),
            .carryin(blink_counter_cry_11),
            .carryout(blink_counter_cry_12),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_13_LC_6_21_5.C_ON=1'b1;
    defparam blink_counter_13_LC_6_21_5.SEQ_MODE=4'b1000;
    defparam blink_counter_13_LC_6_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_13_LC_6_21_5 (
            .in0(_gnd_net_),
            .in1(N__9539),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(blink_counterZ0Z_13),
            .ltout(),
            .carryin(blink_counter_cry_12),
            .carryout(blink_counter_cry_13),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_14_LC_6_21_6.C_ON=1'b1;
    defparam blink_counter_14_LC_6_21_6.SEQ_MODE=4'b1000;
    defparam blink_counter_14_LC_6_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_14_LC_6_21_6 (
            .in0(_gnd_net_),
            .in1(N__9530),
            .in2(_gnd_net_),
            .in3(N__9524),
            .lcout(blink_counterZ0Z_14),
            .ltout(),
            .carryin(blink_counter_cry_13),
            .carryout(blink_counter_cry_14),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_15_LC_6_21_7.C_ON=1'b1;
    defparam blink_counter_15_LC_6_21_7.SEQ_MODE=4'b1000;
    defparam blink_counter_15_LC_6_21_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_15_LC_6_21_7 (
            .in0(_gnd_net_),
            .in1(N__9521),
            .in2(_gnd_net_),
            .in3(N__9515),
            .lcout(blink_counterZ0Z_15),
            .ltout(),
            .carryin(blink_counter_cry_14),
            .carryout(blink_counter_cry_15),
            .clk(N__21837),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_16_LC_6_22_0.C_ON=1'b1;
    defparam blink_counter_16_LC_6_22_0.SEQ_MODE=4'b1000;
    defparam blink_counter_16_LC_6_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_16_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(N__9512),
            .in2(_gnd_net_),
            .in3(N__9506),
            .lcout(blink_counterZ0Z_16),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(blink_counter_cry_16),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_17_LC_6_22_1.C_ON=1'b1;
    defparam blink_counter_17_LC_6_22_1.SEQ_MODE=4'b1000;
    defparam blink_counter_17_LC_6_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_17_LC_6_22_1 (
            .in0(_gnd_net_),
            .in1(N__9707),
            .in2(_gnd_net_),
            .in3(N__9701),
            .lcout(blink_counterZ0Z_17),
            .ltout(),
            .carryin(blink_counter_cry_16),
            .carryout(blink_counter_cry_17),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_18_LC_6_22_2.C_ON=1'b1;
    defparam blink_counter_18_LC_6_22_2.SEQ_MODE=4'b1000;
    defparam blink_counter_18_LC_6_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_18_LC_6_22_2 (
            .in0(_gnd_net_),
            .in1(N__9698),
            .in2(_gnd_net_),
            .in3(N__9692),
            .lcout(blink_counterZ0Z_18),
            .ltout(),
            .carryin(blink_counter_cry_17),
            .carryout(blink_counter_cry_18),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_19_LC_6_22_3.C_ON=1'b1;
    defparam blink_counter_19_LC_6_22_3.SEQ_MODE=4'b1000;
    defparam blink_counter_19_LC_6_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_19_LC_6_22_3 (
            .in0(_gnd_net_),
            .in1(N__9689),
            .in2(_gnd_net_),
            .in3(N__9683),
            .lcout(blink_counterZ0Z_19),
            .ltout(),
            .carryin(blink_counter_cry_18),
            .carryout(blink_counter_cry_19),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_20_LC_6_22_4.C_ON=1'b1;
    defparam blink_counter_20_LC_6_22_4.SEQ_MODE=4'b1000;
    defparam blink_counter_20_LC_6_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_20_LC_6_22_4 (
            .in0(_gnd_net_),
            .in1(N__9680),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(blink_counterZ0Z_20),
            .ltout(),
            .carryin(blink_counter_cry_19),
            .carryout(blink_counter_cry_20),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_21_LC_6_22_5.C_ON=1'b1;
    defparam blink_counter_21_LC_6_22_5.SEQ_MODE=4'b1000;
    defparam blink_counter_21_LC_6_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_21_LC_6_22_5 (
            .in0(_gnd_net_),
            .in1(N__9664),
            .in2(_gnd_net_),
            .in3(N__9653),
            .lcout(blink_counterZ0Z_21),
            .ltout(),
            .carryin(blink_counter_cry_20),
            .carryout(blink_counter_cry_21),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_22_LC_6_22_6.C_ON=1'b1;
    defparam blink_counter_22_LC_6_22_6.SEQ_MODE=4'b1000;
    defparam blink_counter_22_LC_6_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_22_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(N__9640),
            .in2(_gnd_net_),
            .in3(N__9629),
            .lcout(blink_counterZ0Z_22),
            .ltout(),
            .carryin(blink_counter_cry_21),
            .carryout(blink_counter_cry_22),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_23_LC_6_22_7.C_ON=1'b1;
    defparam blink_counter_23_LC_6_22_7.SEQ_MODE=4'b1000;
    defparam blink_counter_23_LC_6_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_23_LC_6_22_7 (
            .in0(_gnd_net_),
            .in1(N__9616),
            .in2(_gnd_net_),
            .in3(N__9605),
            .lcout(blink_counterZ0Z_23),
            .ltout(),
            .carryin(blink_counter_cry_22),
            .carryout(blink_counter_cry_23),
            .clk(N__21845),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_24_LC_6_23_0.C_ON=1'b1;
    defparam blink_counter_24_LC_6_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_24_LC_6_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 blink_counter_24_LC_6_23_0 (
            .in0(_gnd_net_),
            .in1(N__9589),
            .in2(_gnd_net_),
            .in3(N__9578),
            .lcout(blink_counterZ0Z_24),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(blink_counter_cry_24),
            .clk(N__21852),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_25_LC_6_23_1.C_ON=1'b0;
    defparam blink_counter_25_LC_6_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_25_LC_6_23_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 blink_counter_25_LC_6_23_1 (
            .in0(_gnd_net_),
            .in1(N__9799),
            .in2(_gnd_net_),
            .in3(N__9815),
            .lcout(blink_counterZ0Z_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21852),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0_LC_6_23_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0_LC_6_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_0_LC_6_23_5 .LUT_INIT=16'b1110000010100100;
    LogicCell40 \c0.tx.r_Bit_Index_0_LC_6_23_5  (
            .in0(N__9722),
            .in1(N__10369),
            .in2(N__9986),
            .in3(N__10328),
            .lcout(\c0.tx.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21852),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNIBPOV_0_LC_6_23_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNIBPOV_0_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNIBPOV_0_LC_6_23_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx.r_SM_Main_RNIBPOV_0_LC_6_23_7  (
            .in0(N__10240),
            .in1(N__10368),
            .in2(_gnd_net_),
            .in3(N__10453),
            .lcout(\c0.tx.o_Tx_Serial12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNIIR5L_0_LC_6_24_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNIIR5L_0_LC_6_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNIIR5L_0_LC_6_24_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.r_SM_Main_RNIIR5L_0_LC_6_24_0  (
            .in0(_gnd_net_),
            .in1(N__10253),
            .in2(_gnd_net_),
            .in3(N__10440),
            .lcout(\c0.tx.N_287 ),
            .ltout(\c0.tx.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_o2_LC_6_24_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_o2_LC_6_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_o2_LC_6_24_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.tx.r_SM_Main_7_1_0__m5_0_o2_LC_6_24_1  (
            .in0(N__9980),
            .in1(N__10021),
            .in2(N__9788),
            .in3(N__10304),
            .lcout(\c0.tx.N_294 ),
            .ltout(\c0.tx.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_2_LC_6_24_2 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_2_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_2_LC_6_24_2 .LUT_INIT=16'b0011000000000011;
    LogicCell40 \c0.tx.r_Bit_Index_2_LC_6_24_2  (
            .in0(_gnd_net_),
            .in1(N__9752),
            .in2(N__9731),
            .in3(N__10046),
            .lcout(\c0.tx.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21859),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_0_LC_6_24_4 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_0_LC_6_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_0_LC_6_24_4 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \c0.tx.r_SM_Main_7_1_0__m5_0_0_LC_6_24_4  (
            .in0(N__10305),
            .in1(N__10254),
            .in2(N__10940),
            .in3(N__10441),
            .lcout(\c0.tx.m5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_RNO_0_1_LC_6_24_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_RNO_0_1_LC_6_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_RNO_0_1_LC_6_24_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.tx.r_Bit_Index_RNO_0_1_LC_6_24_5  (
            .in0(N__9981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10306),
            .lcout(),
            .ltout(\c0.tx.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_1_LC_6_24_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_1_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_1_LC_6_24_6 .LUT_INIT=16'b1010100110001000;
    LogicCell40 \c0.tx.r_Bit_Index_1_LC_6_24_6  (
            .in0(N__10022),
            .in1(N__9721),
            .in2(N__9710),
            .in3(N__10407),
            .lcout(\c0.tx.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21859),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_5_LC_6_24_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_5_LC_6_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_5_LC_6_24_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx_data_RNO_1_5_LC_6_24_7  (
            .in0(N__19361),
            .in1(N__14558),
            .in2(N__10094),
            .in3(N__19238),
            .lcout(\c0.tx_data_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_0_c_LC_6_25_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_LC_6_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_0_c_LC_6_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_0_c_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(N__9883),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_25_0_),
            .carryout(\c0.tx.r_Clock_Count12_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_6_25_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_6_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_6_25_1  (
            .in0(_gnd_net_),
            .in1(N__9860),
            .in2(N__13386),
            .in3(N__9871),
            .lcout(\c0.tx.r_Clock_Count_i_1 ),
            .ltout(),
            .carryin(\c0.tx.r_Clock_Count12_cry_0 ),
            .carryout(\c0.tx.r_Clock_Count12_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_6_25_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_6_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_6_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__9842),
            .in2(N__13394),
            .in3(N__9853),
            .lcout(\c0.tx.r_Clock_Count_i_2 ),
            .ltout(),
            .carryin(\c0.tx.r_Clock_Count12_cry_1 ),
            .carryout(\c0.tx.r_Clock_Count12_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_6_25_3 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_6_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_6_25_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_6_25_3  (
            .in0(N__9835),
            .in1(N__9824),
            .in2(N__13387),
            .in3(_gnd_net_),
            .lcout(\c0.tx.r_Clock_Count_i_3 ),
            .ltout(),
            .carryin(\c0.tx.r_Clock_Count12_cry_2 ),
            .carryout(\c0.tx.r_Clock_Count12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_6_25_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_6_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_6_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_6_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9818),
            .lcout(\c0.tx.r_Clock_Count12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__3_LC_6_25_5 .C_ON=1'b0;
    defparam \c0.data_out_0__3_LC_6_25_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__3_LC_6_25_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_0__3_LC_6_25_5  (
            .in0(N__13361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21863),
            .ce(),
            .sr(N__17347));
    defparam \c0.data_out_0__7_LC_6_25_6 .C_ON=1'b0;
    defparam \c0.data_out_0__7_LC_6_25_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__7_LC_6_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__7_LC_6_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13362),
            .lcout(\c0.d_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21863),
            .ce(),
            .sr(N__17347));
    defparam \c0.data_out_3__3_LC_6_25_7 .C_ON=1'b0;
    defparam \c0.data_out_3__3_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__3_LC_6_25_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__3_LC_6_25_7  (
            .in0(N__13363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21863),
            .ce(),
            .sr(N__17347));
    defparam \c0.data_out_0__2_LC_6_26_0 .C_ON=1'b0;
    defparam \c0.data_out_0__2_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__2_LC_6_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__2_LC_6_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13388),
            .lcout(\c0.d_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21872),
            .ce(),
            .sr(N__17346));
    defparam \c0.data_out_1__7_LC_6_26_2 .C_ON=1'b0;
    defparam \c0.data_out_1__7_LC_6_26_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__7_LC_6_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__7_LC_6_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13390),
            .lcout(\c0.d_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21872),
            .ce(),
            .sr(N__17346));
    defparam \c0.data_out_1__3_LC_6_26_3 .C_ON=1'b0;
    defparam \c0.data_out_1__3_LC_6_26_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__3_LC_6_26_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__3_LC_6_26_3  (
            .in0(N__13389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21872),
            .ce(),
            .sr(N__17346));
    defparam \c0.data_out_2__2_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.data_out_2__2_LC_6_26_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__2_LC_6_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__2_LC_6_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13391),
            .lcout(\c0.d_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21872),
            .ce(),
            .sr(N__17346));
    defparam \c0.data_out_2__5_LC_6_26_5 .C_ON=1'b0;
    defparam \c0.data_out_2__5_LC_6_26_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__5_LC_6_26_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_2__5_LC_6_26_5  (
            .in0(N__13392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21872),
            .ce(),
            .sr(N__17346));
    defparam \c0.data_out_2__7_LC_6_26_6 .C_ON=1'b0;
    defparam \c0.data_out_2__7_LC_6_26_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__7_LC_6_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__7_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13393),
            .lcout(\c0.d_2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21872),
            .ce(),
            .sr(N__17346));
    defparam \c0.d_2_RNIIQK01_7_LC_6_27_0 .C_ON=1'b0;
    defparam \c0.d_2_RNIIQK01_7_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIIQK01_7_LC_6_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIIQK01_7_LC_6_27_0  (
            .in0(N__16541),
            .in1(N__16494),
            .in2(_gnd_net_),
            .in3(N__10510),
            .lcout(\c0.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_1_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_1_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_1_LC_7_20_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_1_LC_7_20_4  (
            .in0(N__21481),
            .in1(N__21396),
            .in2(_gnd_net_),
            .in3(N__21293),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_1_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_1_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_1_LC_7_20_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.rx.r_Rx_Byte_1_LC_7_20_5  (
            .in0(N__11332),
            .in1(N__21228),
            .in2(N__9893),
            .in3(N__21136),
            .lcout(\c0.rx_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21838),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_5_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_5_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_5_LC_7_20_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_5_LC_7_20_6  (
            .in0(N__21137),
            .in1(N__10783),
            .in2(N__21241),
            .in3(N__9890),
            .lcout(\c0.rx_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21838),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_0_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_0_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_0_LC_7_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \c0.rx.r_Bit_Index_0_LC_7_21_0  (
            .in0(N__9937),
            .in1(N__21294),
            .in2(_gnd_net_),
            .in3(N__21145),
            .lcout(\c0.rx.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_RNIRD3K_2_LC_7_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_RNIRD3K_2_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Bit_Index_RNIRD3K_2_LC_7_22_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.r_Bit_Index_RNIRD3K_2_LC_7_22_2  (
            .in0(N__21471),
            .in1(N__21363),
            .in2(_gnd_net_),
            .in3(N__21277),
            .lcout(\c0.rx.un1_r_Rx_Byte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_1_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_1_LC_7_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_1_LC_7_22_3 .LUT_INIT=16'b0000101000000110;
    LogicCell40 \c0.tx.r_SM_Main_1_LC_7_22_3  (
            .in0(N__10397),
            .in1(N__10471),
            .in2(N__10262),
            .in3(N__10320),
            .lcout(\c0.tx.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21853),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_1_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_1_LC_7_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_1_LC_7_22_5 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \c0.rx.r_Bit_Index_1_LC_7_22_5  (
            .in0(N__21278),
            .in1(N__9938),
            .in2(N__21390),
            .in3(N__21132),
            .lcout(\c0.rx.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21853),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_RNIFAME1_0_0_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_RNIFAME1_0_0_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_RNIFAME1_0_0_LC_7_23_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.tx.r_SM_Main_RNIFAME1_0_0_LC_7_23_1  (
            .in0(N__10378),
            .in1(N__10470),
            .in2(N__10255),
            .in3(N__10319),
            .lcout(),
            .ltout(\c0.tx.r_Tx_Active_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_LC_7_23_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_LC_7_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_LC_7_23_2 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \c0.tx.r_Tx_Active_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__10921),
            .in2(N__9911),
            .in3(N__14184),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21860),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_1_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_1_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_1_LC_7_23_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \c0.tx_data_RNO_0_1_LC_7_23_3  (
            .in0(N__19398),
            .in1(N__19205),
            .in2(N__10865),
            .in3(N__14959),
            .lcout(\c0.tx_data_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_1_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_1_LC_7_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_1_LC_7_24_0 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \c0.tx.r_Tx_Data_1_LC_7_24_0  (
            .in0(N__16876),
            .in1(N__9908),
            .in2(N__11039),
            .in3(N__10544),
            .lcout(\c0.tx.r_Tx_DataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21864),
            .ce(N__10942),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_3_LC_7_24_1 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_3_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_3_LC_7_24_1 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_3_LC_7_24_1  (
            .in0(N__9902),
            .in1(N__10043),
            .in2(N__10061),
            .in3(N__10017),
            .lcout(),
            .ltout(\c0.tx.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_1_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_1_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_1_LC_7_24_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_1_LC_7_24_2  (
            .in0(N__10018),
            .in1(N__10955),
            .in2(N__9896),
            .in3(N__10076),
            .lcout(\c0.tx.N_354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_3_LC_7_24_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_3_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_3_LC_7_24_3 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \c0.tx_data_RNO_2_3_LC_7_24_3  (
            .in0(N__10052),
            .in1(N__17567),
            .in2(N__16882),
            .in3(N__10826),
            .lcout(),
            .ltout(\c0.tx_data_1_0_i_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_3_LC_7_24_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_3_LC_7_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_3_LC_7_24_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx.r_Tx_Data_3_LC_7_24_4  (
            .in0(N__16877),
            .in1(N__14705),
            .in2(N__10079),
            .in3(N__10535),
            .lcout(\c0.tx.r_Tx_DataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21864),
            .ce(N__10942),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_5_LC_7_24_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_5_LC_7_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_5_LC_7_24_5 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \c0.tx.r_Tx_Data_5_LC_7_24_5  (
            .in0(N__16875),
            .in1(N__11090),
            .in2(N__10070),
            .in3(N__9944),
            .lcout(\c0.tx.r_Tx_DataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21864),
            .ce(N__10942),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_3_LC_7_25_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_3_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_3_LC_7_25_1 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \c0.tx_data_RNO_4_3_LC_7_25_1  (
            .in0(N__19410),
            .in1(N__19209),
            .in2(N__11903),
            .in3(N__15332),
            .lcout(\c0.tx_data_RNO_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_4_LC_7_25_2 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_4_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_4_LC_7_25_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_4_LC_7_25_2  (
            .in0(N__10112),
            .in1(N__10044),
            .in2(N__10103),
            .in3(N__10019),
            .lcout(),
            .ltout(\c0.tx.r_Tx_Data_pmux_3_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_2_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_2_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_2_LC_7_25_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_2_LC_7_25_3  (
            .in0(N__10020),
            .in1(N__10985),
            .in2(N__9995),
            .in3(N__10973),
            .lcout(),
            .ltout(\c0.tx.N_357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_RNO_0_LC_7_25_4 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_RNO_0_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_RNO_0_LC_7_25_4 .LUT_INIT=16'b0000000001000111;
    LogicCell40 \c0.tx.o_Tx_Serial_RNO_0_LC_7_25_4  (
            .in0(N__9992),
            .in1(N__9985),
            .in2(N__9959),
            .in3(N__10472),
            .lcout(\c0.tx.N_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_5_LC_7_25_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_5_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_5_LC_7_25_6 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx_data_RNO_3_5_LC_7_25_6  (
            .in0(N__15170),
            .in1(N__11257),
            .in2(N__19232),
            .in3(N__19397),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_5_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_5_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_5_LC_7_25_7 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_5_LC_7_25_7  (
            .in0(N__16868),
            .in1(N__17554),
            .in2(N__9947),
            .in3(N__12746),
            .lcout(\c0.tx_data_1_0_i_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_0_LC_7_26_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_0_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_0_LC_7_26_1 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_1_0_LC_7_26_1  (
            .in0(N__12839),
            .in1(N__17566),
            .in2(N__13436),
            .in3(N__16913),
            .lcout(),
            .ltout(\c0.tx_data_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_0_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_0_LC_7_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_0_LC_7_26_2 .LUT_INIT=16'b1111011110110011;
    LogicCell40 \c0.tx.r_Tx_Data_0_LC_7_26_2  (
            .in0(N__16883),
            .in1(N__11570),
            .in2(N__10115),
            .in3(N__11777),
            .lcout(\c0.tx.r_Tx_DataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21879),
            .ce(N__10943),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_4_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_4_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_4_LC_7_26_3 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \c0.tx.r_Tx_Data_4_LC_7_26_3  (
            .in0(N__16881),
            .in1(N__10145),
            .in2(N__10880),
            .in3(N__11186),
            .lcout(\c0.tx.r_Tx_DataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21879),
            .ce(N__10943),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__5_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.data_out_7__5_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__5_LC_7_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_7__5_LC_7_27_1  (
            .in0(N__10484),
            .in1(N__12038),
            .in2(_gnd_net_),
            .in3(N__12971),
            .lcout(\c0.data_out_7_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21887),
            .ce(N__17298),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__3_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.data_out_4__3_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__3_LC_7_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__3_LC_7_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10652),
            .lcout(\c0.d_2_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21887),
            .ce(N__17298),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__4_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.data_out_4__4_LC_7_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__4_LC_7_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__4_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10631),
            .lcout(\c0.d_2_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21897),
            .ce(N__17297),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__3_LC_9_16_2 .C_ON=1'b0;
    defparam \c0.data_in_0__3_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__3_LC_9_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__3_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13927),
            .lcout(\c0.data_in_0_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21825),
            .ce(N__22151),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_2_c_RNO_LC_9_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_2_c_RNO_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_2_c_RNO_LC_9_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_2_c_RNO_LC_9_17_0  (
            .in0(N__13887),
            .in1(N__14082),
            .in2(N__12361),
            .in3(N__13659),
            .lcout(\c0.i12_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__4_LC_9_17_1 .C_ON=1'b0;
    defparam \c0.data_in_1__4_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__4_LC_9_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_1__4_LC_9_17_1  (
            .in0(N__16197),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_1_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21834),
            .ce(N__22150),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__7_LC_9_17_3 .C_ON=1'b0;
    defparam \c0.data_in_1__7_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__7_LC_9_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__7_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15946),
            .lcout(\c0.data_in_1_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21834),
            .ce(N__22150),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__4_LC_9_17_6 .C_ON=1'b0;
    defparam \c0.data_in_2__4_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__4_LC_9_17_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_2__4_LC_9_17_6  (
            .in0(N__11443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_2_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21834),
            .ce(N__22150),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_5_c_RNO_LC_9_17_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_5_c_RNO_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_5_c_RNO_LC_9_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_5_c_RNO_LC_9_17_7  (
            .in0(N__18121),
            .in1(N__11419),
            .in2(N__16201),
            .in3(N__13755),
            .lcout(\c0.i12_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__0_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0__0_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__0_LC_9_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__0_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18301),
            .lcout(\c0.data_in_0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21839),
            .ce(N__22152),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__1_LC_9_18_1 .C_ON=1'b0;
    defparam \c0.data_in_2__1_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__1_LC_9_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__1_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13847),
            .lcout(\c0.data_in_2_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21839),
            .ce(N__22152),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__0_LC_9_18_2 .C_ON=1'b0;
    defparam \c0.data_in_2__0_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__0_LC_9_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__0_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18674),
            .lcout(\c0.data_in_2_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21839),
            .ce(N__22152),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__5_LC_9_18_3 .C_ON=1'b0;
    defparam \c0.data_in_1__5_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__5_LC_9_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__5_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13867),
            .lcout(\c0.data_in_1_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21839),
            .ce(N__22152),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__0_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.data_in_1__0_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__0_LC_9_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__0_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13660),
            .lcout(\c0.data_in_1_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21839),
            .ce(N__22152),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__5_LC_9_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0__5_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__5_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__5_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13891),
            .lcout(\c0.data_in_0_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21839),
            .ce(N__22152),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__7_LC_9_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0__7_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__7_LC_9_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__7_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12360),
            .lcout(\c0.data_in_0_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21847),
            .ce(N__22155),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__2_LC_9_19_2 .C_ON=1'b0;
    defparam \c0.data_in_1__2_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__2_LC_9_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__2_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16227),
            .lcout(\c0.data_in_1_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21847),
            .ce(N__22155),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__3_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.data_in_1__3_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__3_LC_9_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__3_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15424),
            .lcout(\c0.data_in_1_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21847),
            .ce(N__22155),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__3_LC_9_19_5 .C_ON=1'b0;
    defparam \c0.data_in_7__3_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__3_LC_9_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_7__3_LC_9_19_5  (
            .in0(N__10130),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_7_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21847),
            .ce(N__22155),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__1_LC_9_19_6 .C_ON=1'b0;
    defparam \c0.data_in_1__1_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__1_LC_9_19_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_in_1__1_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__13756),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_1_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21847),
            .ce(N__22155),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__2_LC_9_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0__2_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__2_LC_9_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__2_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16645),
            .lcout(\c0.data_in_0_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21847),
            .ce(N__22155),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_3_LC_9_20_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_3_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_3_LC_9_20_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_3_LC_9_20_5  (
            .in0(N__21494),
            .in1(N__21411),
            .in2(_gnd_net_),
            .in3(N__21315),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_3_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_3_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_3_LC_9_20_6 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.rx.r_Rx_Byte_3_LC_9_20_6  (
            .in0(N__10129),
            .in1(N__21227),
            .in2(N__10133),
            .in3(N__21146),
            .lcout(\c0.rx_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21854),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_2_LC_9_21_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_2_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_2_LC_9_21_2 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \c0.tx2_data_RNO_3_2_LC_9_21_2  (
            .in0(N__16628),
            .in1(N__18925),
            .in2(N__19563),
            .in3(N__12500),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_2_LC_9_21_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_2_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_2_LC_9_21_3 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \c0.tx2_data_RNO_2_2_LC_9_21_3  (
            .in0(N__10772),
            .in1(N__20354),
            .in2(N__10118),
            .in3(N__20939),
            .lcout(\c0.tx2_data_1_0_i_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__4_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.data_out_3__4_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__4_LC_9_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__4_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13330),
            .lcout(\c0.d_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21865),
            .ce(),
            .sr(N__17348));
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_a2_0_LC_9_23_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_a2_0_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_7_1_0__m5_0_a2_0_LC_9_23_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.tx.r_SM_Main_7_1_0__m5_0_a2_0_LC_9_23_2  (
            .in0(N__10398),
            .in1(N__14207),
            .in2(N__10239),
            .in3(N__10468),
            .lcout(\c0.tx.r_Tx_Data_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_5_6_LC_9_23_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_5_6_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_5_6_LC_9_23_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.tx_data_RNO_5_6_LC_9_23_4  (
            .in0(N__11703),
            .in1(N__19158),
            .in2(N__11995),
            .in3(N__17561),
            .lcout(\c0.m115_amcf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2_LC_9_23_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_2_LC_9_23_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \c0.tx.r_SM_Main_2_LC_9_23_5  (
            .in0(N__10469),
            .in1(N__10209),
            .in2(N__10408),
            .in3(N__10327),
            .lcout(\c0.tx.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21873),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_4_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_4_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_4_LC_9_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_6__RNO_0_4_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__11912),
            .in2(_gnd_net_),
            .in3(N__13016),
            .lcout(),
            .ltout(\c0.nextCRC16_3_3_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4_LC_9_24_1 .C_ON=1'b0;
    defparam \c0.data_out_6__4_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__4_LC_9_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__4_LC_9_24_1  (
            .in0(N__10160),
            .in1(N__12934),
            .in2(N__10163),
            .in3(N__12110),
            .lcout(\c0.data_out_6_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21880),
            .ce(N__17300),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_1_4_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_1_4_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_1_4_LC_9_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_1_4_LC_9_24_2  (
            .in0(N__12144),
            .in1(N__14657),
            .in2(N__13432),
            .in3(N__10812),
            .lcout(\c0.nextCRC16_3_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_4_LC_9_24_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_4_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_4_LC_9_24_3 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \c0.tx_data_RNO_0_4_LC_9_24_3  (
            .in0(N__19362),
            .in1(N__10154),
            .in2(N__15017),
            .in3(N__19204),
            .lcout(\c0.tx_data_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__6_LC_9_24_4 .C_ON=1'b0;
    defparam \c0.data_out_4__6_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__6_LC_9_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__6_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10610),
            .lcout(\c0.d_2_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21880),
            .ce(N__17300),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__1_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.data_out_5__1_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__1_LC_9_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__1_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10577),
            .lcout(\c0.d_2_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21880),
            .ce(N__17300),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_1_LC_9_24_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_1_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_1_LC_9_24_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_4_1_LC_9_24_6  (
            .in0(N__19203),
            .in1(N__12794),
            .in2(N__12148),
            .in3(N__19363),
            .lcout(),
            .ltout(\c0.tx_data_RNO_4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_1_LC_9_24_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_1_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_1_LC_9_24_7 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \c0.tx_data_RNO_2_1_LC_9_24_7  (
            .in0(N__16867),
            .in1(N__17562),
            .in2(N__10547),
            .in3(N__12635),
            .lcout(\c0.tx_data_1_0_i_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_3_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_3_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_3_LC_9_25_0 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \c0.tx_data_RNO_0_3_LC_9_25_0  (
            .in0(N__19402),
            .in1(N__19202),
            .in2(N__10520),
            .in3(N__10592),
            .lcout(\c0.tx_data_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_3_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_3_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_3_LC_9_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__RNO_0_3_LC_9_25_1  (
            .in0(N__11955),
            .in1(N__11076),
            .in2(_gnd_net_),
            .in3(N__12106),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__3_LC_9_25_2 .C_ON=1'b0;
    defparam \c0.data_out_6__3_LC_9_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__3_LC_9_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__3_LC_9_25_2  (
            .in0(N__10813),
            .in1(N__12770),
            .in2(N__10523),
            .in3(N__11258),
            .lcout(\c0.data_out_6_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21888),
            .ce(N__17299),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_7_LC_9_25_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_7_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_7_LC_9_25_5 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_3_7_LC_9_25_5  (
            .in0(N__19200),
            .in1(N__10511),
            .in2(N__12938),
            .in3(N__19403),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_7_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_7_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_7_LC_9_25_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_7_LC_9_25_6  (
            .in0(N__16842),
            .in1(N__17553),
            .in2(N__10493),
            .in3(N__10490),
            .lcout(\c0.tx_data_1_0_i_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_7_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_7_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_7_LC_9_25_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_4_7_LC_9_25_7  (
            .in0(N__19201),
            .in1(N__15286),
            .in2(N__15208),
            .in3(N__19401),
            .lcout(\c0.tx_data_RNO_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNI1DHT_19_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.d_2_RNI1DHT_19_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNI1DHT_19_LC_9_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNI1DHT_19_LC_9_26_1  (
            .in0(N__17418),
            .in1(N__17379),
            .in2(_gnd_net_),
            .in3(N__10591),
            .lcout(\c0.N_74 ),
            .ltout(\c0.N_74_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNITDBK1_47_LC_9_26_2 .C_ON=1'b0;
    defparam \c0.d_2_RNITDBK1_47_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNITDBK1_47_LC_9_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.d_2_RNITDBK1_47_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__15195),
            .in2(N__10595),
            .in3(N__15166),
            .lcout(\c0.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__3_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.data_out_2__3_LC_9_26_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__3_LC_9_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__3_LC_9_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13300),
            .lcout(\c0.d_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21898),
            .ce(),
            .sr(N__17343));
    defparam \c0.d_2_RNINVK01_8_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.d_2_RNINVK01_8_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNINVK01_8_LC_9_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNINVK01_8_LC_9_26_5  (
            .in0(N__10814),
            .in1(N__11249),
            .in2(_gnd_net_),
            .in3(N__11788),
            .lcout(\c0.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__0_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.data_out_1__0_LC_9_26_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__0_LC_9_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__0_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13299),
            .lcout(\c0.d_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21898),
            .ce(),
            .sr(N__17343));
    defparam \c0.data_0_LC_9_27_0 .C_ON=1'b1;
    defparam \c0.data_0_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_0_LC_9_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_0_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__11809),
            .in2(_gnd_net_),
            .in3(N__10580),
            .lcout(\c0.dataZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\c0.data_cry_0 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_1_LC_9_27_1 .C_ON=1'b1;
    defparam \c0.data_1_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_1_LC_9_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_1_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__10573),
            .in2(_gnd_net_),
            .in3(N__10562),
            .lcout(\c0.dataZ0Z_1 ),
            .ltout(),
            .carryin(\c0.data_cry_0 ),
            .carryout(\c0.data_cry_1 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_2_LC_9_27_2 .C_ON=1'b1;
    defparam \c0.data_2_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_2_LC_9_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_2_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__11113),
            .in2(_gnd_net_),
            .in3(N__10559),
            .lcout(\c0.dataZ0Z_2 ),
            .ltout(),
            .carryin(\c0.data_cry_1 ),
            .carryout(\c0.data_cry_2 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_3_LC_9_27_3 .C_ON=1'b1;
    defparam \c0.data_3_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_3_LC_9_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_3_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__11149),
            .in2(_gnd_net_),
            .in3(N__10556),
            .lcout(\c0.dataZ0Z_3 ),
            .ltout(),
            .carryin(\c0.data_cry_2 ),
            .carryout(\c0.data_cry_3 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_4_LC_9_27_4 .C_ON=1'b1;
    defparam \c0.data_4_LC_9_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_4_LC_9_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_4_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__11221),
            .in2(_gnd_net_),
            .in3(N__10553),
            .lcout(\c0.dataZ0Z_4 ),
            .ltout(),
            .carryin(\c0.data_cry_3 ),
            .carryout(\c0.data_cry_4 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_5_LC_9_27_5 .C_ON=1'b1;
    defparam \c0.data_5_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_5_LC_9_27_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_5_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__11281),
            .in2(_gnd_net_),
            .in3(N__10550),
            .lcout(\c0.dataZ0Z_5 ),
            .ltout(),
            .carryin(\c0.data_cry_4 ),
            .carryout(\c0.data_cry_5 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_6_LC_9_27_6 .C_ON=1'b1;
    defparam \c0.data_6_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_6_LC_9_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_6_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__11125),
            .in2(_gnd_net_),
            .in3(N__10667),
            .lcout(\c0.dataZ0Z_6 ),
            .ltout(),
            .carryin(\c0.data_cry_5 ),
            .carryout(\c0.data_cry_6 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_7_LC_9_27_7 .C_ON=1'b1;
    defparam \c0.data_7_LC_9_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_7_LC_9_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_7_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__11161),
            .in2(_gnd_net_),
            .in3(N__10664),
            .lcout(\c0.dataZ0Z_7 ),
            .ltout(),
            .carryin(\c0.data_cry_6 ),
            .carryout(\c0.data_cry_7 ),
            .clk(N__21906),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_8_LC_9_28_0 .C_ON=1'b1;
    defparam \c0.data_8_LC_9_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_8_LC_9_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_8_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__11869),
            .in2(_gnd_net_),
            .in3(N__10661),
            .lcout(\c0.dataZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\c0.data_cry_8 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_9_LC_9_28_1 .C_ON=1'b1;
    defparam \c0.data_9_LC_9_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_9_LC_9_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_9_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__11209),
            .in2(_gnd_net_),
            .in3(N__10658),
            .lcout(\c0.dataZ0Z_9 ),
            .ltout(),
            .carryin(\c0.data_cry_8 ),
            .carryout(\c0.data_cry_9 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_10_LC_9_28_2 .C_ON=1'b1;
    defparam \c0.data_10_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_10_LC_9_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_10_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__11137),
            .in2(_gnd_net_),
            .in3(N__10655),
            .lcout(\c0.dataZ0Z_10 ),
            .ltout(),
            .carryin(\c0.data_cry_9 ),
            .carryout(\c0.data_cry_10 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_11_LC_9_28_3 .C_ON=1'b1;
    defparam \c0.data_11_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_11_LC_9_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_11_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__10645),
            .in2(_gnd_net_),
            .in3(N__10634),
            .lcout(\c0.dataZ0Z_11 ),
            .ltout(),
            .carryin(\c0.data_cry_10 ),
            .carryout(\c0.data_cry_11 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_12_LC_9_28_4 .C_ON=1'b1;
    defparam \c0.data_12_LC_9_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_12_LC_9_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_12_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(N__10627),
            .in2(_gnd_net_),
            .in3(N__10616),
            .lcout(\c0.dataZ0Z_12 ),
            .ltout(),
            .carryin(\c0.data_cry_11 ),
            .carryout(\c0.data_cry_12 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_13_LC_9_28_5 .C_ON=1'b1;
    defparam \c0.data_13_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_13_LC_9_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_13_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(N__11269),
            .in2(_gnd_net_),
            .in3(N__10613),
            .lcout(\c0.dataZ0Z_13 ),
            .ltout(),
            .carryin(\c0.data_cry_12 ),
            .carryout(\c0.data_cry_13 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_14_LC_9_28_6 .C_ON=1'b1;
    defparam \c0.data_14_LC_9_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_14_LC_9_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_14_LC_9_28_6  (
            .in0(_gnd_net_),
            .in1(N__10606),
            .in2(_gnd_net_),
            .in3(N__10691),
            .lcout(\c0.dataZ0Z_14 ),
            .ltout(),
            .carryin(\c0.data_cry_13 ),
            .carryout(\c0.data_cry_14 ),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_15_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.data_15_LC_9_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_15_LC_9_28_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_15_LC_9_28_7  (
            .in0(_gnd_net_),
            .in1(N__12244),
            .in2(_gnd_net_),
            .in3(N__10688),
            .lcout(\c0.dataZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21914),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__1_LC_9_30_1 .C_ON=1'b0;
    defparam \c0.data_out_3__1_LC_9_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__1_LC_9_30_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__1_LC_9_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.d_2_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21929),
            .ce(),
            .sr(N__17339));
    defparam \c0.FRAME_MATCHER_i12_0_c_RNO_LC_10_16_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_0_c_RNO_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_0_c_RNO_LC_10_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_0_c_RNO_LC_10_16_3  (
            .in0(N__12166),
            .in1(N__12373),
            .in2(N__13585),
            .in3(N__15472),
            .lcout(\c0.i12_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__1_LC_10_16_4 .C_ON=1'b0;
    defparam \c0.data_in_0__1_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__1_LC_10_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__1_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15976),
            .lcout(\c0.data_in_0_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21829),
            .ce(N__22154),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__4_LC_10_16_6 .C_ON=1'b0;
    defparam \c0.data_in_0__4_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__4_LC_10_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__4_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14086),
            .lcout(\c0.data_in_0_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21829),
            .ce(N__22154),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_0_c_LC_10_17_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_0_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_0_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_0_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10685),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\c0.i12_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_1_c_LC_10_17_1 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_1_c_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_1_c_LC_10_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_1_c_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10709),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_0 ),
            .carryout(\c0.i12_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_2_c_LC_10_17_2 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_2_c_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_2_c_LC_10_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_2_c_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10676),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_1 ),
            .carryout(\c0.i12_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_3_c_LC_10_17_3 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_3_c_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_3_c_LC_10_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_3_c_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10700),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_2 ),
            .carryout(\c0.i12_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_4_c_LC_10_17_4 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_4_c_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_4_c_LC_10_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_4_c_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10742),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_3 ),
            .carryout(\c0.i12_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_5_c_LC_10_17_5 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_5_c_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_5_c_LC_10_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_5_c_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10721),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_4 ),
            .carryout(\c0.i12_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_6_c_LC_10_17_6 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_6_c_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_6_c_LC_10_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_6_c_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10733),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_5 ),
            .carryout(\c0.i12_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_LC_10_17_7 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i12_7_c_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_LC_10_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11198),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.i12_6 ),
            .carryout(\c0.i12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_THRU_LUT4_0_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.i12_THRU_LUT4_0_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_THRU_LUT4_0_LC_10_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.i12_THRU_LUT4_0_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10712),
            .lcout(\c0.i12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_3_LC_10_18_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_3_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_3_LC_10_18_2 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \c0.tx2_data_RNO_2_3_LC_10_18_2  (
            .in0(N__20334),
            .in1(N__17759),
            .in2(N__14111),
            .in3(N__17870),
            .lcout(\c0.tx2_data_1_iv_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_1_c_RNO_LC_10_18_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_1_c_RNO_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_1_c_RNO_LC_10_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_1_c_RNO_LC_10_18_3  (
            .in0(N__18297),
            .in1(N__15960),
            .in2(N__13923),
            .in3(N__17956),
            .lcout(\c0.i12_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_4  (
            .in0(N__15939),
            .in1(N__13863),
            .in2(N__16231),
            .in3(N__15423),
            .lcout(\c0.i12_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_3_LC_10_18_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_3_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_3_LC_10_18_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \c0.tx2_data_RNO_3_3_LC_10_18_5  (
            .in0(N__20902),
            .in1(N__13550),
            .in2(_gnd_net_),
            .in3(N__15406),
            .lcout(\c0.tx2_data_1_iv_3_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_18_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_18_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_18_6  (
            .in0(N__16258),
            .in1(N__13678),
            .in2(N__12409),
            .in3(N__16644),
            .lcout(\c0.i12_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__2_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.data_in_2__2_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__2_LC_10_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_2__2_LC_10_19_1  (
            .in0(N__16737),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_2_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21848),
            .ce(N__22156),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__3_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.data_in_2__3_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__3_LC_10_19_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_2__3_LC_10_19_2  (
            .in0(N__13804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_2_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21848),
            .ce(N__22156),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__5_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.data_in_2__5_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__5_LC_10_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__5_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11396),
            .lcout(\c0.data_in_2_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21848),
            .ce(N__22156),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__7_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.data_in_2__7_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__7_LC_10_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__7_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12331),
            .lcout(\c0.data_in_2_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21848),
            .ce(N__22156),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_19_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_19_7  (
            .in0(N__18666),
            .in1(N__13839),
            .in2(N__16741),
            .in3(N__13803),
            .lcout(\c0.i12_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__1_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.data_in_4__1_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__1_LC_10_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__1_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13819),
            .lcout(\c0.data_in_4_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__3_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.data_in_3__3_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__3_LC_10_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__3_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15844),
            .lcout(\c0.data_in_3_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__1_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.data_in_3__1_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__1_LC_10_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__1_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16078),
            .lcout(\c0.data_in_3_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__0_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.data_in_3__0_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__0_LC_10_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__0_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11320),
            .lcout(\c0.data_in_3_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__0_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.data_in_4__0_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__0_LC_10_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__0_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15913),
            .lcout(\c0.data_in_4_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__0_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.data_in_5__0_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__0_LC_10_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__0_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18782),
            .lcout(\c0.data_in_5_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__5_LC_10_20_7 .C_ON=1'b0;
    defparam \c0.data_in_7__5_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__5_LC_10_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__5_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10787),
            .lcout(\c0.data_in_7_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21855),
            .ce(N__22158),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_2_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_2_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_2_LC_10_21_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx2_data_RNO_1_2_LC_10_21_0  (
            .in0(N__22088),
            .in1(N__21992),
            .in2(N__19564),
            .in3(N__18923),
            .lcout(\c0.tx2_data_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_2_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_2_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_2_LC_10_21_1 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \c0.tx2_data_RNO_4_2_LC_10_21_1  (
            .in0(N__18921),
            .in1(N__16181),
            .in2(N__19539),
            .in3(N__16721),
            .lcout(\c0.tx2_data_RNO_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_2_LC_10_21_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_2_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_2_LC_10_21_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx2_data_RNO_0_2_LC_10_21_3  (
            .in0(N__18924),
            .in1(N__18411),
            .in2(N__19540),
            .in3(N__14165),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_2_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_2_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_2_LC_10_21_4 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \c0.tx2.r_Tx_Data_2_LC_10_21_4  (
            .in0(N__20357),
            .in1(N__10766),
            .in2(N__10760),
            .in3(N__10757),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21861),
            .ce(N__20745),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_1_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_1_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_1_LC_10_21_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx2_data_RNO_1_1_LC_10_21_6  (
            .in0(N__16670),
            .in1(N__19523),
            .in2(N__22040),
            .in3(N__18922),
            .lcout(\c0.tx2_data_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_3_LC_10_21_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_3_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_3_LC_10_21_7 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \c0.tx2.r_Tx_Data_3_LC_10_21_7  (
            .in0(N__14120),
            .in1(N__10751),
            .in2(N__12188),
            .in3(N__20356),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21861),
            .ce(N__20745),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_3_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_3_LC_10_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_3_LC_10_22_1 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.tx2.r_Clock_Count_3_LC_10_22_1  (
            .in0(N__14435),
            .in1(N__16436),
            .in2(N__14292),
            .in3(N__11555),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21866),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_7_LC_10_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_7_LC_10_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_7_LC_10_22_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.rx.r_Rx_Byte_7_LC_10_22_2  (
            .in0(N__10849),
            .in1(N__21122),
            .in2(N__18826),
            .in3(N__21218),
            .lcout(\c0.rx_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21866),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNI13HR_0_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNI13HR_0_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNI13HR_0_LC_10_22_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.tx2.r_SM_Main_RNI13HR_0_LC_10_22_4  (
            .in0(N__16366),
            .in1(N__14433),
            .in2(_gnd_net_),
            .in3(N__14354),
            .lcout(\c0.tx2.o_Tx_Serial12 ),
            .ltout(\c0.tx2.o_Tx_Serial12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_2_LC_10_22_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_2_LC_10_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_2_LC_10_22_5 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.tx2.r_Clock_Count_2_LC_10_22_5  (
            .in0(N__14434),
            .in1(N__11357),
            .in2(N__10829),
            .in3(N__16435),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21866),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_3_LC_10_22_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_3_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_3_LC_10_22_6 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx_data_RNO_3_3_LC_10_22_6  (
            .in0(N__12064),
            .in1(N__16516),
            .in2(N__19234),
            .in3(N__19411),
            .lcout(\c0.tx_data_RNO_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_2_LC_10_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_2_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_2_LC_10_22_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_2_LC_10_22_7  (
            .in0(N__21485),
            .in1(N__21391),
            .in2(_gnd_net_),
            .in3(N__21308),
            .lcout(\c0.rx.r_Rx_Bytece_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__6_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.data_out_0__6_LC_10_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__6_LC_10_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__6_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13249),
            .lcout(\c0.d_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21874),
            .ce(),
            .sr(N__17345));
    defparam \c0.data_out_2__4_LC_10_23_2 .C_ON=1'b0;
    defparam \c0.data_out_2__4_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__4_LC_10_23_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_2__4_LC_10_23_2  (
            .in0(N__13250),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21874),
            .ce(),
            .sr(N__17345));
    defparam \c0.data_out_2__6_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.data_out_2__6_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__6_LC_10_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__6_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13251),
            .lcout(\c0.d_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21874),
            .ce(),
            .sr(N__17345));
    defparam \c0.tx_data_RNO_4_6_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_6_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_6_LC_10_23_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx_data_RNO_4_6_LC_10_23_5  (
            .in0(N__15060),
            .in1(N__17540),
            .in2(_gnd_net_),
            .in3(N__10811),
            .lcout(),
            .ltout(\c0.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_6_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_6_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_6_LC_10_23_6 .LUT_INIT=16'b0001010111111111;
    LogicCell40 \c0.tx_data_RNO_2_6_LC_10_23_6  (
            .in0(N__11009),
            .in1(N__19162),
            .in2(N__11000),
            .in3(N__19412),
            .lcout(\c0.tx_data_1_0_i_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_6_LC_10_24_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_6_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_6_LC_10_24_0 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx_data_RNO_1_6_LC_10_24_0  (
            .in0(N__17563),
            .in1(N__14511),
            .in2(N__11748),
            .in3(N__16908),
            .lcout(),
            .ltout(\c0.tx_data_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_6_LC_10_24_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_6_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_6_LC_10_24_1 .LUT_INIT=16'b1011000110111011;
    LogicCell40 \c0.tx.r_Tx_Data_6_LC_10_24_1  (
            .in0(N__16869),
            .in1(N__10997),
            .in2(N__10988),
            .in3(N__16958),
            .lcout(\c0.tx.r_Tx_DataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21881),
            .ce(N__10941),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_2_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_2_LC_10_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_2_LC_10_24_2 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \c0.tx.r_Tx_Data_2_LC_10_24_2  (
            .in0(N__11615),
            .in1(N__16871),
            .in2(N__11021),
            .in3(N__14666),
            .lcout(\c0.tx.r_Tx_DataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21881),
            .ce(N__10941),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_7_LC_10_24_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_7_LC_10_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_7_LC_10_24_3 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \c0.tx.r_Tx_Data_7_LC_10_24_3  (
            .in0(N__16870),
            .in1(N__11045),
            .in2(N__14681),
            .in3(N__10961),
            .lcout(\c0.tx.r_Tx_DataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21881),
            .ce(N__10941),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_0_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_0_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_0_LC_10_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__RNO_0_0_LC_10_24_4  (
            .in0(N__11739),
            .in1(N__11256),
            .in2(_gnd_net_),
            .in3(N__17435),
            .lcout(\c0.nextCRC16_3_0_a2_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_24_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_24_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_24_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_4_LC_10_25_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_4_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_4_LC_10_25_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_1_4_LC_10_25_1  (
            .in0(N__19372),
            .in1(N__11171),
            .in2(N__19237),
            .in3(N__13092),
            .lcout(\c0.tx_data_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.data_out_6__1_LC_10_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__1_LC_10_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__1_LC_10_25_3  (
            .in0(N__11605),
            .in1(N__11849),
            .in2(N__11653),
            .in3(N__11078),
            .lcout(\c0.data_out_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21889),
            .ce(N__17295),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_5_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_5_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_5_LC_10_25_4 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.tx_data_RNO_0_5_LC_10_25_4  (
            .in0(N__11604),
            .in1(N__19373),
            .in2(N__12887),
            .in3(N__19218),
            .lcout(\c0.tx_data_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_7_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_7_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_7_LC_10_25_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_0_7_LC_10_25_5  (
            .in0(N__19374),
            .in1(N__12851),
            .in2(N__19235),
            .in3(N__11077),
            .lcout(\c0.tx_data_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_1_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_1_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_1_LC_10_25_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.tx_data_RNO_1_1_LC_10_25_6  (
            .in0(N__11956),
            .in1(N__19371),
            .in2(N__13127),
            .in3(N__19222),
            .lcout(\c0.tx_data_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_2_LC_10_25_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_2_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_2_LC_10_25_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx_data_RNO_1_2_LC_10_25_7  (
            .in0(N__19375),
            .in1(N__11102),
            .in2(N__19236),
            .in3(N__13003),
            .lcout(\c0.tx_data_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__4_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.data_out_1__4_LC_10_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__4_LC_10_26_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__4_LC_10_26_0  (
            .in0(N__13298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21899),
            .ce(),
            .sr(N__17342));
    defparam \c0.data_out_6__RNO_2_7_LC_10_26_1 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_2_7_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_2_7_LC_10_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_2_7_LC_10_26_1  (
            .in0(N__14603),
            .in1(N__12124),
            .in2(N__13011),
            .in3(N__12098),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_7_LC_10_26_2 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_7_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_7_LC_10_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_0_7_LC_10_26_2  (
            .in0(N__11957),
            .in1(N__11907),
            .in2(N__11012),
            .in3(N__13046),
            .lcout(\c0.nextCRC16_3_0_a2_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__2_LC_10_26_4 .C_ON=1'b0;
    defparam \c0.data_out_3__2_LC_10_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__2_LC_10_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__2_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.d_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21899),
            .ce(),
            .sr(N__17342));
    defparam \c0.tx_data_RNO_3_4_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_4_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_4_LC_10_26_5 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx_data_RNO_3_4_LC_10_26_5  (
            .in0(N__14860),
            .in1(N__16566),
            .in2(N__19233),
            .in3(N__19400),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_4_LC_10_26_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_4_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_4_LC_10_26_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \c0.tx_data_RNO_2_4_LC_10_26_6  (
            .in0(N__16843),
            .in1(N__17564),
            .in2(N__11189),
            .in3(N__11177),
            .lcout(\c0.tx_data_1_0_i_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_4_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_4_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_4_LC_10_26_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_4_4_LC_10_26_7  (
            .in0(N__19213),
            .in1(N__12125),
            .in2(N__12020),
            .in3(N__19399),
            .lcout(\c0.tx_data_RNO_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__4_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.data_out_7__4_LC_10_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__4_LC_10_27_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__4_LC_10_27_0  (
            .in0(N__12002),
            .in1(N__12838),
            .in2(N__14518),
            .in3(N__17378),
            .lcout(\c0.data_out_7_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__7_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.data_out_5__7_LC_10_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__7_LC_10_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__7_LC_10_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11162),
            .lcout(\c0.d_2_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__3_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.data_out_5__3_LC_10_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__3_LC_10_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__3_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11150),
            .lcout(\c0.d_2_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__2_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.data_out_4__2_LC_10_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__2_LC_10_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__2_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11138),
            .lcout(\c0.d_2_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__6_LC_10_27_4 .C_ON=1'b0;
    defparam \c0.data_out_5__6_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__6_LC_10_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__6_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11126),
            .lcout(\c0.d_2_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__2_LC_10_27_5 .C_ON=1'b0;
    defparam \c0.data_out_5__2_LC_10_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__2_LC_10_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__2_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11114),
            .lcout(\c0.d_2_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__2_LC_10_27_6 .C_ON=1'b0;
    defparam \c0.data_out_7__2_LC_10_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__2_LC_10_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__2_LC_10_27_6  (
            .in0(N__14557),
            .in1(N__14916),
            .in2(N__14519),
            .in3(N__12071),
            .lcout(\c0.data_out_7_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__5_LC_10_27_7 .C_ON=1'b0;
    defparam \c0.data_out_5__5_LC_10_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__5_LC_10_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__5_LC_10_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11282),
            .lcout(\c0.d_2_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21907),
            .ce(N__17293),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__5_LC_10_28_1 .C_ON=1'b0;
    defparam \c0.data_out_4__5_LC_10_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__5_LC_10_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__5_LC_10_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11270),
            .lcout(\c0.d_2_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21915),
            .ce(N__17291),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__4_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.data_out_5__4_LC_10_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__4_LC_10_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__4_LC_10_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11222),
            .lcout(\c0.d_2_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21915),
            .ce(N__17291),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__1_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.data_out_4__1_LC_10_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__1_LC_10_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__1_LC_10_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11210),
            .lcout(\c0.d_2_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21915),
            .ce(N__17291),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__6_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.data_out_1__6_LC_10_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__6_LC_10_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__6_LC_10_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13349),
            .lcout(\c0.d_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21923),
            .ce(),
            .sr(N__17338));
    defparam \c0.data_in_0__6_LC_11_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0__6_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__6_LC_11_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_0__6_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11418),
            .lcout(\c0.data_in_0_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21835),
            .ce(N__22157),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNO_LC_11_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNO_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNO_LC_11_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNO_LC_11_17_0  (
            .in0(N__11388),
            .in1(N__11436),
            .in2(N__13705),
            .in3(N__12324),
            .lcout(\c0.i12_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__4_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.data_in_3__4_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__4_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__4_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18511),
            .lcout(\c0.data_in_3_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__5_LC_11_17_2 .C_ON=1'b0;
    defparam \c0.data_in_3__5_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__5_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__5_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20009),
            .lcout(\c0.data_in_3_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__6_LC_11_17_3 .C_ON=1'b0;
    defparam \c0.data_in_3__6_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__6_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__6_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20555),
            .lcout(\c0.data_in_3_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__7_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.data_in_3__7_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__7_LC_11_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_3__7_LC_11_17_4  (
            .in0(N__18848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_3_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__6_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.data_in_2__6_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__6_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_2__6_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13701),
            .lcout(\c0.data_in_2_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__6_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.data_in_1__6_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__6_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_1__6_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18114),
            .lcout(\c0.data_in_1_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__4_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.data_in_4__4_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__4_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__4_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18719),
            .lcout(\c0.data_in_4_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21841),
            .ce(N__22153),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_2_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_2_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_2_LC_11_18_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \c0.wait_for_transmission_RNO_2_LC_11_18_0  (
            .in0(N__19493),
            .in1(N__20333),
            .in2(N__20901),
            .in3(N__18896),
            .lcout(\c0.N_72_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNI0CLC_0_0_LC_11_18_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNI0CLC_0_0_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNI0CLC_0_0_LC_11_18_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \c0.byte_transmit_counter2_RNI0CLC_0_0_LC_11_18_1  (
            .in0(N__20332),
            .in1(N__20861),
            .in2(_gnd_net_),
            .in3(N__19488),
            .lcout(),
            .ltout(\c0.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_active_RNIU1BT1_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.tx2_active_RNIU1BT1_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_active_RNIU1BT1_LC_11_18_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.tx2_active_RNIU1BT1_LC_11_18_2  (
            .in0(N__19758),
            .in1(N__12232),
            .in2(N__11294),
            .in3(N__18895),
            .lcout(\c0.N_247_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_0_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_0_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_0_LC_11_18_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.wait_for_transmission_RNO_0_LC_11_18_3  (
            .in0(N__12233),
            .in1(N__19759),
            .in2(_gnd_net_),
            .in3(N__11291),
            .lcout(),
            .ltout(\c0.N_249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_LC_11_18_4 .SEQ_MODE=4'b1001;
    defparam \c0.wait_for_transmission_LC_11_18_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \c0.wait_for_transmission_LC_11_18_4  (
            .in0(N__19807),
            .in1(N__11300),
            .in2(N__11285),
            .in3(N__12284),
            .lcout(\c0.wait_for_transmissionZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21849),
            .ce(),
            .sr(N__20045));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_11_18_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_11_18_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_11_18_5  (
            .in0(N__19793),
            .in1(N__17725),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_frame_0__0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_0_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_0_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_0_LC_11_18_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \c0.tx2_data_RNO_0_0_LC_11_18_6  (
            .in0(N__18910),
            .in1(N__15601),
            .in2(N__19502),
            .in3(N__15902),
            .lcout(\c0.tx2_data_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_1_LC_11_18_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_1_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_1_LC_11_18_7 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \c0.tx2_data_RNO_0_1_LC_11_18_7  (
            .in0(N__18897),
            .in1(N__15782),
            .in2(N__16067),
            .in3(N__19492),
            .lcout(\c0.tx2_data_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIM5UG_0_19_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIM5UG_0_19_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIM5UG_0_19_LC_11_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIM5UG_0_19_LC_11_19_0  (
            .in0(N__15595),
            .in1(N__15401),
            .in2(N__19961),
            .in3(N__17903),
            .lcout(\c0.g3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__0_LC_11_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__0_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__0_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__0_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11321),
            .lcout(\c0.d_4_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21856),
            .ce(N__21594),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_4_LC_11_19_2 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_4_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_4_LC_11_19_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.wait_for_transmission_RNO_4_LC_11_19_2  (
            .in0(N__17744),
            .in1(N__18143),
            .in2(N__18536),
            .in3(N__17724),
            .lcout(\c0.g0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIM5UG_19_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIM5UG_19_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIM5UG_19_LC_11_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIM5UG_19_LC_11_19_3  (
            .in0(N__17905),
            .in1(N__19954),
            .in2(N__15407),
            .in3(N__15597),
            .lcout(\c0.g3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_5_LC_11_19_4 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_5_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_5_LC_11_19_4 .LUT_INIT=16'b0001001010000100;
    LogicCell40 \c0.wait_for_transmission_RNO_5_LC_11_19_4  (
            .in0(N__15869),
            .in1(N__17691),
            .in2(N__13565),
            .in3(N__17660),
            .lcout(),
            .ltout(\c0.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_1_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_1_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_1_LC_11_19_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \c0.wait_for_transmission_RNO_1_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__11345),
            .in2(N__11309),
            .in3(N__11306),
            .lcout(\c0.byte_transmit_counter2_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_6_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_6_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_6_LC_11_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.wait_for_transmission_RNO_6_LC_11_19_6  (
            .in0(N__15596),
            .in1(N__15402),
            .in2(N__19962),
            .in3(N__17904),
            .lcout(),
            .ltout(\c0.g3_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_3_LC_11_19_7 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_3_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_3_LC_11_19_7 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \c0.wait_for_transmission_RNO_3_LC_11_19_7  (
            .in0(N__15698),
            .in1(N__15734),
            .in2(N__11348),
            .in3(N__15818),
            .lcout(\c0.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__2_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.data_in_4__2_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__2_LC_11_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__2_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11371),
            .lcout(\c0.data_in_4_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__3_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.data_in_6__3_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__3_LC_11_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__3_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14065),
            .lcout(\c0.data_in_6_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__2_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.data_in_3__2_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__2_LC_11_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_3__2_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13939),
            .lcout(\c0.data_in_3_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__1_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.data_in_5__1_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__1_LC_11_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__1_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18809),
            .lcout(\c0.data_in_5_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__2_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.data_in_5__2_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__2_LC_11_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__2_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22115),
            .lcout(\c0.data_in_5_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__1_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.data_in_7__1_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__1_LC_11_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__1_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11339),
            .lcout(\c0.data_in_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__3_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.data_in_4__3_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__3_LC_11_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__3_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14446),
            .lcout(\c0.data_in_4_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__3_LC_11_20_7 .C_ON=1'b0;
    defparam \c0.data_in_5__3_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__3_LC_11_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__3_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20631),
            .lcout(\c0.data_in_5_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21862),
            .ce(N__22159),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIBANL_28_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIBANL_28_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIBANL_28_LC_11_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIBANL_28_LC_11_21_0  (
            .in0(N__17015),
            .in1(N__18956),
            .in2(N__14008),
            .in3(N__12598),
            .lcout(\c0.un1_data_in_7__2_0_a2_0_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__4_LC_11_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__4_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__4_LC_11_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__4_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11444),
            .lcout(\c0.d_4_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21867),
            .ce(N__21599),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__6_LC_11_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__6_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__6_LC_11_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__6_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11420),
            .lcout(\c0.d_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21867),
            .ce(N__21599),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__5_LC_11_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__5_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__5_LC_11_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__5_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11395),
            .lcout(\c0.d_4_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21867),
            .ce(N__21599),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI7BIA_29_LC_11_21_4 .C_ON=1'b0;
    defparam \c0.d_4_RNI7BIA_29_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI7BIA_29_LC_11_21_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.d_4_RNI7BIA_29_LC_11_21_4  (
            .in0(N__22200),
            .in1(_gnd_net_),
            .in2(N__17023),
            .in3(N__17127),
            .lcout(\c0.un1_data_in_6__7_0_a2_17_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__4_LC_11_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__4_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__4_LC_11_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__4_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18718),
            .lcout(\c0.d_4_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21867),
            .ce(N__21599),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__2_LC_11_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__2_LC_11_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__2_LC_11_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__2_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11372),
            .lcout(\c0.d_4_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21867),
            .ce(N__21599),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_RNO_0_0_LC_11_22_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count_RNO_0_0_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count_RNO_0_0_LC_11_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx2.r_Clock_Count_RNO_0_0_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__11528),
            .in2(N__11549),
            .in3(N__11548),
            .lcout(\c0.tx2.r_Clock_Count_RNO_0_0_0 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\c0.tx2.un1_r_Clock_Count_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_RNO_0_1_LC_11_22_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count_RNO_0_1_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count_RNO_0_1_LC_11_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx2.r_Clock_Count_RNO_0_1_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__11498),
            .in2(_gnd_net_),
            .in3(N__11360),
            .lcout(\c0.tx2.r_Clock_Count_RNO_0_0_1 ),
            .ltout(),
            .carryin(\c0.tx2.un1_r_Clock_Count_cry_0 ),
            .carryout(\c0.tx2.un1_r_Clock_Count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_RNO_0_2_LC_11_22_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count_RNO_0_2_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count_RNO_0_2_LC_11_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.tx2.r_Clock_Count_RNO_0_2_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__11480),
            .in2(_gnd_net_),
            .in3(N__11351),
            .lcout(\c0.tx2.r_Clock_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\c0.tx2.un1_r_Clock_Count_cry_1 ),
            .carryout(\c0.tx2.un1_r_Clock_Count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_RNO_0_3_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_RNO_0_3_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count_RNO_0_3_LC_11_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.tx2.r_Clock_Count_RNO_0_3_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__11462),
            .in2(_gnd_net_),
            .in3(N__11558),
            .lcout(\c0.tx2.r_Clock_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNINID81_0_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNINID81_0_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNINID81_0_LC_11_22_4 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.tx2.r_SM_Main_RNINID81_0_LC_11_22_4  (
            .in0(N__16365),
            .in1(N__14350),
            .in2(N__14432),
            .in3(N__16420),
            .lcout(\c0.tx2.r_Clock_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_11_22_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_11_22_5  (
            .in0(N__13348),
            .in1(N__11527),
            .in2(_gnd_net_),
            .in3(N__11510),
            .lcout(\c0.tx2.r_Clock_Count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_0_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_0_LC_11_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_0_LC_11_22_6 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \c0.tx2.r_Clock_Count_0_LC_11_22_6  (
            .in0(N__14419),
            .in1(N__11534),
            .in2(N__14293),
            .in3(N__16421),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count_1_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count_1_LC_11_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count_1_LC_11_22_7 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.tx2.r_Clock_Count_1_LC_11_22_7  (
            .in0(N__16422),
            .in1(N__14420),
            .in2(N__14291),
            .in3(N__11516),
            .lcout(\c0.tx2.r_Clock_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21875),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_LC_11_23_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_0_c_LC_11_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_0_c_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__11509),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\c0.tx2.r_Clock_Count12_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_11_23_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_11_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__11486),
            .in2(N__13301),
            .in3(N__11497),
            .lcout(\c0.tx2.r_Clock_Count_i_1 ),
            .ltout(),
            .carryin(\c0.tx2.r_Clock_Count12_cry_0 ),
            .carryout(\c0.tx2.r_Clock_Count12_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_11_23_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_11_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__11468),
            .in2(N__13303),
            .in3(N__11479),
            .lcout(\c0.tx2.r_Clock_Count_i_2 ),
            .ltout(),
            .carryin(\c0.tx2.r_Clock_Count12_cry_1 ),
            .carryout(\c0.tx2.r_Clock_Count12_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_11_23_3 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_11_23_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_11_23_3  (
            .in0(N__11461),
            .in1(N__11450),
            .in2(N__13302),
            .in3(_gnd_net_),
            .lcout(\c0.tx2.r_Clock_Count_i_3 ),
            .ltout(),
            .carryin(\c0.tx2.r_Clock_Count12_cry_2 ),
            .carryout(\c0.tx2.r_Clock_Count12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_11_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11657),
            .lcout(\c0.tx2.r_Clock_Count12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__1_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.data_out_1__1_LC_11_23_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__1_LC_11_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_1__1_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13260),
            .lcout(\c0.d_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21882),
            .ce(),
            .sr(N__17344));
    defparam \c0.data_out_1__2_LC_11_23_7 .C_ON=1'b0;
    defparam \c0.data_out_1__2_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__2_LC_11_23_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__2_LC_11_23_7  (
            .in0(N__13261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21882),
            .ce(),
            .sr(N__17344));
    defparam \c0.data_out_6__2_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.data_out_6__2_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__2_LC_11_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__2_LC_11_24_0  (
            .in0(N__12932),
            .in1(N__12790),
            .in2(N__11762),
            .in3(N__11654),
            .lcout(\c0.data_out_6_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21890),
            .ce(N__17296),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_2_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_2_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_2_LC_11_24_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx_data_RNO_0_2_LC_11_24_2  (
            .in0(N__15106),
            .in1(N__19185),
            .in2(N__11624),
            .in3(N__19370),
            .lcout(\c0.tx_data_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__7_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.data_out_7__7_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__7_LC_11_24_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__7_LC_11_24_5  (
            .in0(N__11709),
            .in1(N__11609),
            .in2(N__16478),
            .in3(N__11675),
            .lcout(\c0.data_out_7_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21890),
            .ce(N__17296),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_0_LC_11_25_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_0_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_0_LC_11_25_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \c0.tx_data_RNO_4_0_LC_11_25_0  (
            .in0(N__15135),
            .in1(N__16808),
            .in2(N__12105),
            .in3(N__17521),
            .lcout(),
            .ltout(\c0.tx_data_1_iv_i_m2_0_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_0_LC_11_25_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_0_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_0_LC_11_25_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx_data_RNO_3_0_LC_11_25_1  (
            .in0(N__16809),
            .in1(N__11798),
            .in2(N__11576),
            .in3(N__11822),
            .lcout(),
            .ltout(\c0.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_0_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_0_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_0_LC_11_25_2 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \c0.tx_data_RNO_2_0_LC_11_25_2  (
            .in0(_gnd_net_),
            .in1(N__19396),
            .in2(N__11573),
            .in3(N__19214),
            .lcout(\c0.tx_data_1_iv_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__0_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.data_out_6__0_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__0_LC_11_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__0_LC_11_25_3  (
            .in0(N__15023),
            .in1(N__11723),
            .in2(N__11858),
            .in3(N__11848),
            .lcout(\c0.data_out_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21900),
            .ce(N__17294),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__0_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.data_out_5__0_LC_11_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__0_LC_11_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_5__0_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11816),
            .lcout(\c0.d_2_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21900),
            .ce(N__17294),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__0_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.data_out_7__0_LC_11_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__0_LC_11_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__0_LC_11_25_6  (
            .in0(N__11768),
            .in1(N__12701),
            .in2(N__13190),
            .in3(N__13147),
            .lcout(\c0.data_out_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21900),
            .ce(N__17294),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_0_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_0_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_0_LC_11_26_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx_data_RNO_0_0_LC_11_26_0  (
            .in0(N__11792),
            .in1(N__17565),
            .in2(N__13064),
            .in3(N__16909),
            .lcout(\c0.tx_data_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_0_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_0_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_0_LC_11_26_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.data_out_7__RNO_0_0_LC_11_26_1  (
            .in0(N__15098),
            .in1(_gnd_net_),
            .in2(N__15246),
            .in3(N__12034),
            .lcout(\c0.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_0_2_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_0_2_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_0_2_LC_11_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__RNO_0_2_LC_11_26_2  (
            .in0(N__16568),
            .in1(N__11750),
            .in2(_gnd_net_),
            .in3(N__13418),
            .lcout(\c0.nextCRC16_3_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_2_0_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_2_0_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_2_0_LC_11_26_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.data_out_7__RNO_2_0_LC_11_26_4  (
            .in0(N__15308),
            .in1(_gnd_net_),
            .in2(N__15062),
            .in3(N__12828),
            .lcout(\c0.nextCRC16_3_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIQ3DA1_20_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.d_2_RNIQ3DA1_20_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIQ3DA1_20_LC_11_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIQ3DA1_20_LC_11_26_5  (
            .in0(N__11749),
            .in1(N__15021),
            .in2(N__13425),
            .in3(N__11716),
            .lcout(),
            .ltout(\c0.nextCRC16_3_0_a2_6_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIKDAK6_20_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.d_2_RNIKDAK6_20_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIKDAK6_20_LC_11_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIKDAK6_20_LC_11_26_6  (
            .in0(N__12769),
            .in1(N__11687),
            .in2(N__11678),
            .in3(N__11671),
            .lcout(\c0.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIM3JT_12_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.d_2_RNIM3JT_12_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIM3JT_12_LC_11_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIM3JT_12_LC_11_26_7  (
            .in0(N__12149),
            .in1(N__12123),
            .in2(_gnd_net_),
            .in3(N__12097),
            .lcout(\c0.N_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__RNO_1_7_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.data_out_6__RNO_1_7_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__RNO_1_7_LC_11_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__RNO_1_7_LC_11_27_0  (
            .in0(N__12967),
            .in1(N__14550),
            .in2(N__14921),
            .in3(N__14501),
            .lcout(\c0.nextCRC16_3_0_a2_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_2_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_2_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_2_LC_11_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_0_2_LC_11_27_1  (
            .in0(N__15055),
            .in1(N__12820),
            .in2(N__11996),
            .in3(N__13070),
            .lcout(\c0.nextCRC16_3_0_a2_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNI6EK01_3_LC_11_27_3 .C_ON=1'b0;
    defparam \c0.d_2_RNI6EK01_3_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNI6EK01_3_LC_11_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNI6EK01_3_LC_11_27_3  (
            .in0(N__15126),
            .in1(N__15350),
            .in2(_gnd_net_),
            .in3(N__12065),
            .lcout(\c0.N_75 ),
            .ltout(\c0.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIJ2812_44_LC_11_27_4 .C_ON=1'b0;
    defparam \c0.d_2_RNIJ2812_44_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIJ2812_44_LC_11_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIJ2812_44_LC_11_27_4  (
            .in0(N__15247),
            .in1(N__15105),
            .in2(N__12023),
            .in3(N__12013),
            .lcout(\c0.N_95 ),
            .ltout(\c0.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIJDOU2_14_LC_11_27_5 .C_ON=1'b0;
    defparam \c0.d_2_RNIJDOU2_14_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIJDOU2_14_LC_11_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIJDOU2_14_LC_11_27_5  (
            .in0(N__15056),
            .in1(N__11991),
            .in2(N__11960),
            .in3(N__12821),
            .lcout(\c0.nextCRC16_3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNII92R1_27_LC_11_27_7 .C_ON=1'b0;
    defparam \c0.d_2_RNII92R1_27_LC_11_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNII92R1_27_LC_11_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNII92R1_27_LC_11_27_7  (
            .in0(N__11954),
            .in1(N__11911),
            .in2(N__14731),
            .in3(N__14569),
            .lcout(\c0.N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__0_LC_11_28_2 .C_ON=1'b0;
    defparam \c0.data_out_4__0_LC_11_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__0_LC_11_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__0_LC_11_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11873),
            .lcout(\c0.d_2_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21924),
            .ce(N__17289),
            .sr(_gnd_net_));
    defparam \c0.data_out_4__7_LC_11_28_3 .C_ON=1'b0;
    defparam \c0.data_out_4__7_LC_11_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_4__7_LC_11_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_4__7_LC_11_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12248),
            .lcout(\c0.d_2_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21924),
            .ce(N__17289),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_LC_12_16_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_LC_12_16_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.tx2.r_Tx_Active_LC_12_16_6  (
            .in0(N__20749),
            .in1(N__12231),
            .in2(_gnd_net_),
            .in3(N__12647),
            .lcout(\c0.tx2_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_5_7_LC_12_17_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_5_7_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_5_7_LC_12_17_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \c0.tx2_data_RNO_5_7_LC_12_17_0  (
            .in0(N__20924),
            .in1(N__12206),
            .in2(_gnd_net_),
            .in3(N__18218),
            .lcout(\c0.tx2_data_1_iv_5_1_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_7_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_7_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_7_LC_12_17_1 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \c0.tx2_data_RNO_4_7_LC_12_17_1  (
            .in0(N__18044),
            .in1(N__20925),
            .in2(N__20411),
            .in3(N__18335),
            .lcout(),
            .ltout(\c0.tx2_data_1_iv_5_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_7_LC_12_17_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_7_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_7_LC_12_17_2 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \c0.tx2_data_RNO_2_7_LC_12_17_2  (
            .in0(N__12215),
            .in1(N__20408),
            .in2(N__12209),
            .in3(N__20339),
            .lcout(\c0.tx2_data_1_iv_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__7_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__7_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__7_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__7_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22205),
            .lcout(\c0.data_in_frame_6_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21850),
            .ce(N__21586),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_3_LC_12_17_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_3_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_3_LC_12_17_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.tx2_data_RNO_1_3_LC_12_17_4  (
            .in0(N__12200),
            .in1(N__20407),
            .in2(_gnd_net_),
            .in3(N__20338),
            .lcout(\c0.tx2_data_1_iv_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__3_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__3_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__3_LC_12_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__3_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12173),
            .lcout(\c0.d_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21850),
            .ce(N__21586),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNI94LS6_LC_12_18_0 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNI94LS6_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNI94LS6_LC_12_18_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \c0.wait_for_transmission_RNI94LS6_LC_12_18_0  (
            .in0(N__19792),
            .in1(N__12155),
            .in2(_gnd_net_),
            .in3(N__13478),
            .lcout(\c0.wait_for_transmission_RNI94LSZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIT2KP_20_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIT2KP_20_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIT2KP_20_LC_12_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIT2KP_20_LC_12_18_1  (
            .in0(N__19726),
            .in1(N__18334),
            .in2(N__18781),
            .in3(N__14158),
            .lcout(),
            .ltout(\c0.un1_data_in_6__0_0_a2_5_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI2LMH1_6_LC_12_18_2 .C_ON=1'b0;
    defparam \c0.d_4_RNI2LMH1_6_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI2LMH1_6_LC_12_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI2LMH1_6_LC_12_18_2  (
            .in0(N__18004),
            .in1(N__18182),
            .in2(N__12308),
            .in3(N__15460),
            .lcout(\c0.un1_data_in_6__0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI4CPT_18_LC_12_18_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI4CPT_18_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI4CPT_18_LC_12_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI4CPT_18_LC_12_18_3  (
            .in0(N__13545),
            .in1(N__16180),
            .in2(N__21980),
            .in3(N__16063),
            .lcout(),
            .ltout(\c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIHG3O1_16_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIHG3O1_16_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIHG3O1_16_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.d_4_RNIHG3O1_16_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__12422),
            .in2(N__12305),
            .in3(N__12467),
            .lcout(),
            .ltout(\c0.un1_data_in_7__4_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIK1Q66_10_LC_12_18_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIK1Q66_10_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIK1Q66_10_LC_12_18_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \c0.d_4_RNIK1Q66_10_LC_12_18_5  (
            .in0(N__14132),
            .in1(N__15995),
            .in2(N__12302),
            .in3(N__12299),
            .lcout(\c0.wait_for_transmission4_12_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIF73E2_14_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIF73E2_14_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIF73E2_14_LC_12_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIF73E2_14_LC_12_19_0  (
            .in0(N__17184),
            .in1(N__16717),
            .in2(N__14024),
            .in3(N__13783),
            .lcout(),
            .ltout(\c0.d_4_RNIF73E2Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIMKFE3_14_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIMKFE3_14_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIMKFE3_14_LC_12_19_1 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.d_4_RNIMKFE3_14_LC_12_19_1  (
            .in0(N__12434),
            .in1(_gnd_net_),
            .in2(N__12293),
            .in3(N__14803),
            .lcout(),
            .ltout(\c0.d_4_RNIMKFE3Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIOL9I8_10_LC_12_19_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIOL9I8_10_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIOL9I8_10_LC_12_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.d_4_RNIOL9I8_10_LC_12_19_2  (
            .in0(N__15550),
            .in1(N__16103),
            .in2(N__12290),
            .in3(N__15811),
            .lcout(),
            .ltout(\c0.un1_data_in_6__7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIB4H0M_43_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIB4H0M_43_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIB4H0M_43_LC_12_19_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.d_4_RNIB4H0M_43_LC_12_19_3  (
            .in0(N__17627),
            .in1(N__17605),
            .in2(N__12287),
            .in3(N__17587),
            .lcout(\c0.wait_for_transmission4_12 ),
            .ltout(\c0.wait_for_transmission4_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI61KS81_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI61KS81_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI61KS81_LC_12_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNI61KS81_LC_12_19_4  (
            .in0(N__12265),
            .in1(N__13442),
            .in2(N__12251),
            .in3(N__13454),
            .lcout(\c0.tx2_transmit_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIFCG72_32_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIFCG72_32_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIFCG72_32_LC_12_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.d_4_RNIFCG72_32_LC_12_19_5  (
            .in0(N__15594),
            .in1(N__12386),
            .in2(_gnd_net_),
            .in3(N__12392),
            .lcout(\c0.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI46QL_16_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI46QL_16_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI46QL_16_LC_12_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI46QL_16_LC_12_20_0  (
            .in0(N__13635),
            .in1(N__17128),
            .in2(N__13969),
            .in3(N__12491),
            .lcout(\c0.un1_data_in_7__4_0_a2_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__2_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__2_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__2_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__2_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12413),
            .lcout(\c0.d_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21868),
            .ce(N__21595),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNID6K21_0_15_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNID6K21_0_15_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNID6K21_0_15_LC_12_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNID6K21_0_15_LC_12_20_2  (
            .in0(N__17901),
            .in1(N__12487),
            .in2(N__17941),
            .in3(N__12600),
            .lcout(\c0.d_4_RNID6K21_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNID6K21_15_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.d_4_RNID6K21_15_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNID6K21_15_LC_12_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.d_4_RNID6K21_15_LC_12_20_3  (
            .in0(N__12599),
            .in1(N__17937),
            .in2(N__12496),
            .in3(N__17902),
            .lcout(\c0.d_4_RNID6K21Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__1_LC_12_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__1_LC_12_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__1_LC_12_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__1_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12380),
            .lcout(\c0.d_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21868),
            .ce(N__21595),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__7_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__7_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__7_LC_12_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__7_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12362),
            .lcout(\c0.d_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21868),
            .ce(N__21595),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__7_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__7_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__7_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__7_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12332),
            .lcout(\c0.d_4_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21868),
            .ce(N__21595),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI9UF4_32_LC_12_20_7 .C_ON=1'b0;
    defparam \c0.d_4_RNI9UF4_32_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI9UF4_32_LC_12_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_4_RNI9UF4_32_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__15593),
            .in2(_gnd_net_),
            .in3(N__17900),
            .lcout(\c0.N_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__RNI74HC_1_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.data_in_7__RNI74HC_1_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_7__RNI74HC_1_LC_12_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_in_7__RNI74HC_1_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__22056),
            .in2(_gnd_net_),
            .in3(N__17125),
            .lcout(),
            .ltout(\c0.un1_data_in_7__1_0_a2_24_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI716J_16_LC_12_21_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI716J_16_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI716J_16_LC_12_21_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.d_4_RNI716J_16_LC_12_21_1  (
            .in0(N__18412),
            .in1(N__13642),
            .in2(N__12503),
            .in3(N__17171),
            .lcout(\c0.wait_for_transmission4_13_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNID6C91_1_LC_12_21_3 .C_ON=1'b0;
    defparam \c0.d_4_RNID6C91_1_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNID6C91_1_LC_12_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNID6C91_1_LC_12_21_3  (
            .in0(N__12492),
            .in1(N__12463),
            .in2(N__15723),
            .in3(N__12601),
            .lcout(),
            .ltout(\c0.un1_data_in_7__1_0_a2_24_a2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI8S283_14_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.d_4_RNI8S283_14_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI8S283_14_LC_12_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI8S283_14_LC_12_21_4  (
            .in0(N__14009),
            .in1(N__12452),
            .in2(N__12446),
            .in3(N__12440),
            .lcout(\c0.wait_for_transmission4_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIJ6E4_27_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIJ6E4_27_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIJ6E4_27_LC_12_21_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.d_4_RNIJ6E4_27_LC_12_21_5  (
            .in0(N__17798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18957),
            .lcout(),
            .ltout(\c0.un1_data_in_7__1_0_a2_24_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIVMA91_17_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIVMA91_17_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIVMA91_17_LC_12_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIVMA91_17_LC_12_21_6  (
            .in0(N__13546),
            .in1(N__13738),
            .in2(N__12443),
            .in3(N__15618),
            .lcout(\c0.un1_data_in_7__1_0_a2_24_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNITCRC_29_LC_12_21_7 .C_ON=1'b0;
    defparam \c0.d_4_RNITCRC_29_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNITCRC_29_LC_12_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNITCRC_29_LC_12_21_7  (
            .in0(N__17126),
            .in1(N__22201),
            .in2(N__18423),
            .in3(N__17022),
            .lcout(\c0.d_4_RNITCRCZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_0_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_0_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_0_LC_12_22_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \c0.tx2_data_RNO_4_0_LC_12_22_0  (
            .in0(N__18928),
            .in1(N__18648),
            .in2(N__19574),
            .in3(N__13643),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_0_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_0_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_0_LC_12_22_1 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \c0.tx2_data_RNO_2_0_LC_12_22_1  (
            .in0(N__20342),
            .in1(N__13601),
            .in2(N__12425),
            .in3(N__20941),
            .lcout(),
            .ltout(\c0.tx2_data_1_0_i_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_0_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_0_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_0_LC_12_22_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \c0.tx2.r_Tx_Data_0_LC_12_22_2  (
            .in0(N__12539),
            .in1(N__12623),
            .in2(N__12611),
            .in3(N__20344),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21883),
            .ce(N__20741),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_1_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_1_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_1_LC_12_22_3 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2_data_RNO_3_1_LC_12_22_3  (
            .in0(N__19572),
            .in1(N__18257),
            .in2(N__12608),
            .in3(N__18927),
            .lcout(),
            .ltout(\c0.tx2_data_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_1_LC_12_22_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_1_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_1_LC_12_22_4 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \c0.tx2_data_RNO_2_1_LC_12_22_4  (
            .in0(N__20942),
            .in1(N__12545),
            .in2(N__12575),
            .in3(N__20343),
            .lcout(),
            .ltout(\c0.tx2_data_1_0_i_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_1_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_1_LC_12_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_1_LC_12_22_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \c0.tx2.r_Tx_Data_1_LC_12_22_5  (
            .in0(N__20345),
            .in1(N__12572),
            .in2(N__12560),
            .in3(N__12557),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21883),
            .ce(N__20741),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_1_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_1_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_1_LC_12_22_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \c0.tx2_data_RNO_4_1_LC_12_22_6  (
            .in0(N__18926),
            .in1(N__13739),
            .in2(N__19573),
            .in3(N__16031),
            .lcout(\c0.tx2_data_RNO_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_0_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_0_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_0_LC_12_22_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx2_data_RNO_1_0_LC_12_22_7  (
            .in0(N__16754),
            .in1(N__19568),
            .in2(N__16583),
            .in3(N__18929),
            .lcout(\c0.tx2_data_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_2_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_2_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_2_LC_12_23_0 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_2_LC_12_23_0  (
            .in0(N__16306),
            .in1(N__12533),
            .in2(N__14744),
            .in3(N__12515),
            .lcout(\c0.tx2.N_349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_4_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_4_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_4_LC_12_23_1 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_4_LC_12_23_1  (
            .in0(N__12521),
            .in1(N__14225),
            .in2(N__20768),
            .in3(N__16304),
            .lcout(\c0.tx2.r_Tx_Data_pmux_3_i_m2_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_3_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_3_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_3_LC_12_23_2 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_3_LC_12_23_2  (
            .in0(N__16305),
            .in1(N__16982),
            .in2(N__14233),
            .in3(N__12509),
            .lcout(),
            .ltout(\c0.tx2.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_1_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_1_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_1_LC_12_23_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_1_LC_12_23_3  (
            .in0(N__17081),
            .in1(N__12695),
            .in2(N__12683),
            .in3(N__16307),
            .lcout(),
            .ltout(\c0.tx2.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_RNO_0_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_RNO_0_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_RNO_0_LC_12_23_4 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \c0.tx2.o_Tx_Serial_RNO_0_LC_12_23_4  (
            .in0(N__16461),
            .in1(N__12680),
            .in2(N__12674),
            .in3(N__14343),
            .lcout(),
            .ltout(\c0.tx2.N_279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_LC_12_23_5 .SEQ_MODE=4'b1001;
    defparam \c0.tx2.o_Tx_Serial_LC_12_23_5 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \c0.tx2.o_Tx_Serial_LC_12_23_5  (
            .in0(N__14408),
            .in1(N__12664),
            .in2(N__12671),
            .in3(N__16349),
            .lcout(PIN_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21891),
            .ce(),
            .sr(N__14287));
    defparam \c0.tx2.r_SM_Main_RNINID81_0_0_LC_12_23_7 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNINID81_0_0_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNINID81_0_0_LC_12_23_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.tx2.r_SM_Main_RNINID81_0_0_LC_12_23_7  (
            .in0(N__14342),
            .in1(N__16348),
            .in2(N__14429),
            .in3(N__16423),
            .lcout(\c0.tx2.r_Tx_Active_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_2_LC_12_24_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.tx2.r_SM_Main_2_LC_12_24_1  (
            .in0(N__16352),
            .in1(N__14349),
            .in2(N__14431),
            .in3(N__16434),
            .lcout(\c0.tx2.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21901),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_1_LC_12_24_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_1_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_1_LC_12_24_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_3_1_LC_12_24_2  (
            .in0(N__19168),
            .in1(N__14889),
            .in2(N__17392),
            .in3(N__19322),
            .lcout(\c0.tx_data_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_0_LC_12_24_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_0_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_0_LC_12_24_3 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \c0.tx2.r_SM_Main_7_1_0__m5_0_0_LC_12_24_3  (
            .in0(N__14409),
            .in1(N__14347),
            .in2(N__20715),
            .in3(N__16432),
            .lcout(),
            .ltout(\c0.tx2.m5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_0_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_0_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_0_LC_12_24_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \c0.tx2.r_SM_Main_0_LC_12_24_4  (
            .in0(N__14234),
            .in1(N__16350),
            .in2(N__12626),
            .in3(N__14300),
            .lcout(\c0.tx2.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21901),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_1_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_1_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_1_LC_12_24_5 .LUT_INIT=16'b0000101000000110;
    LogicCell40 \c0.tx2.r_SM_Main_1_LC_12_24_5  (
            .in0(N__16351),
            .in1(N__14348),
            .in2(N__14430),
            .in3(N__16433),
            .lcout(\c0.tx2.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21901),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIGMI01_10_LC_12_24_6 .C_ON=1'b0;
    defparam \c0.d_2_RNIGMI01_10_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIGMI01_10_LC_12_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIGMI01_10_LC_12_24_6  (
            .in0(N__12933),
            .in1(N__14641),
            .in2(_gnd_net_),
            .in3(N__12786),
            .lcout(\c0.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_5_LC_12_24_7 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_5_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_5_LC_12_24_7 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \c0.tx_data_RNO_4_5_LC_12_24_7  (
            .in0(N__19321),
            .in1(N__19169),
            .in2(N__13037),
            .in3(N__12731),
            .lcout(\c0.tx_data_RNO_4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIFMJ01_45_LC_12_25_1 .C_ON=1'b0;
    defparam \c0.d_2_RNIFMJ01_45_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIFMJ01_45_LC_12_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_2_RNIFMJ01_45_LC_12_25_1  (
            .in0(N__12730),
            .in1(N__14939),
            .in2(_gnd_net_),
            .in3(N__14843),
            .lcout(\c0.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__4_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.data_out_0__4_LC_12_25_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__4_LC_12_25_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_0__4_LC_12_25_2  (
            .in0(N__13351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(),
            .sr(N__17341));
    defparam \c0.data_out_2__1_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.data_out_2__1_LC_12_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__1_LC_12_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_2__1_LC_12_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13352),
            .lcout(\c0.d_2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(),
            .sr(N__17341));
    defparam \c0.data_out_3__5_LC_12_25_4 .C_ON=1'b0;
    defparam \c0.data_out_3__5_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__5_LC_12_25_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__5_LC_12_25_4  (
            .in0(N__13353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(),
            .sr(N__17341));
    defparam \c0.data_out_0__1_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.data_out_0__1_LC_12_25_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_0__1_LC_12_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__1_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13350),
            .lcout(\c0.d_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(),
            .sr(N__17341));
    defparam \c0.data_out_3__6_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.data_out_3__6_LC_12_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__6_LC_12_25_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_3__6_LC_12_25_6  (
            .in0(N__13354),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(),
            .sr(N__17341));
    defparam \c0.data_out_7__RNO_1_0_LC_12_25_7 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_0_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_0_LC_12_25_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_0_LC_12_25_7  (
            .in0(N__14899),
            .in1(N__12707),
            .in2(N__14505),
            .in3(N__12944),
            .lcout(\c0.nextCRC16_3_0_a2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_2_RNIK3C71_13_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.d_2_RNIK3C71_13_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIK3C71_13_LC_12_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_2_RNIK3C71_13_LC_12_26_0  (
            .in0(N__13094),
            .in1(N__13004),
            .in2(N__14629),
            .in3(N__13029),
            .lcout(\c0.nextCRC16_3_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__5_LC_12_26_2 .C_ON=1'b0;
    defparam \c0.data_out_1__5_LC_12_26_2 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_1__5_LC_12_26_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_1__5_LC_12_26_2  (
            .in0(N__13356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21916),
            .ce(),
            .sr(N__17340));
    defparam \c0.data_out_7__RNO_1_2_LC_12_26_4 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_2_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_2_LC_12_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_2_LC_12_26_4  (
            .in0(N__13093),
            .in1(N__15360),
            .in2(N__14628),
            .in3(N__13060),
            .lcout(\c0.nextCRC16_3_0_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__0_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.data_out_0__0_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__0_LC_12_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__0_LC_12_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13355),
            .lcout(\c0.d_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21916),
            .ce(),
            .sr(N__17340));
    defparam \c0.d_2_RNIIJMM_15_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.d_2_RNIIJMM_15_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_2_RNIIJMM_15_LC_12_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.d_2_RNIIJMM_15_LC_12_26_6  (
            .in0(_gnd_net_),
            .in1(N__15282),
            .in2(_gnd_net_),
            .in3(N__13059),
            .lcout(\c0.nextCRC16_3_4_0 ),
            .ltout(\c0.nextCRC16_3_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_3_0_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_3_0_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_3_0_LC_12_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_3_0_LC_12_26_7  (
            .in0(N__13030),
            .in1(N__13012),
            .in2(N__12974),
            .in3(N__12960),
            .lcout(\c0.nextCRC16_3_0_a2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__5_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.data_out_6__5_LC_12_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__5_LC_12_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__5_LC_12_27_1  (
            .in0(N__14618),
            .in1(N__12919),
            .in2(_gnd_net_),
            .in3(N__13179),
            .lcout(\c0.data_out_6_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21925),
            .ce(N__17290),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__7_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.data_out_6__7_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__7_LC_12_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_6__7_LC_12_27_4  (
            .in0(N__12872),
            .in1(N__13159),
            .in2(N__12866),
            .in3(N__13143),
            .lcout(\c0.data_out_6_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21925),
            .ce(N__17290),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__0_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.data_out_2__0_LC_12_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_2__0_LC_12_28_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_out_2__0_LC_12_28_0  (
            .in0(N__13358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21930),
            .ce(),
            .sr(N__17337));
    defparam \c0.data_out_3__7_LC_12_28_1 .C_ON=1'b0;
    defparam \c0.data_out_3__7_LC_12_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__7_LC_12_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__7_LC_12_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13359),
            .lcout(\c0.d_2_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21930),
            .ce(),
            .sr(N__17337));
    defparam \c0.data_out_3__0_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.data_out_3__0_LC_12_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__0_LC_12_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_3__0_LC_12_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.d_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21930),
            .ce(),
            .sr(N__17337));
    defparam \c0.data_out_0__5_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.data_out_0__5_LC_12_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__5_LC_12_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_out_0__5_LC_12_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13357),
            .lcout(\c0.d_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21930),
            .ce(),
            .sr(N__17337));
    defparam \c0.data_out_7__1_LC_12_29_2 .C_ON=1'b0;
    defparam \c0.data_out_7__1_LC_12_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__1_LC_12_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__1_LC_12_29_2  (
            .in0(N__13186),
            .in1(N__13163),
            .in2(N__14825),
            .in3(N__13148),
            .lcout(\c0.data_out_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21931),
            .ce(N__17287),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_5_LC_13_17_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_5_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_5_LC_13_17_0 .LUT_INIT=16'b0101110101111111;
    LogicCell40 \c0.tx2_data_RNO_0_5_LC_13_17_0  (
            .in0(N__17856),
            .in1(N__20926),
            .in2(N__13112),
            .in3(N__13510),
            .lcout(\c0.tx2_data_1_0_i_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__5_LC_13_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__5_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__5_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__5_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19967),
            .lcout(\c0.data_in_frame_7_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21857),
            .ce(N__21583),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__5_LC_13_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__5_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__5_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__5_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19985),
            .lcout(\c0.d_4_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21857),
            .ce(N__21583),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_7_LC_13_17_3 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_7_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_7_LC_13_17_3 .LUT_INIT=16'b0011101101111111;
    LogicCell40 \c0.tx2_data_RNO_0_7_LC_13_17_3  (
            .in0(N__20927),
            .in1(N__17857),
            .in2(N__13103),
            .in3(N__15524),
            .lcout(\c0.tx2_data_1_0_i_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__7_LC_13_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__7_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__7_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__7_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22238),
            .lcout(\c0.data_in_frame_7_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21857),
            .ce(N__21583),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__7_LC_13_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__7_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__7_LC_13_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_5__7_LC_13_17_5  (
            .in0(N__20666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21857),
            .ce(N__21583),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_10_LC_13_17_6 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_10_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_10_LC_13_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.wait_for_transmission_RNO_10_LC_13_17_6  (
            .in0(N__17999),
            .in1(N__15390),
            .in2(N__15527),
            .in3(N__15456),
            .lcout(),
            .ltout(\c0.wait_for_transmission_RNOZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_8_LC_13_17_7 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_8_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_8_LC_13_17_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.wait_for_transmission_RNO_8_LC_13_17_7  (
            .in0(N__15557),
            .in1(N__16247),
            .in2(N__13568),
            .in3(N__18590),
            .lcout(\c0.g0_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI5L571_45_LC_13_18_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI5L571_45_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI5L571_45_LC_13_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI5L571_45_LC_13_18_0  (
            .in0(N__13725),
            .in1(N__13544),
            .in2(N__13514),
            .in3(N__15628),
            .lcout(\c0.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI8A8H_26_LC_13_18_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI8A8H_26_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI8A8H_26_LC_13_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI8A8H_26_LC_13_18_1  (
            .in0(N__18429),
            .in1(N__16716),
            .in2(N__13496),
            .in3(N__17188),
            .lcout(),
            .ltout(\c0.un1_data_in_6__7_0_a2_17_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI6CFJ4_26_LC_13_18_2 .C_ON=1'b0;
    defparam \c0.d_4_RNI6CFJ4_26_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI6CFJ4_26_LC_13_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI6CFJ4_26_LC_13_18_2  (
            .in0(N__13782),
            .in1(N__14799),
            .in2(N__13481),
            .in3(N__15808),
            .lcout(\c0.un1_data_in_6__7_0_a2_17_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIU7HB6_19_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIU7HB6_19_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIU7HB6_19_LC_13_18_4 .LUT_INIT=16'b0100000000000100;
    LogicCell40 \c0.d_4_RNIU7HB6_19_LC_13_18_4  (
            .in0(N__18062),
            .in1(N__15680),
            .in2(N__13472),
            .in3(N__15809),
            .lcout(\c0.g0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIIVJN_13_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIIVJN_13_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIIVJN_13_LC_13_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIIVJN_13_LC_13_18_5  (
            .in0(N__15644),
            .in1(N__16715),
            .in2(N__15780),
            .in3(N__17062),
            .lcout(),
            .ltout(\c0.un1_data_in_7__0_0_a2_1_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIG1RP4_13_LC_13_18_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIG1RP4_13_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIG1RP4_13_LC_13_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIG1RP4_13_LC_13_18_6  (
            .in0(N__13781),
            .in1(N__14798),
            .in2(N__13448),
            .in3(N__15807),
            .lcout(\c0.un1_data_in_7__0_0_a2_1_a2_5_0 ),
            .ltout(\c0.un1_data_in_7__0_0_a2_1_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIN2KLB_14_LC_13_18_7 .C_ON=1'b0;
    defparam \c0.d_4_RNIN2KLB_14_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIN2KLB_14_LC_13_18_7 .LUT_INIT=16'b0000001111000000;
    LogicCell40 \c0.d_4_RNIN2KLB_14_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__17705),
            .in2(N__13445),
            .in3(N__17692),
            .lcout(\c0.tx2_transmit_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIN7VG_17_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIN7VG_17_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIN7VG_17_LC_13_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIN7VG_17_LC_13_19_0  (
            .in0(N__13962),
            .in1(N__13731),
            .in2(N__14064),
            .in3(N__15526),
            .lcout(),
            .ltout(\c0.un1_data_in_7__3_0_a2_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIORVS2_43_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIORVS2_43_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIORVS2_43_LC_13_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIORVS2_43_LC_13_19_1  (
            .in0(N__17035),
            .in1(N__15671),
            .in2(N__13787),
            .in3(N__13784),
            .lcout(\c0.un1_data_in_7__3_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__1_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__1_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__1_LC_13_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__1_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13763),
            .lcout(\c0.d_4_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21869),
            .ce(N__21589),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__6_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__6_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__6_LC_13_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__6_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13709),
            .lcout(\c0.d_4_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21869),
            .ce(N__21589),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIA0HJ_0_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIA0HJ_0_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIA0HJ_0_LC_13_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNIA0HJ_0_LC_13_19_4  (
            .in0(N__13961),
            .in1(N__13629),
            .in2(_gnd_net_),
            .in3(N__13609),
            .lcout(\c0.N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__0_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__0_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__0_LC_13_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__0_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13685),
            .lcout(\c0.d_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21869),
            .ce(N__21589),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__0_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__0_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__0_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__0_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13667),
            .lcout(\c0.d_4_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21869),
            .ce(N__21589),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_0_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_0_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_0_LC_13_19_7 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \c0.tx2_data_RNO_3_0_LC_13_19_7  (
            .in0(N__18281),
            .in1(N__19541),
            .in2(N__13613),
            .in3(N__18911),
            .lcout(\c0.tx2_data_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__4_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__4_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__4_LC_13_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__4_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13589),
            .lcout(\c0.d_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__2_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__2_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__2_LC_13_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__2_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13943),
            .lcout(\c0.d_4_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__3_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__3_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__3_LC_13_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__3_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13928),
            .lcout(\c0.d_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__5_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__5_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__5_LC_13_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__5_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13898),
            .lcout(\c0.d_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__5_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__5_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__5_LC_13_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__5_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13871),
            .lcout(\c0.d_4_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__1_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__1_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__1_LC_13_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__1_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13846),
            .lcout(\c0.d_4_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__1_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__1_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__1_LC_13_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__1_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13823),
            .lcout(\c0.d_4_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__3_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__3_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__3_LC_13_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__3_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13808),
            .lcout(\c0.d_4_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__21592),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_6_LC_13_21_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_6_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_6_LC_13_21_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \c0.tx2_data_RNO_3_6_LC_13_21_1  (
            .in0(N__20928),
            .in1(N__18092),
            .in2(_gnd_net_),
            .in3(N__15461),
            .lcout(),
            .ltout(\c0.tx2_data_1_iv_3_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_6_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_6_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_6_LC_13_21_2 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \c0.tx2_data_RNO_1_6_LC_13_21_2  (
            .in0(N__20410),
            .in1(_gnd_net_),
            .in2(N__13790),
            .in3(N__20340),
            .lcout(\c0.tx2_data_1_iv_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI1VL6_13_LC_13_21_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI1VL6_13_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI1VL6_13_LC_13_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI1VL6_13_LC_13_21_3  (
            .in0(N__17055),
            .in1(N__15760),
            .in2(_gnd_net_),
            .in3(N__16691),
            .lcout(\c0.N_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIH9JJ_4_LC_13_21_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIH9JJ_4_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIH9JJ_4_LC_13_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNIH9JJ_4_LC_13_21_4  (
            .in0(N__14150),
            .in1(N__16049),
            .in2(_gnd_net_),
            .in3(N__19687),
            .lcout(\c0.N_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNII9QU3_14_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.d_4_RNII9QU3_14_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNII9QU3_14_LC_13_21_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.d_4_RNII9QU3_14_LC_13_21_5  (
            .in0(N__14022),
            .in1(N__15551),
            .in2(_gnd_net_),
            .in3(N__16099),
            .lcout(\c0.d_4_RNII9QU3Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI675O1_33_LC_13_21_6 .C_ON=1'b0;
    defparam \c0.d_4_RNI675O1_33_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI675O1_33_LC_13_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI675O1_33_LC_13_21_6  (
            .in0(N__14151),
            .in1(N__15497),
            .in2(N__16277),
            .in3(N__16050),
            .lcout(\c0.un1_data_in_7__7_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_3_LC_13_21_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_3_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_3_LC_13_21_7 .LUT_INIT=16'b0011010111111111;
    LogicCell40 \c0.tx2_data_RNO_0_3_LC_13_21_7  (
            .in0(N__18005),
            .in1(N__20612),
            .in2(N__20940),
            .in3(N__20409),
            .lcout(\c0.tx2_data_1_0_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_5_3_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_5_3_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_5_3_LC_13_22_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \c0.tx2_data_RNO_5_3_LC_13_22_1  (
            .in0(N__20932),
            .in1(N__14030),
            .in2(_gnd_net_),
            .in3(N__15660),
            .lcout(\c0.tx2_data_1_iv_4_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__4_LC_13_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__4_LC_13_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__4_LC_13_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__4_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14093),
            .lcout(\c0.d_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21892),
            .ce(N__21597),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__3_LC_13_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__3_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__3_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__3_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14066),
            .lcout(\c0.data_in_frame_7_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21892),
            .ce(N__21597),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_6_LC_13_22_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_6_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_6_LC_13_22_5 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \c0.tx2_data_RNO_4_6_LC_13_22_5  (
            .in0(N__20933),
            .in1(N__14023),
            .in2(N__17869),
            .in3(N__13970),
            .lcout(),
            .ltout(\c0.tx2_data_1_iv_4_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_6_LC_13_22_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_6_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_6_LC_13_22_6 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \c0.tx2_data_RNO_2_6_LC_13_22_6  (
            .in0(N__18449),
            .in1(N__17865),
            .in2(N__14456),
            .in3(N__20341),
            .lcout(\c0.tx2_data_1_iv_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__3_LC_13_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__3_LC_13_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__3_LC_13_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__3_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14453),
            .lcout(\c0.d_4_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21892),
            .ce(N__21597),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_a2_0_LC_13_23_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_a2_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_a2_0_LC_13_23_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx2.r_SM_Main_7_1_0__m5_0_a2_0_LC_13_23_0  (
            .in0(N__19763),
            .in1(N__16346),
            .in2(N__14421),
            .in3(N__14341),
            .lcout(\c0.tx2.r_Tx_Data_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_0_LC_13_23_1 .LUT_INIT=16'b1110000011000010;
    LogicCell40 \c0.tx2.r_Bit_Index_0_LC_13_23_1  (
            .in0(N__16347),
            .in1(N__16381),
            .in2(N__16463),
            .in3(N__16438),
            .lcout(\c0.tx2.r_Bit_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_RNIMCBI_0_LC_13_23_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_RNIMCBI_0_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_RNIMCBI_0_LC_13_23_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx2.r_SM_Main_RNIMCBI_0_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__14398),
            .in2(_gnd_net_),
            .in3(N__14340),
            .lcout(\c0.tx2.N_257 ),
            .ltout(\c0.tx2.N_257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_o2_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_o2_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_7_1_0__m5_0_o2_LC_13_23_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.tx2.r_SM_Main_7_1_0__m5_0_o2_LC_13_23_3  (
            .in0(N__16457),
            .in1(N__16302),
            .in2(N__14303),
            .in3(N__16437),
            .lcout(\c0.tx2.N_261 ),
            .ltout(\c0.tx2.N_261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_2_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_2_LC_13_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_2_LC_13_23_4 .LUT_INIT=16'b0011000000000011;
    LogicCell40 \c0.tx2.r_Bit_Index_2_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__14294),
            .in2(N__14237),
            .in3(N__14232),
            .lcout(\c0.tx2.r_Bit_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_LC_13_23_5 .C_ON=1'b0;
    defparam \c0.tx_transmit_LC_13_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_LC_13_23_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.tx_transmit_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__14200),
            .in2(_gnd_net_),
            .in3(N__14186),
            .lcout(\c0.tx_transmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21902),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_RNI6GJO_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.tx_active_RNI6GJO_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx_active_RNI6GJO_LC_13_23_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.tx_active_RNI6GJO_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__14199),
            .in2(_gnd_net_),
            .in3(N__14185),
            .lcout(\c0.byte_transmit_counter15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_6_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_6_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_6_LC_13_24_0 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \c0.tx2.r_Tx_Data_6_LC_13_24_0  (
            .in0(N__20600),
            .in1(N__14765),
            .in2(N__14756),
            .in3(N__20355),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21909),
            .ce(N__20750),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_3_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_3_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_3_LC_13_24_1 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \c0.tx_data_RNO_1_3_LC_13_24_1  (
            .in0(N__19312),
            .in1(N__14465),
            .in2(N__14735),
            .in3(N__19172),
            .lcout(\c0.tx_data_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_1_7_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_1_7_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_1_7_LC_13_24_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \c0.tx_data_RNO_1_7_LC_13_24_3  (
            .in0(N__19313),
            .in1(N__19173),
            .in2(N__14693),
            .in3(N__15365),
            .lcout(\c0.tx_data_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_2_LC_13_24_4 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_2_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_2_LC_13_24_4 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx_data_RNO_3_2_LC_13_24_4  (
            .in0(N__19170),
            .in1(N__17434),
            .in2(N__15257),
            .in3(N__19314),
            .lcout(),
            .ltout(\c0.tx_data_RNO_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_2_2_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_2_2_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_2_2_LC_13_24_5 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \c0.tx_data_RNO_2_2_LC_13_24_5  (
            .in0(N__17520),
            .in1(N__16782),
            .in2(N__14669),
            .in3(N__14582),
            .lcout(\c0.tx_data_1_0_i_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_4_2_LC_13_24_6 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_4_2_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_4_2_LC_13_24_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx_data_RNO_4_2_LC_13_24_6  (
            .in0(N__19171),
            .in1(N__14653),
            .in2(N__14630),
            .in3(N__19311),
            .lcout(\c0.tx_data_RNO_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNIRD6P_0_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNIRD6P_0_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNIRD6P_0_LC_13_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter_RNIRD6P_0_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__16781),
            .in2(_gnd_net_),
            .in3(N__17475),
            .lcout(\c0.N_201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__6_LC_13_25_1 .C_ON=1'b0;
    defparam \c0.data_out_6__6_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__6_LC_13_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_6__6_LC_13_25_1  (
            .in0(N__15331),
            .in1(N__14974),
            .in2(_gnd_net_),
            .in3(N__14576),
            .lcout(\c0.data_out_6_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21917),
            .ce(N__17292),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__3_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.data_out_7__3_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__3_LC_13_25_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__3_LC_13_25_2  (
            .in0(N__14546),
            .in1(N__14500),
            .in2(N__14912),
            .in3(N__15176),
            .lcout(\c0.data_out_7_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21917),
            .ce(N__17292),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_1_3_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_3_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_3_LC_13_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_3_LC_13_26_2  (
            .in0(N__15142),
            .in1(N__15361),
            .in2(N__15330),
            .in3(N__15287),
            .lcout(),
            .ltout(\c0.un105_newcrc_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_3_LC_13_26_3 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_3_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_3_LC_13_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_0_3_LC_13_26_3  (
            .in0(N__15239),
            .in1(N__15209),
            .in2(N__15179),
            .in3(N__14940),
            .lcout(\c0.un105_newcrc_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_1_6_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_1_6_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_1_6_LC_13_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_1_6_LC_13_27_2  (
            .in0(N__15159),
            .in1(N__15143),
            .in2(N__15110),
            .in3(N__14856),
            .lcout(\c0.un144_newcrc_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_6_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_6_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_6_LC_13_27_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_7__RNO_0_6_LC_13_27_5  (
            .in0(N__15061),
            .in1(N__15022),
            .in2(_gnd_net_),
            .in3(N__16515),
            .lcout(\c0.un144_newcrc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_1_LC_13_29_7 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_1_LC_13_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_1_LC_13_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_7__RNO_0_1_LC_13_29_7  (
            .in0(N__14978),
            .in1(N__14960),
            .in2(N__14920),
            .in3(N__14861),
            .lcout(\c0.nextCRC16_3_0_a2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI22UN_24_LC_14_17_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI22UN_24_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI22UN_24_LC_14_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI22UN_24_LC_14_17_0  (
            .in0(N__18649),
            .in1(N__20534),
            .in2(N__14816),
            .in3(N__16132),
            .lcout(\c0.un1_data_in_6__4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__RNIFRNC_4_LC_14_17_1 .C_ON=1'b0;
    defparam \c0.data_in_6__RNIFRNC_4_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_6__RNIFRNC_4_LC_14_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_6__RNIFRNC_4_LC_14_17_1  (
            .in0(N__16619),
            .in1(N__15781),
            .in2(N__22271),
            .in3(N__16708),
            .lcout(\c0.un1_data_in_6__4_0_a2_5_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI9IAQ1_31_LC_14_17_2 .C_ON=1'b0;
    defparam \c0.d_4_RNI9IAQ1_31_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI9IAQ1_31_LC_14_17_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.d_4_RNI9IAQ1_31_LC_14_17_2  (
            .in0(N__18347),
            .in1(N__14807),
            .in2(N__14780),
            .in3(N__17917),
            .lcout(),
            .ltout(\c0.wait_for_transmission4_12_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI7HDA4_24_LC_14_17_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI7HDA4_24_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI7HDA4_24_LC_14_17_3 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \c0.d_4_RNI7HDA4_24_LC_14_17_3  (
            .in0(N__15563),
            .in1(N__15638),
            .in2(N__15632),
            .in3(N__15629),
            .lcout(\c0.wait_for_transmission4_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__RNIBJH41_6_LC_14_17_4 .C_ON=1'b0;
    defparam \c0.data_in_7__RNIBJH41_6_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_7__RNIBJH41_6_LC_14_17_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_in_7__RNIBJH41_6_LC_14_17_4  (
            .in0(N__16151),
            .in1(N__17995),
            .in2(N__19877),
            .in3(N__15605),
            .lcout(\c0.un1_data_in_7__6_0_a2_5_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_11_LC_14_17_5 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_11_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_11_LC_14_17_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.wait_for_transmission_RNO_11_LC_14_17_5  (
            .in0(N__16620),
            .in1(N__16030),
            .in2(_gnd_net_),
            .in3(N__18253),
            .lcout(\c0.wait_for_transmission_RNOZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI4SA91_10_LC_14_18_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI4SA91_10_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI4SA91_10_LC_14_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI4SA91_10_LC_14_18_0  (
            .in0(N__16029),
            .in1(N__18252),
            .in2(N__16627),
            .in3(N__15490),
            .lcout(\c0.un1_data_in_6__7_0_a2_17_a2_4_1 ),
            .ltout(\c0.un1_data_in_6__7_0_a2_17_a2_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIV4MJ3_24_LC_14_18_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIV4MJ3_24_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIV4MJ3_24_LC_14_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIV4MJ3_24_LC_14_18_1  (
            .in0(N__16150),
            .in1(N__18572),
            .in2(N__15530),
            .in3(N__15862),
            .lcout(\c0.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIJLQL_47_LC_14_18_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIJLQL_47_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIJLQL_47_LC_14_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIJLQL_47_LC_14_18_2  (
            .in0(N__17991),
            .in1(N__15383),
            .in2(N__15525),
            .in3(N__15452),
            .lcout(\c0.N_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__6_LC_14_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__6_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__6_LC_14_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__6_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15479),
            .lcout(\c0.d_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21870),
            .ce(N__21584),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__3_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__3_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__3_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__3_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15431),
            .lcout(\c0.d_4_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21870),
            .ce(N__21584),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIQCTH_24_LC_14_18_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIQCTH_24_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIQCTH_24_LC_14_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIQCTH_24_LC_14_18_6  (
            .in0(N__20533),
            .in1(N__18178),
            .in2(N__18650),
            .in3(N__16124),
            .lcout(\c0.un1_data_in_6__7_0_a2_17_a2_4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__3_LC_14_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__3_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__3_LC_14_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__3_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15851),
            .lcout(\c0.d_4_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21870),
            .ce(N__21584),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIO7RC_28_LC_14_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIO7RC_28_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIO7RC_28_LC_14_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIO7RC_28_LC_14_19_0  (
            .in0(N__20588),
            .in1(N__18967),
            .in2(N__15898),
            .in3(N__15670),
            .lcout(),
            .ltout(\c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI15AH_12_LC_14_19_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI15AH_12_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI15AH_12_LC_14_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.d_4_RNI15AH_12_LC_14_19_1  (
            .in0(N__17180),
            .in1(_gnd_net_),
            .in2(N__15833),
            .in3(N__18431),
            .lcout(\c0.un1_data_in_6__6_0_a2_0_a2_3 ),
            .ltout(\c0.un1_data_in_6__6_0_a2_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNITU3G2_19_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.d_4_RNITU3G2_19_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNITU3G2_19_LC_14_19_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \c0.d_4_RNITU3G2_19_LC_14_19_2  (
            .in0(N__15830),
            .in1(N__15732),
            .in2(N__15821),
            .in3(N__15810),
            .lcout(\c0.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIN4PC_27_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIN4PC_27_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIN4PC_27_LC_14_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIN4PC_27_LC_14_19_3  (
            .in0(N__16018),
            .in1(N__15761),
            .in2(N__19928),
            .in3(N__17800),
            .lcout(),
            .ltout(\c0.un1_data_in_6__5_0_a2_5_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI23VN_12_LC_14_19_4 .C_ON=1'b0;
    defparam \c0.d_4_RNI23VN_12_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI23VN_12_LC_14_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI23VN_12_LC_14_19_4  (
            .in0(N__18430),
            .in1(N__17179),
            .in2(N__15737),
            .in3(N__16125),
            .lcout(\c0.un1_data_in_6__5 ),
            .ltout(\c0.un1_data_in_6__5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIOEM13_24_LC_14_19_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIOEM13_24_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIOEM13_24_LC_14_19_5 .LUT_INIT=16'b0000000000001001;
    LogicCell40 \c0.d_4_RNIOEM13_24_LC_14_19_5  (
            .in0(N__15733),
            .in1(N__15694),
            .in2(N__15683),
            .in3(N__18188),
            .lcout(\c0.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIH0UG_27_LC_14_19_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIH0UG_27_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIH0UG_27_LC_14_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIH0UG_27_LC_14_19_6  (
            .in0(N__17799),
            .in1(N__15669),
            .in2(N__18746),
            .in3(N__17178),
            .lcout(\c0.un1_data_in_7__0_0_a2_1_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI21N6_11_LC_14_19_7 .C_ON=1'b0;
    defparam \c0.d_4_RNI21N6_11_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI21N6_11_LC_14_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI21N6_11_LC_14_19_7  (
            .in0(N__15890),
            .in1(N__18209),
            .in2(_gnd_net_),
            .in3(N__17770),
            .lcout(\c0.d_4_RNI21N6Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIQ7PC_23_LC_14_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIQ7PC_23_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIQ7PC_23_LC_14_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIQ7PC_23_LC_14_20_0  (
            .in0(N__18036),
            .in1(N__20532),
            .in2(N__20641),
            .in3(N__20158),
            .lcout(),
            .ltout(\c0.un1_data_in_6__3_0_a2_5_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIRKQ41_10_LC_14_20_1 .C_ON=1'b0;
    defparam \c0.d_4_RNIRKQ41_10_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIRKQ41_10_LC_14_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.d_4_RNIRKQ41_10_LC_14_20_1  (
            .in0(N__15983),
            .in1(N__16615),
            .in2(N__16034),
            .in3(N__16025),
            .lcout(\c0.un1_data_in_6__3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIPIKJ_39_LC_14_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIPIKJ_39_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIPIKJ_39_LC_14_20_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.d_4_RNIPIKJ_39_LC_14_20_2  (
            .in0(N__18248),
            .in1(N__15891),
            .in2(_gnd_net_),
            .in3(N__18211),
            .lcout(\c0.un1_data_in_6__3_0_a2_5_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__1_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__1_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__1_LC_14_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__1_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15977),
            .lcout(\c0.d_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__21590),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__7_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__7_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__7_LC_14_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__7_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15947),
            .lcout(\c0.d_4_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__21590),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__7_LC_14_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__7_LC_14_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__7_LC_14_20_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_4__7_LC_14_20_5  (
            .in0(N__18841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__21590),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__0_LC_14_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__0_LC_14_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__0_LC_14_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__0_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15917),
            .lcout(\c0.d_4_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__21590),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__5_LC_14_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__5_LC_14_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__5_LC_14_20_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_in_frame_4__5_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__20002),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21884),
            .ce(N__21590),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI6FQT_21_LC_14_21_0 .C_ON=1'b0;
    defparam \c0.d_4_RNI6FQT_21_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI6FQT_21_LC_14_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNI6FQT_21_LC_14_21_0  (
            .in0(N__20470),
            .in1(N__20430),
            .in2(N__22227),
            .in3(N__18492),
            .lcout(\c0.un1_data_in_7__7_0_a2_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__5_LC_14_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__5_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__5_LC_14_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__5_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16268),
            .lcout(\c0.d_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21893),
            .ce(N__21593),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_9_LC_14_21_2 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_9_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_9_LC_14_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.wait_for_transmission_RNO_9_LC_14_21_2  (
            .in0(N__19713),
            .in1(N__20469),
            .in2(N__18371),
            .in3(N__16167),
            .lcout(\c0.wait_for_transmission_RNOZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__2_LC_14_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__2_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__2_LC_14_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__2_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16235),
            .lcout(\c0.d_4_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21893),
            .ce(N__21593),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__4_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__4_LC_14_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__4_LC_14_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__4_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16208),
            .lcout(\c0.d_4_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21893),
            .ce(N__21593),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_5__6_LC_14_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_5__6_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_5__6_LC_14_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_5__6_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19895),
            .lcout(\c0.d_4_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21893),
            .ce(N__21593),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIABPL_18_LC_14_21_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIABPL_18_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIABPL_18_LC_14_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIABPL_18_LC_14_21_6  (
            .in0(N__19712),
            .in1(N__20468),
            .in2(N__18370),
            .in3(N__16166),
            .lcout(\c0.N_124 ),
            .ltout(\c0.N_124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIPF9J2_37_LC_14_21_7 .C_ON=1'b0;
    defparam \c0.d_4_RNIPF9J2_37_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIPF9J2_37_LC_14_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIPF9J2_37_LC_14_21_7  (
            .in0(N__18680),
            .in1(N__18582),
            .in2(N__16136),
            .in3(N__16133),
            .lcout(\c0.d_4_RNIPF9J2Z0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__1_LC_14_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__1_LC_14_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__1_LC_14_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__1_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16085),
            .lcout(\c0.d_4_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21903),
            .ce(N__21596),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__0_LC_14_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__0_LC_14_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__0_LC_14_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__0_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18765),
            .lcout(\c0.data_in_frame_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21903),
            .ce(N__21596),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__2_LC_14_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__2_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__2_LC_14_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_3__2_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16745),
            .lcout(\c0.d_4_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21903),
            .ce(N__21596),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__1_LC_14_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__1_LC_14_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__1_LC_14_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__1_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18801),
            .lcout(\c0.data_in_frame_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21903),
            .ce(N__21596),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__2_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__2_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__2_LC_14_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__2_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16655),
            .lcout(\c0.d_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21903),
            .ce(N__21596),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__0_LC_14_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__0_LC_14_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__0_LC_14_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__0_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18738),
            .lcout(\c0.data_in_frame_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21903),
            .ce(N__21596),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__RNO_0_7_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.data_out_7__RNO_0_7_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_7__RNO_0_7_LC_14_23_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.data_out_7__RNO_0_7_LC_14_23_1  (
            .in0(N__16567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16523),
            .lcout(\c0.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_6_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_6_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_6_LC_14_23_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_6_LC_14_23_4  (
            .in0(N__21413),
            .in1(N__21497),
            .in2(_gnd_net_),
            .in3(N__21324),
            .lcout(\c0.rx.r_Rx_Bytece_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_RNO_0_1_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_RNO_0_1_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_RNO_0_1_LC_14_23_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.tx2.r_Bit_Index_RNO_0_1_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__16462),
            .in2(_gnd_net_),
            .in3(N__16439),
            .lcout(),
            .ltout(\c0.tx2.N_258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_1_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_1_LC_14_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_1_LC_14_23_7 .LUT_INIT=16'b1100100110001000;
    LogicCell40 \c0.tx2.r_Bit_Index_1_LC_14_23_7  (
            .in0(N__16382),
            .in1(N__16303),
            .in2(N__16370),
            .in3(N__16367),
            .lcout(\c0.tx2.r_Bit_IndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21910),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_3_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_3_LC_14_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_3_LC_14_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_3_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21918),
            .ce(N__19030),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_6_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_6_LC_14_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_6_LC_14_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_6_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21918),
            .ce(N__19030),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_3_6_LC_14_24_2 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_3_6_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_3_6_LC_14_24_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx_data_RNO_3_6_LC_14_24_2  (
            .in0(N__19077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19287),
            .lcout(),
            .ltout(\c0.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_data_RNO_0_6_LC_14_24_3 .C_ON=1'b0;
    defparam \c0.tx_data_RNO_0_6_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx_data_RNO_0_6_LC_14_24_3 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \c0.tx_data_RNO_0_6_LC_14_24_3  (
            .in0(N__16967),
            .in1(N__17357),
            .in2(N__16961),
            .in3(N__17503),
            .lcout(\c0.N_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNIA0ET3_2_LC_14_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNIA0ET3_2_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNIA0ET3_2_LC_14_24_4 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \c0.byte_transmit_counter_RNIA0ET3_2_LC_14_24_4  (
            .in0(N__19019),
            .in1(N__19423),
            .in2(N__19114),
            .in3(N__19286),
            .lcout(\c0.data_out_0__1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNI3M6P_3_LC_14_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNI3M6P_3_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNI3M6P_3_LC_14_24_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.byte_transmit_counter_RNI3M6P_3_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__16931),
            .in2(_gnd_net_),
            .in3(N__16925),
            .lcout(),
            .ltout(\c0.m2_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNIQP0V1_4_LC_14_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNIQP0V1_4_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNIQP0V1_4_LC_14_24_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.byte_transmit_counter_RNIQP0V1_4_LC_14_24_6  (
            .in0(N__19040),
            .in1(N__18695),
            .in2(N__16919),
            .in3(N__17573),
            .lcout(\c0.N_129_mux ),
            .ltout(\c0.N_129_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_RNI92KB2_2_LC_14_24_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_RNI92KB2_2_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_RNI92KB2_2_LC_14_24_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.byte_transmit_counter_RNI92KB2_2_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16916),
            .in3(N__19076),
            .lcout(\c0.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1_LC_14_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1_LC_14_25_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \c0.byte_transmit_counter_1_LC_14_25_0  (
            .in0(N__16807),
            .in1(N__17505),
            .in2(_gnd_net_),
            .in3(N__19319),
            .lcout(\c0.byte_transmit_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21926),
            .ce(N__19034),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4_LC_14_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_4_LC_14_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_4_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21926),
            .ce(N__19034),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0_LC_14_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0_LC_14_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_0_LC_14_25_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.byte_transmit_counter_0_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__17504),
            .in2(_gnd_net_),
            .in3(N__19318),
            .lcout(\c0.byte_transmit_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21926),
            .ce(N__19034),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__6_LC_14_27_1 .C_ON=1'b0;
    defparam \c0.data_out_7__6_LC_14_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__6_LC_14_27_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_7__6_LC_14_27_1  (
            .in0(N__17441),
            .in1(N__17433),
            .in2(N__17402),
            .in3(N__17393),
            .lcout(\c0.data_out_7_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21932),
            .ce(N__17288),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_4_LC_15_16_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_4_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_4_LC_15_16_0 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \c0.tx2_data_RNO_1_4_LC_15_16_0  (
            .in0(N__20327),
            .in1(N__17192),
            .in2(N__17858),
            .in3(N__17138),
            .lcout(\c0.tx2_data_1_0_i_1_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_7_LC_15_17_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_7_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_7_LC_15_17_0 .LUT_INIT=16'b0111111101110111;
    LogicCell40 \c0.tx2.r_Tx_Data_7_LC_15_17_0  (
            .in0(N__17102),
            .in1(N__17876),
            .in2(N__17093),
            .in3(N__20277),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21871),
            .ce(N__20734),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_5_LC_15_17_1 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_5_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_5_LC_15_17_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \c0.tx2_data_RNO_3_5_LC_15_17_1  (
            .in0(N__20845),
            .in1(N__17835),
            .in2(N__20326),
            .in3(N__17066),
            .lcout(),
            .ltout(\c0.data_in_frame_1__m_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_5_LC_15_17_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_5_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_5_LC_15_17_2 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \c0.tx2_data_RNO_1_5_LC_15_17_2  (
            .in0(N__17042),
            .in1(N__20275),
            .in2(N__16997),
            .in3(N__18985),
            .lcout(),
            .ltout(\c0.tx2_data_1_iv_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_5_LC_15_17_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_5_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_5_LC_15_17_3 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \c0.tx2.r_Tx_Data_5_LC_15_17_3  (
            .in0(N__20276),
            .in1(N__16994),
            .in2(N__16985),
            .in3(N__20189),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21871),
            .ce(N__20734),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_7_LC_15_17_4 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_7_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_7_LC_15_17_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \c0.tx2_data_RNO_3_7_LC_15_17_4  (
            .in0(N__17945),
            .in1(N__20270),
            .in2(N__17850),
            .in3(N__20844),
            .lcout(),
            .ltout(\c0.data_in_frame_1__m_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_1_7_LC_15_17_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_1_7_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_1_7_LC_15_17_5 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \c0.tx2_data_RNO_1_7_LC_15_17_5  (
            .in0(N__20274),
            .in1(N__18986),
            .in2(N__17921),
            .in3(N__17918),
            .lcout(\c0.tx2_data_1_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIJBBP_6_LC_15_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIJBBP_6_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIJBBP_6_LC_15_17_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \c0.byte_transmit_counter2_RNIJBBP_6_LC_15_17_6  (
            .in0(N__19480),
            .in1(N__19607),
            .in2(N__19648),
            .in3(N__19738),
            .lcout(\c0.N_205 ),
            .ltout(\c0.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_3_LC_15_17_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_3_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_3_LC_15_17_7 .LUT_INIT=16'b0010111101111111;
    LogicCell40 \c0.tx2_data_RNO_4_3_LC_15_17_7  (
            .in0(N__20846),
            .in1(N__17807),
            .in2(N__17780),
            .in3(N__17777),
            .lcout(\c0.tx2_data_1_iv_4_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI25GA4_LC_15_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI25GA4_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNI25GA4_LC_15_18_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNI25GA4_LC_15_18_0  (
            .in0(N__18011),
            .in1(N__18139),
            .in2(N__17743),
            .in3(N__17726),
            .lcout(),
            .ltout(\c0.g1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i12_7_c_RNIP740G_LC_15_18_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNIP740G_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.FRAME_MATCHER_i12_7_c_RNIP740G_LC_15_18_1 .LUT_INIT=16'b0010000001000000;
    LogicCell40 \c0.FRAME_MATCHER_i12_7_c_RNIP740G_LC_15_18_1  (
            .in0(N__17704),
            .in1(N__17693),
            .in2(N__17663),
            .in3(N__17653),
            .lcout(),
            .ltout(\c0.i12_7_c_RNIP740G_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIM68GI_19_LC_15_18_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIM68GI_19_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIM68GI_19_LC_15_18_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.d_4_RNIM68GI_19_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17636),
            .in3(N__17633),
            .lcout(),
            .ltout(\c0.g1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI9LFUV_43_LC_15_18_3 .C_ON=1'b0;
    defparam \c0.d_4_RNI9LFUV_43_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI9LFUV_43_LC_15_18_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \c0.d_4_RNI9LFUV_43_LC_15_18_3  (
            .in0(N__17620),
            .in1(N__17609),
            .in2(N__17591),
            .in3(N__17588),
            .lcout(\c0.d_4_RNI9LFUVZ0Z_43 ),
            .ltout(\c0.d_4_RNI9LFUVZ0Z_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNI9PP5B1_LC_15_18_4 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNI9PP5B1_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNI9PP5B1_LC_15_18_4 .LUT_INIT=16'b0000010010101011;
    LogicCell40 \c0.wait_for_transmission_RNI9PP5B1_LC_15_18_4  (
            .in0(N__19803),
            .in1(N__19849),
            .in2(N__18068),
            .in3(N__19825),
            .lcout(\c0.wait_for_transmission_RNI9PP5BZ0Z1 ),
            .ltout(\c0.wait_for_transmission_RNI9PP5BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0_LC_15_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_0_LC_15_18_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.byte_transmit_counter2_0_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18065),
            .in3(N__19486),
            .lcout(\c0.byte_transmit_counter2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21877),
            .ce(),
            .sr(N__20053));
    defparam \c0.byte_transmit_counter2_1_LC_15_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_1_LC_15_18_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \c0.byte_transmit_counter2_1_LC_15_18_6  (
            .in0(N__19485),
            .in1(N__20859),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\c0.byte_transmit_counter2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21877),
            .ce(),
            .sr(N__20053));
    defparam \c0.byte_transmit_counter2_2_LC_15_18_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2_LC_15_18_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \c0.byte_transmit_counter2_2_LC_15_18_7  (
            .in0(N__20860),
            .in1(N__20289),
            .in2(N__20087),
            .in3(N__19487),
            .lcout(\c0.byte_transmit_counter2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21877),
            .ce(),
            .sr(N__20053));
    defparam \c0.d_4_RNIBUMH1_0_37_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIBUMH1_0_37_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIBUMH1_0_37_LC_15_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIBUMH1_0_37_LC_15_19_0  (
            .in0(N__18550),
            .in1(N__20159),
            .in2(N__18500),
            .in3(N__18050),
            .lcout(\c0.un1_data_in_6__1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNINGK21_0_21_LC_15_19_1 .C_ON=1'b0;
    defparam \c0.d_4_RNINGK21_0_21_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNINGK21_0_21_LC_15_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNINGK21_0_21_LC_15_19_1  (
            .in0(N__18322),
            .in1(N__18035),
            .in2(N__18280),
            .in3(N__20443),
            .lcout(\c0.g0_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNINGK21_21_LC_15_19_2 .C_ON=1'b0;
    defparam \c0.d_4_RNINGK21_21_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNINGK21_21_LC_15_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNINGK21_21_LC_15_19_2  (
            .in0(N__20442),
            .in1(N__18272),
            .in2(N__18040),
            .in3(N__18321),
            .lcout(\c0.N_126 ),
            .ltout(\c0.N_126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIBUMH1_37_LC_15_19_3 .C_ON=1'b0;
    defparam \c0.d_4_RNIBUMH1_37_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIBUMH1_37_LC_15_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIBUMH1_37_LC_15_19_3  (
            .in0(N__20160),
            .in1(N__18496),
            .in2(N__18014),
            .in3(N__18549),
            .lcout(\c0.un1_data_in_6__1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__RNI15IA_1_LC_15_19_4 .C_ON=1'b0;
    defparam \c0.data_in_6__RNI15IA_1_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_6__RNI15IA_1_LC_15_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_in_6__RNI15IA_1_LC_15_19_4  (
            .in0(N__18003),
            .in1(N__20528),
            .in2(_gnd_net_),
            .in3(N__18805),
            .lcout(\c0.un1_data_in_6__1_0_a2_4_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__7_LC_15_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__7_LC_15_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__7_LC_15_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_0__7_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17960),
            .lcout(\c0.d_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21885),
            .ce(N__21585),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_1__0_LC_15_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_1__0_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_1__0_LC_15_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_1__0_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18308),
            .lcout(\c0.d_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21885),
            .ce(N__21585),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNISRG61_39_LC_15_19_7 .C_ON=1'b0;
    defparam \c0.d_4_RNISRG61_39_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNISRG61_39_LC_15_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNISRG61_39_LC_15_19_7  (
            .in0(N__18273),
            .in1(N__18241),
            .in2(N__22110),
            .in3(N__18210),
            .lcout(\c0.un1_data_in_6__2_0_a2_6_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIK7NH1_0_24_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.d_4_RNIK7NH1_0_24_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIK7NH1_0_24_LC_15_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIK7NH1_0_24_LC_15_20_0  (
            .in0(N__18155),
            .in1(N__20506),
            .in2(N__18644),
            .in3(N__18177),
            .lcout(\c0.un1_data_in_6__2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI76N6_22_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.d_4_RNI76N6_22_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI76N6_22_LC_15_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI76N6_22_LC_15_20_1  (
            .in0(N__20156),
            .in1(N__18482),
            .in2(_gnd_net_),
            .in3(N__18083),
            .lcout(\c0.N_107 ),
            .ltout(\c0.N_107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIK7NH1_24_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.d_4_RNIK7NH1_24_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIK7NH1_24_LC_15_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIK7NH1_24_LC_15_20_2  (
            .in0(N__18154),
            .in1(N__18627),
            .in2(N__18146),
            .in3(N__20507),
            .lcout(\c0.un1_data_in_6__2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_2__6_LC_15_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_2__6_LC_15_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_2__6_LC_15_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_2__6_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18122),
            .lcout(\c0.d_4_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21894),
            .ce(N__21587),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIU6U8_22_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.d_4_RNIU6U8_22_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIU6U8_22_LC_15_20_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.d_4_RNIU6U8_22_LC_15_20_4  (
            .in0(N__18084),
            .in1(N__18626),
            .in2(N__18495),
            .in3(N__20504),
            .lcout(\c0.d_4_RNIU6U8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIU6U8_0_22_LC_15_20_5 .C_ON=1'b0;
    defparam \c0.d_4_RNIU6U8_0_22_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIU6U8_0_22_LC_15_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.d_4_RNIU6U8_0_22_LC_15_20_5  (
            .in0(N__20505),
            .in1(N__18486),
            .in2(N__18640),
            .in3(N__18085),
            .lcout(),
            .ltout(\c0.d_4_RNIU6U8_0Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNIMI4K_37_LC_15_20_6 .C_ON=1'b0;
    defparam \c0.d_4_RNIMI4K_37_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNIMI4K_37_LC_15_20_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.d_4_RNIMI4K_37_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__18689),
            .in2(N__18683),
            .in3(N__20157),
            .lcout(\c0.d_4_RNIMI4KZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_3__0_LC_15_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_3__0_LC_15_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_3__0_LC_15_20_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_3__0_LC_15_20_7  (
            .in0(N__18673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21894),
            .ce(N__21587),
            .sr(_gnd_net_));
    defparam \c0.wait_for_transmission_RNO_7_LC_15_21_0 .C_ON=1'b0;
    defparam \c0.wait_for_transmission_RNO_7_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.wait_for_transmission_RNO_7_LC_15_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.wait_for_transmission_RNO_7_LC_15_21_0  (
            .in0(N__20161),
            .in1(N__18493),
            .in2(N__18589),
            .in3(N__18554),
            .lcout(\c0.un1_data_in_6__1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__4_LC_15_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__4_LC_15_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__4_LC_15_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_4__4_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18521),
            .lcout(\c0.d_4_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21904),
            .ce(N__21591),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_4_LC_15_21_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_4_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_4_LC_15_21_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \c0.tx2_data_RNO_4_4_LC_15_21_2  (
            .in0(N__18455),
            .in1(N__18494),
            .in2(_gnd_net_),
            .in3(N__20919),
            .lcout(\c0.tx2_data_1_iv_5_1_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__4_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__4_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__4_LC_15_21_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_in_frame_6__4_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__22263),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_frame_6_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21904),
            .ce(N__21591),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_5_6_LC_15_21_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_5_6_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_5_6_LC_15_21_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \c0.tx2_data_RNO_5_6_LC_15_21_5  (
            .in0(N__20920),
            .in1(N__18437),
            .in2(_gnd_net_),
            .in3(N__18369),
            .lcout(\c0.tx2_data_1_iv_4_1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__6_LC_15_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__6_LC_15_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__6_LC_15_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__6_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19870),
            .lcout(\c0.data_in_frame_7_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21904),
            .ce(N__21591),
            .sr(_gnd_net_));
    defparam \c0.d_4_RNI09QE_46_LC_15_21_7 .C_ON=1'b0;
    defparam \c0.d_4_RNI09QE_46_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.d_4_RNI09QE_46_LC_15_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.d_4_RNI09QE_46_LC_15_21_7  (
            .in0(N__22017),
            .in1(N__18419),
            .in2(_gnd_net_),
            .in3(N__18368),
            .lcout(\c0.un1_data_in_7__2_0_a2_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__4_LC_15_22_0 .C_ON=1'b0;
    defparam \c0.data_in_7__4_LC_15_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__4_LC_15_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__4_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21509),
            .lcout(\c0.data_in_7_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__2_LC_15_22_1 .C_ON=1'b0;
    defparam \c0.data_in_7__2_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__2_LC_15_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__2_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21526),
            .lcout(\c0.data_in_7_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__7_LC_15_22_2 .C_ON=1'b0;
    defparam \c0.data_in_4__7_LC_15_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__7_LC_15_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__7_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20665),
            .lcout(\c0.data_in_4_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__7_LC_15_22_3 .C_ON=1'b0;
    defparam \c0.data_in_7__7_LC_15_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__7_LC_15_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__7_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18827),
            .lcout(\c0.data_in_7_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__1_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.data_in_6__1_LC_15_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__1_LC_15_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__1_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22069),
            .lcout(\c0.data_in_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__0_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.data_in_6__0_LC_15_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__0_LC_15_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__0_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18742),
            .lcout(\c0.data_in_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__0_LC_15_22_6 .C_ON=1'b0;
    defparam \c0.data_in_7__0_LC_15_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__0_LC_15_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__0_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21071),
            .lcout(\c0.data_in_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__4_LC_15_22_7 .C_ON=1'b0;
    defparam \c0.data_in_5__4_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__4_LC_15_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__4_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22270),
            .lcout(\c0.data_in_5_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21911),
            .ce(N__22161),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5_LC_15_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5_LC_15_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_5_LC_15_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_5_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21919),
            .ce(N__19029),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_2_LC_15_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_2_LC_15_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_2_LC_15_23_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \c0.byte_transmit_counter_2_LC_15_23_2  (
            .in0(N__19113),
            .in1(N__19430),
            .in2(_gnd_net_),
            .in3(N__19320),
            .lcout(\c0.byte_transmit_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21919),
            .ce(N__19029),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_7_LC_15_23_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_7_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_7_LC_15_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.byte_transmit_counter_7_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\c0.byte_transmit_counterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21919),
            .ce(N__19029),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__5_LC_15_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__5_LC_15_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__5_LC_15_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__5_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19927),
            .lcout(\c0.data_in_frame_6_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21927),
            .ce(N__21598),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_3_LC_16_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_3_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_3_LC_16_17_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \c0.byte_transmit_counter2_3_LC_16_17_0  (
            .in0(N__21059),
            .in1(N__21039),
            .in2(_gnd_net_),
            .in3(N__20082),
            .lcout(\c0.byte_transmit_counter2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21878),
            .ce(),
            .sr(N__20046));
    defparam \c0.tx2_data_RNO_2_4_LC_16_18_0 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_4_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_4_LC_16_18_0 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \c0.tx2_data_RNO_2_4_LC_16_18_0  (
            .in0(N__20388),
            .in1(N__19676),
            .in2(N__18998),
            .in3(N__20279),
            .lcout(\c0.tx2_data_1_iv_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIJFIT_0_LC_16_18_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIJFIT_0_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIJFIT_0_LC_16_18_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.byte_transmit_counter2_RNIJFIT_0_LC_16_18_1  (
            .in0(N__20831),
            .in1(N__19482),
            .in2(_gnd_net_),
            .in3(N__18873),
            .lcout(\c0.N_207 ),
            .ltout(\c0.N_207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_4_LC_16_18_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_4_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_4_LC_16_18_2 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \c0.tx2_data_RNO_0_4_LC_16_18_2  (
            .in0(N__21944),
            .in1(N__20278),
            .in2(N__18971),
            .in3(N__18968),
            .lcout(\c0.tx2_data_1_0_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIBNLC_7_LC_16_18_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIBNLC_7_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIBNLC_7_LC_16_18_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.byte_transmit_counter2_RNIBNLC_7_LC_16_18_3  (
            .in0(N__21032),
            .in1(N__19666),
            .in2(_gnd_net_),
            .in3(N__21005),
            .lcout(\c0.m2_e_0_2 ),
            .ltout(\c0.m2_e_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIK84L_6_LC_16_18_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIK84L_6_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIK84L_6_LC_16_18_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \c0.byte_transmit_counter2_RNIK84L_6_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__19630),
            .in2(N__18932),
            .in3(N__19599),
            .lcout(\c0.N_71_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_LC_16_18_5 .C_ON=1'b0;
    defparam \c0.tx2_transmit_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_LC_16_18_5 .LUT_INIT=16'b0011000000111001;
    LogicCell40 \c0.tx2_transmit_LC_16_18_5  (
            .in0(N__19850),
            .in1(N__19826),
            .in2(N__19811),
            .in3(N__19769),
            .lcout(\c0.tx2_transmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21886),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNIJBBP_0_6_LC_16_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNIJBBP_0_6_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNIJBBP_0_6_LC_16_18_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.byte_transmit_counter2_RNIJBBP_0_6_LC_16_18_6  (
            .in0(N__19481),
            .in1(N__19739),
            .in2(N__19649),
            .in3(N__19600),
            .lcout(\c0.N_203 ),
            .ltout(\c0.N_203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_3_4_LC_16_18_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_3_4_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_3_4_LC_16_18_7 .LUT_INIT=16'b0010111101111111;
    LogicCell40 \c0.tx2_data_RNO_3_4_LC_16_18_7  (
            .in0(N__20832),
            .in1(N__19727),
            .in2(N__19697),
            .in3(N__19694),
            .lcout(\c0.tx2_data_1_iv_5_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNO_1_7_LC_16_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNO_1_7_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNO_1_7_LC_16_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.byte_transmit_counter2_RNO_1_7_LC_16_19_0  (
            .in0(N__20858),
            .in1(N__21009),
            .in2(N__20325),
            .in3(N__21040),
            .lcout(),
            .ltout(\c0.un1_m4_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_7_LC_16_19_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_7_LC_16_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_7_LC_16_19_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \c0.byte_transmit_counter2_7_LC_16_19_1  (
            .in0(N__19655),
            .in1(N__19667),
            .in2(N__19670),
            .in3(N__20086),
            .lcout(\c0.byte_transmit_counter2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21895),
            .ce(),
            .sr(N__20054));
    defparam \c0.byte_transmit_counter2_RNO_0_7_LC_16_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNO_0_7_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNO_0_7_LC_16_19_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.byte_transmit_counter2_RNO_0_7_LC_16_19_2  (
            .in0(N__19484),
            .in1(N__19637),
            .in2(_gnd_net_),
            .in3(N__19604),
            .lcout(\c0.un1_m4_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_6_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_6_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_6_LC_16_19_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \c0.byte_transmit_counter2_6_LC_16_19_3  (
            .in0(N__20983),
            .in1(N__19606),
            .in2(N__19647),
            .in3(N__20085),
            .lcout(\c0.byte_transmit_counter2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21895),
            .ce(),
            .sr(N__20054));
    defparam \c0.byte_transmit_counter2_5_LC_16_19_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_5_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_5_LC_16_19_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \c0.byte_transmit_counter2_5_LC_16_19_5  (
            .in0(N__19605),
            .in1(_gnd_net_),
            .in2(N__20984),
            .in3(N__20084),
            .lcout(\c0.byte_transmit_counter2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21895),
            .ce(),
            .sr(N__20054));
    defparam \c0.byte_transmit_counter2_RNI0CLC_0_LC_16_19_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNI0CLC_0_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNI0CLC_0_LC_16_19_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.byte_transmit_counter2_RNI0CLC_0_LC_16_19_6  (
            .in0(N__19483),
            .in1(_gnd_net_),
            .in2(N__20324),
            .in3(N__20843),
            .lcout(\c0.un1_byte_transmit_counter2_1_ac0_3_out ),
            .ltout(\c0.un1_byte_transmit_counter2_1_ac0_3_out_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4_LC_16_19_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4_LC_16_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_4_LC_16_19_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \c0.byte_transmit_counter2_4_LC_16_19_7  (
            .in0(N__21041),
            .in1(N__21010),
            .in2(N__20090),
            .in3(N__20083),
            .lcout(\c0.byte_transmit_counter2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21895),
            .ce(),
            .sr(N__20054));
    defparam \c0.data_in_4__5_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.data_in_4__5_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__5_LC_16_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__5_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19978),
            .lcout(\c0.data_in_4_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__5_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.data_in_5__5_LC_16_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__5_LC_16_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__5_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19914),
            .lcout(\c0.data_in_5_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__5_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.data_in_6__5_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__5_LC_16_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__5_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19963),
            .lcout(\c0.data_in_6_Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__2_LC_16_20_3 .C_ON=1'b0;
    defparam \c0.data_in_6__2_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__2_LC_16_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__2_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22018),
            .lcout(\c0.data_in_6_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_4__6_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.data_in_4__6_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_4__6_LC_16_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_4__6_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19888),
            .lcout(\c0.data_in_4_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__6_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.data_in_5__6_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__6_LC_16_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_5__6_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20583),
            .lcout(\c0.data_in_5_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__6_LC_16_20_6 .C_ON=1'b0;
    defparam \c0.data_in_6__6_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__6_LC_16_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__6_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19869),
            .lcout(\c0.data_in_6_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_7__6_LC_16_20_7 .C_ON=1'b0;
    defparam \c0.data_in_7__6_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_7__6_LC_16_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_7__6_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20108),
            .lcout(\c0.data_in_7_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21905),
            .ce(N__22160),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__3_LC_16_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__3_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__3_LC_16_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__3_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20642),
            .lcout(\c0.data_in_frame_6_Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21912),
            .ce(N__21588),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_0_6_LC_16_21_2 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_0_6_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_0_6_LC_16_21_2 .LUT_INIT=16'b0011101101111111;
    LogicCell40 \c0.tx2_data_RNO_0_6_LC_16_21_2  (
            .in0(N__20923),
            .in1(N__20390),
            .in2(N__20564),
            .in3(N__20515),
            .lcout(\c0.tx2_data_1_0_i_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__6_LC_16_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__6_LC_16_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__6_LC_16_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__6_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20584),
            .lcout(\c0.data_in_frame_6_Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21912),
            .ce(N__21588),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_4__6_LC_16_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_4__6_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_4__6_LC_16_21_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.data_in_frame_4__6_LC_16_21_4  (
            .in0(N__20545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.d_4_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21912),
            .ce(N__21588),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_4_5_LC_16_21_5 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_4_5_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_4_5_LC_16_21_5 .LUT_INIT=16'b0101111101110111;
    LogicCell40 \c0.tx2_data_RNO_4_5_LC_16_21_5  (
            .in0(N__20389),
            .in1(N__20474),
            .in2(N__20450),
            .in3(N__20922),
            .lcout(),
            .ltout(\c0.tx2_data_1_iv_5_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_2_5_LC_16_21_6 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_2_5_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_2_5_LC_16_21_6 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \c0.tx2_data_RNO_2_5_LC_16_21_6  (
            .in0(N__20126),
            .in1(N__20391),
            .in2(N__20360),
            .in3(N__20328),
            .lcout(\c0.tx2_data_1_iv_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_data_RNO_5_5_LC_16_21_7 .C_ON=1'b0;
    defparam \c0.tx2_data_RNO_5_5_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2_data_RNO_5_5_LC_16_21_7 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \c0.tx2_data_RNO_5_5_LC_16_21_7  (
            .in0(N__20177),
            .in1(N__20921),
            .in2(_gnd_net_),
            .in3(N__20168),
            .lcout(\c0.tx2_data_1_iv_5_1_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_6_LC_16_22_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_6_LC_16_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_6_LC_16_22_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_6_LC_16_22_1  (
            .in0(N__21245),
            .in1(N__20120),
            .in2(N__20107),
            .in3(N__21144),
            .lcout(\c0.rx_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21920),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_2_LC_16_22_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_2_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_2_LC_16_22_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.rx.r_Rx_Byte_2_LC_16_22_2  (
            .in0(N__21142),
            .in1(N__21536),
            .in2(N__21527),
            .in3(N__21243),
            .lcout(\c0.rx_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21920),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_4_LC_16_22_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_4_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_4_LC_16_22_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_4_LC_16_22_3  (
            .in0(N__21326),
            .in1(_gnd_net_),
            .in2(N__21412),
            .in3(N__21496),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_4_LC_16_22_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_4_LC_16_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_4_LC_16_22_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \c0.rx.r_Rx_Byte_4_LC_16_22_4  (
            .in0(N__21143),
            .in1(N__21508),
            .in2(N__21512),
            .in3(N__21244),
            .lcout(\c0.rx_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21920),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_RNO_0_0_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_RNO_0_0_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_Rx_Byte_RNO_0_0_LC_16_22_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \c0.rx.r_Rx_Byte_RNO_0_0_LC_16_22_6  (
            .in0(N__21495),
            .in1(N__21403),
            .in2(_gnd_net_),
            .in3(N__21325),
            .lcout(),
            .ltout(\c0.rx.r_Rx_Bytece_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_0_LC_16_22_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_0_LC_16_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_0_LC_16_22_7 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_0_LC_16_22_7  (
            .in0(N__21242),
            .in1(N__21070),
            .in2(N__21149),
            .in3(N__21141),
            .lcout(\c0.rx_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21920),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_RNI5P3L_4_LC_17_17_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_RNI5P3L_4_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_RNI5P3L_4_LC_17_17_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.byte_transmit_counter2_RNI5P3L_4_LC_17_17_7  (
            .in0(N__21058),
            .in1(N__21033),
            .in2(_gnd_net_),
            .in3(N__21011),
            .lcout(\c0.un1_byte_transmit_counter2_1_ac0_7_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_4_LC_17_18_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_4_LC_17_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_4_LC_17_18_6 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \c0.tx2.r_Tx_Data_4_LC_17_18_6  (
            .in0(N__20969),
            .in1(N__20963),
            .in2(N__20957),
            .in3(N__20878),
            .lcout(\c0.tx2.r_Tx_DataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21896),
            .ce(N__20733),
            .sr(_gnd_net_));
    defparam \c0.data_in_5__7_LC_17_20_0 .C_ON=1'b0;
    defparam \c0.data_in_5__7_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_5__7_LC_17_20_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.data_in_5__7_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__22190),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_5_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21913),
            .ce(N__22162),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__4_LC_17_21_0 .C_ON=1'b0;
    defparam \c0.data_in_6__4_LC_17_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__4_LC_17_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__4_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21975),
            .lcout(\c0.data_in_6_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21921),
            .ce(N__22163),
            .sr(_gnd_net_));
    defparam \c0.data_in_6__7_LC_17_21_1 .C_ON=1'b0;
    defparam \c0.data_in_6__7_LC_17_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_6__7_LC_17_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_6__7_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22234),
            .lcout(\c0.data_in_6_Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21921),
            .ce(N__22163),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_6__2_LC_18_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_6__2_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_6__2_LC_18_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_6__2_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22111),
            .lcout(\c0.data_in_frame_6_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21922),
            .ce(N__21581),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__1_LC_18_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__1_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__1_LC_18_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__1_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22073),
            .lcout(\c0.data_in_frame_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21928),
            .ce(N__21582),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__2_LC_18_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__2_LC_18_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__2_LC_18_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__2_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22022),
            .lcout(\c0.data_in_frame_7_Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21928),
            .ce(N__21582),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_7__4_LC_18_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_7__4_LC_18_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_7__4_LC_18_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.data_in_frame_7__4_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21976),
            .lcout(\c0.data_in_frame_7_Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21928),
            .ce(N__21582),
            .sr(_gnd_net_));
endmodule // top
