// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 19 2019 16:12:29

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    output PIN_9;
    input PIN_8;
    input PIN_7;
    inout PIN_6;
    inout PIN_5;
    inout PIN_4;
    output PIN_3;
    output PIN_24;
    output PIN_23;
    output PIN_22;
    input PIN_21;
    input PIN_20;
    output PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    inout PIN_11;
    inout PIN_10;
    output PIN_1;
    output LED;
    input CLK;

    wire N__101572;
    wire N__101571;
    wire N__101570;
    wire N__101563;
    wire N__101562;
    wire N__101561;
    wire N__101554;
    wire N__101553;
    wire N__101552;
    wire N__101545;
    wire N__101544;
    wire N__101543;
    wire N__101536;
    wire N__101535;
    wire N__101534;
    wire N__101527;
    wire N__101526;
    wire N__101525;
    wire N__101518;
    wire N__101517;
    wire N__101516;
    wire N__101509;
    wire N__101508;
    wire N__101507;
    wire N__101500;
    wire N__101499;
    wire N__101498;
    wire N__101491;
    wire N__101490;
    wire N__101489;
    wire N__101482;
    wire N__101481;
    wire N__101480;
    wire N__101473;
    wire N__101472;
    wire N__101471;
    wire N__101464;
    wire N__101463;
    wire N__101462;
    wire N__101455;
    wire N__101454;
    wire N__101453;
    wire N__101446;
    wire N__101445;
    wire N__101444;
    wire N__101437;
    wire N__101436;
    wire N__101435;
    wire N__101428;
    wire N__101427;
    wire N__101426;
    wire N__101419;
    wire N__101418;
    wire N__101417;
    wire N__101410;
    wire N__101409;
    wire N__101408;
    wire N__101391;
    wire N__101388;
    wire N__101387;
    wire N__101384;
    wire N__101381;
    wire N__101380;
    wire N__101377;
    wire N__101374;
    wire N__101373;
    wire N__101370;
    wire N__101367;
    wire N__101364;
    wire N__101361;
    wire N__101358;
    wire N__101349;
    wire N__101348;
    wire N__101347;
    wire N__101344;
    wire N__101343;
    wire N__101342;
    wire N__101341;
    wire N__101338;
    wire N__101337;
    wire N__101336;
    wire N__101335;
    wire N__101334;
    wire N__101331;
    wire N__101328;
    wire N__101325;
    wire N__101322;
    wire N__101321;
    wire N__101318;
    wire N__101315;
    wire N__101312;
    wire N__101307;
    wire N__101304;
    wire N__101299;
    wire N__101296;
    wire N__101295;
    wire N__101294;
    wire N__101291;
    wire N__101286;
    wire N__101281;
    wire N__101278;
    wire N__101277;
    wire N__101274;
    wire N__101271;
    wire N__101270;
    wire N__101267;
    wire N__101262;
    wire N__101255;
    wire N__101252;
    wire N__101249;
    wire N__101246;
    wire N__101243;
    wire N__101240;
    wire N__101235;
    wire N__101232;
    wire N__101229;
    wire N__101226;
    wire N__101221;
    wire N__101214;
    wire N__101205;
    wire N__101204;
    wire N__101203;
    wire N__101202;
    wire N__101201;
    wire N__101198;
    wire N__101197;
    wire N__101196;
    wire N__101191;
    wire N__101190;
    wire N__101189;
    wire N__101188;
    wire N__101185;
    wire N__101182;
    wire N__101179;
    wire N__101176;
    wire N__101173;
    wire N__101170;
    wire N__101165;
    wire N__101162;
    wire N__101159;
    wire N__101156;
    wire N__101151;
    wire N__101148;
    wire N__101145;
    wire N__101142;
    wire N__101137;
    wire N__101134;
    wire N__101131;
    wire N__101128;
    wire N__101119;
    wire N__101112;
    wire N__101111;
    wire N__101110;
    wire N__101107;
    wire N__101102;
    wire N__101101;
    wire N__101100;
    wire N__101099;
    wire N__101096;
    wire N__101093;
    wire N__101090;
    wire N__101089;
    wire N__101084;
    wire N__101079;
    wire N__101076;
    wire N__101073;
    wire N__101070;
    wire N__101067;
    wire N__101058;
    wire N__101055;
    wire N__101054;
    wire N__101051;
    wire N__101050;
    wire N__101047;
    wire N__101046;
    wire N__101045;
    wire N__101042;
    wire N__101039;
    wire N__101038;
    wire N__101035;
    wire N__101032;
    wire N__101029;
    wire N__101024;
    wire N__101021;
    wire N__101018;
    wire N__101011;
    wire N__101006;
    wire N__101001;
    wire N__101000;
    wire N__100999;
    wire N__100992;
    wire N__100991;
    wire N__100990;
    wire N__100987;
    wire N__100986;
    wire N__100983;
    wire N__100980;
    wire N__100977;
    wire N__100974;
    wire N__100965;
    wire N__100962;
    wire N__100959;
    wire N__100958;
    wire N__100957;
    wire N__100954;
    wire N__100953;
    wire N__100950;
    wire N__100947;
    wire N__100944;
    wire N__100941;
    wire N__100940;
    wire N__100937;
    wire N__100930;
    wire N__100929;
    wire N__100926;
    wire N__100923;
    wire N__100920;
    wire N__100917;
    wire N__100914;
    wire N__100911;
    wire N__100908;
    wire N__100905;
    wire N__100896;
    wire N__100895;
    wire N__100890;
    wire N__100887;
    wire N__100884;
    wire N__100881;
    wire N__100880;
    wire N__100879;
    wire N__100878;
    wire N__100875;
    wire N__100874;
    wire N__100871;
    wire N__100868;
    wire N__100867;
    wire N__100866;
    wire N__100863;
    wire N__100860;
    wire N__100857;
    wire N__100852;
    wire N__100847;
    wire N__100836;
    wire N__100833;
    wire N__100832;
    wire N__100827;
    wire N__100826;
    wire N__100825;
    wire N__100824;
    wire N__100821;
    wire N__100818;
    wire N__100815;
    wire N__100812;
    wire N__100807;
    wire N__100806;
    wire N__100801;
    wire N__100798;
    wire N__100795;
    wire N__100792;
    wire N__100789;
    wire N__100782;
    wire N__100781;
    wire N__100780;
    wire N__100777;
    wire N__100776;
    wire N__100773;
    wire N__100772;
    wire N__100769;
    wire N__100766;
    wire N__100763;
    wire N__100760;
    wire N__100757;
    wire N__100754;
    wire N__100751;
    wire N__100750;
    wire N__100747;
    wire N__100742;
    wire N__100739;
    wire N__100736;
    wire N__100733;
    wire N__100730;
    wire N__100727;
    wire N__100726;
    wire N__100723;
    wire N__100720;
    wire N__100717;
    wire N__100714;
    wire N__100711;
    wire N__100708;
    wire N__100701;
    wire N__100696;
    wire N__100689;
    wire N__100686;
    wire N__100685;
    wire N__100684;
    wire N__100683;
    wire N__100682;
    wire N__100679;
    wire N__100674;
    wire N__100671;
    wire N__100670;
    wire N__100667;
    wire N__100662;
    wire N__100659;
    wire N__100656;
    wire N__100653;
    wire N__100650;
    wire N__100647;
    wire N__100642;
    wire N__100639;
    wire N__100632;
    wire N__100631;
    wire N__100628;
    wire N__100625;
    wire N__100620;
    wire N__100619;
    wire N__100616;
    wire N__100615;
    wire N__100612;
    wire N__100609;
    wire N__100606;
    wire N__100599;
    wire N__100596;
    wire N__100593;
    wire N__100590;
    wire N__100589;
    wire N__100586;
    wire N__100585;
    wire N__100582;
    wire N__100579;
    wire N__100576;
    wire N__100569;
    wire N__100568;
    wire N__100567;
    wire N__100564;
    wire N__100561;
    wire N__100558;
    wire N__100551;
    wire N__100550;
    wire N__100549;
    wire N__100546;
    wire N__100543;
    wire N__100540;
    wire N__100533;
    wire N__100530;
    wire N__100529;
    wire N__100526;
    wire N__100523;
    wire N__100520;
    wire N__100519;
    wire N__100514;
    wire N__100511;
    wire N__100506;
    wire N__100505;
    wire N__100504;
    wire N__100503;
    wire N__100500;
    wire N__100497;
    wire N__100494;
    wire N__100491;
    wire N__100488;
    wire N__100485;
    wire N__100480;
    wire N__100473;
    wire N__100470;
    wire N__100469;
    wire N__100468;
    wire N__100467;
    wire N__100466;
    wire N__100465;
    wire N__100462;
    wire N__100459;
    wire N__100456;
    wire N__100453;
    wire N__100450;
    wire N__100447;
    wire N__100442;
    wire N__100433;
    wire N__100428;
    wire N__100427;
    wire N__100426;
    wire N__100425;
    wire N__100422;
    wire N__100419;
    wire N__100416;
    wire N__100415;
    wire N__100414;
    wire N__100411;
    wire N__100406;
    wire N__100403;
    wire N__100400;
    wire N__100397;
    wire N__100392;
    wire N__100389;
    wire N__100380;
    wire N__100379;
    wire N__100376;
    wire N__100373;
    wire N__100370;
    wire N__100367;
    wire N__100364;
    wire N__100359;
    wire N__100358;
    wire N__100357;
    wire N__100354;
    wire N__100351;
    wire N__100348;
    wire N__100345;
    wire N__100342;
    wire N__100339;
    wire N__100336;
    wire N__100331;
    wire N__100326;
    wire N__100323;
    wire N__100320;
    wire N__100319;
    wire N__100316;
    wire N__100313;
    wire N__100308;
    wire N__100305;
    wire N__100304;
    wire N__100301;
    wire N__100298;
    wire N__100295;
    wire N__100290;
    wire N__100287;
    wire N__100284;
    wire N__100281;
    wire N__100280;
    wire N__100277;
    wire N__100274;
    wire N__100269;
    wire N__100268;
    wire N__100263;
    wire N__100260;
    wire N__100257;
    wire N__100256;
    wire N__100255;
    wire N__100254;
    wire N__100253;
    wire N__100250;
    wire N__100247;
    wire N__100246;
    wire N__100243;
    wire N__100240;
    wire N__100237;
    wire N__100234;
    wire N__100231;
    wire N__100228;
    wire N__100225;
    wire N__100222;
    wire N__100219;
    wire N__100216;
    wire N__100213;
    wire N__100210;
    wire N__100207;
    wire N__100206;
    wire N__100203;
    wire N__100198;
    wire N__100195;
    wire N__100190;
    wire N__100187;
    wire N__100182;
    wire N__100179;
    wire N__100176;
    wire N__100167;
    wire N__100166;
    wire N__100165;
    wire N__100162;
    wire N__100161;
    wire N__100160;
    wire N__100159;
    wire N__100156;
    wire N__100153;
    wire N__100150;
    wire N__100143;
    wire N__100140;
    wire N__100137;
    wire N__100134;
    wire N__100131;
    wire N__100128;
    wire N__100123;
    wire N__100116;
    wire N__100113;
    wire N__100110;
    wire N__100107;
    wire N__100104;
    wire N__100103;
    wire N__100102;
    wire N__100101;
    wire N__100100;
    wire N__100099;
    wire N__100094;
    wire N__100091;
    wire N__100088;
    wire N__100083;
    wire N__100082;
    wire N__100079;
    wire N__100078;
    wire N__100071;
    wire N__100070;
    wire N__100067;
    wire N__100064;
    wire N__100061;
    wire N__100058;
    wire N__100055;
    wire N__100052;
    wire N__100041;
    wire N__100038;
    wire N__100035;
    wire N__100034;
    wire N__100031;
    wire N__100028;
    wire N__100027;
    wire N__100024;
    wire N__100021;
    wire N__100018;
    wire N__100011;
    wire N__100008;
    wire N__100005;
    wire N__100002;
    wire N__99999;
    wire N__99996;
    wire N__99995;
    wire N__99994;
    wire N__99991;
    wire N__99990;
    wire N__99987;
    wire N__99986;
    wire N__99983;
    wire N__99982;
    wire N__99981;
    wire N__99978;
    wire N__99975;
    wire N__99970;
    wire N__99963;
    wire N__99954;
    wire N__99953;
    wire N__99952;
    wire N__99949;
    wire N__99946;
    wire N__99943;
    wire N__99936;
    wire N__99933;
    wire N__99930;
    wire N__99929;
    wire N__99926;
    wire N__99923;
    wire N__99922;
    wire N__99917;
    wire N__99916;
    wire N__99913;
    wire N__99910;
    wire N__99907;
    wire N__99904;
    wire N__99901;
    wire N__99894;
    wire N__99891;
    wire N__99888;
    wire N__99887;
    wire N__99886;
    wire N__99883;
    wire N__99880;
    wire N__99877;
    wire N__99870;
    wire N__99869;
    wire N__99868;
    wire N__99865;
    wire N__99862;
    wire N__99859;
    wire N__99856;
    wire N__99853;
    wire N__99846;
    wire N__99843;
    wire N__99840;
    wire N__99839;
    wire N__99836;
    wire N__99833;
    wire N__99832;
    wire N__99829;
    wire N__99826;
    wire N__99823;
    wire N__99816;
    wire N__99813;
    wire N__99810;
    wire N__99809;
    wire N__99808;
    wire N__99805;
    wire N__99802;
    wire N__99799;
    wire N__99792;
    wire N__99789;
    wire N__99786;
    wire N__99783;
    wire N__99780;
    wire N__99779;
    wire N__99778;
    wire N__99775;
    wire N__99772;
    wire N__99769;
    wire N__99762;
    wire N__99761;
    wire N__99760;
    wire N__99759;
    wire N__99758;
    wire N__99757;
    wire N__99754;
    wire N__99751;
    wire N__99748;
    wire N__99747;
    wire N__99746;
    wire N__99741;
    wire N__99738;
    wire N__99727;
    wire N__99720;
    wire N__99717;
    wire N__99714;
    wire N__99711;
    wire N__99710;
    wire N__99707;
    wire N__99704;
    wire N__99699;
    wire N__99696;
    wire N__99695;
    wire N__99692;
    wire N__99689;
    wire N__99688;
    wire N__99683;
    wire N__99680;
    wire N__99675;
    wire N__99672;
    wire N__99671;
    wire N__99668;
    wire N__99665;
    wire N__99662;
    wire N__99659;
    wire N__99654;
    wire N__99651;
    wire N__99648;
    wire N__99645;
    wire N__99642;
    wire N__99639;
    wire N__99638;
    wire N__99635;
    wire N__99632;
    wire N__99629;
    wire N__99624;
    wire N__99621;
    wire N__99618;
    wire N__99615;
    wire N__99612;
    wire N__99609;
    wire N__99606;
    wire N__99605;
    wire N__99604;
    wire N__99603;
    wire N__99602;
    wire N__99601;
    wire N__99600;
    wire N__99597;
    wire N__99596;
    wire N__99593;
    wire N__99592;
    wire N__99589;
    wire N__99588;
    wire N__99587;
    wire N__99586;
    wire N__99585;
    wire N__99584;
    wire N__99583;
    wire N__99582;
    wire N__99581;
    wire N__99580;
    wire N__99577;
    wire N__99576;
    wire N__99573;
    wire N__99572;
    wire N__99569;
    wire N__99568;
    wire N__99567;
    wire N__99566;
    wire N__99565;
    wire N__99564;
    wire N__99563;
    wire N__99562;
    wire N__99561;
    wire N__99560;
    wire N__99559;
    wire N__99558;
    wire N__99543;
    wire N__99536;
    wire N__99527;
    wire N__99512;
    wire N__99511;
    wire N__99510;
    wire N__99509;
    wire N__99508;
    wire N__99505;
    wire N__99504;
    wire N__99501;
    wire N__99500;
    wire N__99497;
    wire N__99496;
    wire N__99495;
    wire N__99494;
    wire N__99493;
    wire N__99492;
    wire N__99491;
    wire N__99490;
    wire N__99489;
    wire N__99488;
    wire N__99485;
    wire N__99484;
    wire N__99481;
    wire N__99480;
    wire N__99477;
    wire N__99476;
    wire N__99475;
    wire N__99474;
    wire N__99473;
    wire N__99472;
    wire N__99471;
    wire N__99470;
    wire N__99469;
    wire N__99468;
    wire N__99467;
    wire N__99458;
    wire N__99449;
    wire N__99442;
    wire N__99427;
    wire N__99420;
    wire N__99411;
    wire N__99396;
    wire N__99395;
    wire N__99392;
    wire N__99391;
    wire N__99388;
    wire N__99387;
    wire N__99384;
    wire N__99383;
    wire N__99382;
    wire N__99379;
    wire N__99378;
    wire N__99375;
    wire N__99374;
    wire N__99371;
    wire N__99370;
    wire N__99369;
    wire N__99368;
    wire N__99367;
    wire N__99366;
    wire N__99365;
    wire N__99364;
    wire N__99363;
    wire N__99362;
    wire N__99359;
    wire N__99358;
    wire N__99355;
    wire N__99354;
    wire N__99351;
    wire N__99350;
    wire N__99349;
    wire N__99348;
    wire N__99347;
    wire N__99346;
    wire N__99345;
    wire N__99344;
    wire N__99343;
    wire N__99342;
    wire N__99341;
    wire N__99340;
    wire N__99339;
    wire N__99338;
    wire N__99337;
    wire N__99336;
    wire N__99335;
    wire N__99334;
    wire N__99333;
    wire N__99332;
    wire N__99331;
    wire N__99330;
    wire N__99327;
    wire N__99314;
    wire N__99299;
    wire N__99284;
    wire N__99277;
    wire N__99268;
    wire N__99253;
    wire N__99252;
    wire N__99249;
    wire N__99248;
    wire N__99245;
    wire N__99244;
    wire N__99241;
    wire N__99240;
    wire N__99239;
    wire N__99236;
    wire N__99235;
    wire N__99232;
    wire N__99231;
    wire N__99228;
    wire N__99227;
    wire N__99226;
    wire N__99225;
    wire N__99224;
    wire N__99223;
    wire N__99222;
    wire N__99221;
    wire N__99220;
    wire N__99219;
    wire N__99216;
    wire N__99215;
    wire N__99212;
    wire N__99211;
    wire N__99208;
    wire N__99207;
    wire N__99206;
    wire N__99205;
    wire N__99204;
    wire N__99203;
    wire N__99202;
    wire N__99201;
    wire N__99200;
    wire N__99197;
    wire N__99196;
    wire N__99193;
    wire N__99192;
    wire N__99189;
    wire N__99188;
    wire N__99187;
    wire N__99184;
    wire N__99183;
    wire N__99180;
    wire N__99179;
    wire N__99176;
    wire N__99175;
    wire N__99174;
    wire N__99171;
    wire N__99170;
    wire N__99167;
    wire N__99166;
    wire N__99163;
    wire N__99162;
    wire N__99161;
    wire N__99158;
    wire N__99155;
    wire N__99154;
    wire N__99153;
    wire N__99152;
    wire N__99151;
    wire N__99150;
    wire N__99149;
    wire N__99148;
    wire N__99147;
    wire N__99146;
    wire N__99131;
    wire N__99116;
    wire N__99101;
    wire N__99094;
    wire N__99085;
    wire N__99070;
    wire N__99069;
    wire N__99068;
    wire N__99067;
    wire N__99066;
    wire N__99065;
    wire N__99064;
    wire N__99063;
    wire N__99062;
    wire N__99059;
    wire N__99058;
    wire N__99055;
    wire N__99054;
    wire N__99051;
    wire N__99050;
    wire N__99049;
    wire N__99048;
    wire N__99047;
    wire N__99046;
    wire N__99045;
    wire N__99044;
    wire N__99043;
    wire N__99042;
    wire N__99039;
    wire N__99038;
    wire N__99035;
    wire N__99034;
    wire N__99031;
    wire N__99030;
    wire N__99029;
    wire N__99028;
    wire N__99027;
    wire N__99012;
    wire N__98997;
    wire N__98982;
    wire N__98981;
    wire N__98980;
    wire N__98979;
    wire N__98978;
    wire N__98977;
    wire N__98976;
    wire N__98975;
    wire N__98974;
    wire N__98973;
    wire N__98972;
    wire N__98967;
    wire N__98966;
    wire N__98965;
    wire N__98962;
    wire N__98961;
    wire N__98958;
    wire N__98957;
    wire N__98954;
    wire N__98953;
    wire N__98950;
    wire N__98949;
    wire N__98944;
    wire N__98941;
    wire N__98940;
    wire N__98939;
    wire N__98938;
    wire N__98937;
    wire N__98934;
    wire N__98933;
    wire N__98930;
    wire N__98929;
    wire N__98926;
    wire N__98925;
    wire N__98912;
    wire N__98903;
    wire N__98896;
    wire N__98881;
    wire N__98874;
    wire N__98865;
    wire N__98850;
    wire N__98849;
    wire N__98846;
    wire N__98845;
    wire N__98842;
    wire N__98841;
    wire N__98838;
    wire N__98837;
    wire N__98830;
    wire N__98821;
    wire N__98820;
    wire N__98817;
    wire N__98816;
    wire N__98813;
    wire N__98812;
    wire N__98809;
    wire N__98808;
    wire N__98807;
    wire N__98806;
    wire N__98805;
    wire N__98804;
    wire N__98803;
    wire N__98802;
    wire N__98801;
    wire N__98800;
    wire N__98797;
    wire N__98796;
    wire N__98793;
    wire N__98792;
    wire N__98789;
    wire N__98788;
    wire N__98785;
    wire N__98782;
    wire N__98781;
    wire N__98780;
    wire N__98779;
    wire N__98778;
    wire N__98777;
    wire N__98774;
    wire N__98771;
    wire N__98756;
    wire N__98755;
    wire N__98754;
    wire N__98753;
    wire N__98752;
    wire N__98751;
    wire N__98750;
    wire N__98749;
    wire N__98748;
    wire N__98743;
    wire N__98736;
    wire N__98721;
    wire N__98716;
    wire N__98705;
    wire N__98690;
    wire N__98685;
    wire N__98670;
    wire N__98663;
    wire N__98654;
    wire N__98639;
    wire N__98636;
    wire N__98633;
    wire N__98632;
    wire N__98629;
    wire N__98628;
    wire N__98625;
    wire N__98624;
    wire N__98621;
    wire N__98620;
    wire N__98617;
    wire N__98614;
    wire N__98611;
    wire N__98606;
    wire N__98599;
    wire N__98590;
    wire N__98589;
    wire N__98586;
    wire N__98583;
    wire N__98578;
    wire N__98561;
    wire N__98556;
    wire N__98541;
    wire N__98538;
    wire N__98535;
    wire N__98532;
    wire N__98525;
    wire N__98522;
    wire N__98519;
    wire N__98518;
    wire N__98515;
    wire N__98510;
    wire N__98505;
    wire N__98500;
    wire N__98491;
    wire N__98488;
    wire N__98475;
    wire N__98472;
    wire N__98469;
    wire N__98468;
    wire N__98465;
    wire N__98462;
    wire N__98457;
    wire N__98454;
    wire N__98451;
    wire N__98450;
    wire N__98449;
    wire N__98448;
    wire N__98447;
    wire N__98446;
    wire N__98445;
    wire N__98442;
    wire N__98437;
    wire N__98434;
    wire N__98431;
    wire N__98426;
    wire N__98419;
    wire N__98412;
    wire N__98409;
    wire N__98406;
    wire N__98403;
    wire N__98400;
    wire N__98397;
    wire N__98394;
    wire N__98391;
    wire N__98390;
    wire N__98387;
    wire N__98384;
    wire N__98381;
    wire N__98378;
    wire N__98373;
    wire N__98370;
    wire N__98369;
    wire N__98366;
    wire N__98363;
    wire N__98358;
    wire N__98355;
    wire N__98352;
    wire N__98351;
    wire N__98346;
    wire N__98345;
    wire N__98344;
    wire N__98343;
    wire N__98342;
    wire N__98339;
    wire N__98336;
    wire N__98335;
    wire N__98330;
    wire N__98327;
    wire N__98322;
    wire N__98319;
    wire N__98314;
    wire N__98311;
    wire N__98308;
    wire N__98305;
    wire N__98298;
    wire N__98295;
    wire N__98292;
    wire N__98291;
    wire N__98288;
    wire N__98285;
    wire N__98280;
    wire N__98277;
    wire N__98276;
    wire N__98275;
    wire N__98274;
    wire N__98273;
    wire N__98268;
    wire N__98265;
    wire N__98262;
    wire N__98261;
    wire N__98258;
    wire N__98253;
    wire N__98248;
    wire N__98247;
    wire N__98244;
    wire N__98243;
    wire N__98238;
    wire N__98235;
    wire N__98232;
    wire N__98229;
    wire N__98222;
    wire N__98217;
    wire N__98214;
    wire N__98211;
    wire N__98208;
    wire N__98205;
    wire N__98202;
    wire N__98199;
    wire N__98196;
    wire N__98193;
    wire N__98190;
    wire N__98187;
    wire N__98184;
    wire N__98183;
    wire N__98180;
    wire N__98177;
    wire N__98172;
    wire N__98169;
    wire N__98168;
    wire N__98165;
    wire N__98162;
    wire N__98159;
    wire N__98158;
    wire N__98155;
    wire N__98152;
    wire N__98149;
    wire N__98144;
    wire N__98141;
    wire N__98136;
    wire N__98133;
    wire N__98132;
    wire N__98129;
    wire N__98126;
    wire N__98121;
    wire N__98120;
    wire N__98119;
    wire N__98118;
    wire N__98117;
    wire N__98112;
    wire N__98111;
    wire N__98110;
    wire N__98105;
    wire N__98102;
    wire N__98099;
    wire N__98096;
    wire N__98093;
    wire N__98088;
    wire N__98087;
    wire N__98084;
    wire N__98081;
    wire N__98076;
    wire N__98073;
    wire N__98064;
    wire N__98061;
    wire N__98058;
    wire N__98055;
    wire N__98052;
    wire N__98049;
    wire N__98046;
    wire N__98043;
    wire N__98042;
    wire N__98039;
    wire N__98038;
    wire N__98035;
    wire N__98034;
    wire N__98033;
    wire N__98030;
    wire N__98027;
    wire N__98026;
    wire N__98023;
    wire N__98020;
    wire N__98017;
    wire N__98014;
    wire N__98009;
    wire N__98006;
    wire N__98003;
    wire N__98000;
    wire N__97995;
    wire N__97992;
    wire N__97987;
    wire N__97980;
    wire N__97977;
    wire N__97976;
    wire N__97975;
    wire N__97974;
    wire N__97971;
    wire N__97968;
    wire N__97963;
    wire N__97962;
    wire N__97961;
    wire N__97958;
    wire N__97955;
    wire N__97952;
    wire N__97951;
    wire N__97948;
    wire N__97945;
    wire N__97942;
    wire N__97937;
    wire N__97932;
    wire N__97929;
    wire N__97926;
    wire N__97923;
    wire N__97914;
    wire N__97911;
    wire N__97908;
    wire N__97905;
    wire N__97902;
    wire N__97901;
    wire N__97900;
    wire N__97897;
    wire N__97892;
    wire N__97887;
    wire N__97884;
    wire N__97881;
    wire N__97880;
    wire N__97877;
    wire N__97876;
    wire N__97875;
    wire N__97874;
    wire N__97871;
    wire N__97868;
    wire N__97865;
    wire N__97858;
    wire N__97853;
    wire N__97850;
    wire N__97845;
    wire N__97844;
    wire N__97843;
    wire N__97840;
    wire N__97835;
    wire N__97832;
    wire N__97827;
    wire N__97824;
    wire N__97821;
    wire N__97818;
    wire N__97815;
    wire N__97812;
    wire N__97809;
    wire N__97806;
    wire N__97805;
    wire N__97804;
    wire N__97803;
    wire N__97802;
    wire N__97801;
    wire N__97798;
    wire N__97797;
    wire N__97796;
    wire N__97795;
    wire N__97794;
    wire N__97793;
    wire N__97792;
    wire N__97791;
    wire N__97790;
    wire N__97789;
    wire N__97788;
    wire N__97787;
    wire N__97786;
    wire N__97785;
    wire N__97784;
    wire N__97783;
    wire N__97782;
    wire N__97781;
    wire N__97780;
    wire N__97779;
    wire N__97778;
    wire N__97777;
    wire N__97776;
    wire N__97775;
    wire N__97774;
    wire N__97773;
    wire N__97772;
    wire N__97771;
    wire N__97770;
    wire N__97769;
    wire N__97768;
    wire N__97767;
    wire N__97766;
    wire N__97765;
    wire N__97764;
    wire N__97763;
    wire N__97762;
    wire N__97761;
    wire N__97760;
    wire N__97759;
    wire N__97758;
    wire N__97757;
    wire N__97756;
    wire N__97755;
    wire N__97754;
    wire N__97753;
    wire N__97752;
    wire N__97751;
    wire N__97750;
    wire N__97749;
    wire N__97748;
    wire N__97747;
    wire N__97746;
    wire N__97745;
    wire N__97744;
    wire N__97743;
    wire N__97742;
    wire N__97741;
    wire N__97740;
    wire N__97739;
    wire N__97738;
    wire N__97737;
    wire N__97736;
    wire N__97735;
    wire N__97734;
    wire N__97733;
    wire N__97732;
    wire N__97731;
    wire N__97730;
    wire N__97729;
    wire N__97728;
    wire N__97727;
    wire N__97726;
    wire N__97725;
    wire N__97724;
    wire N__97723;
    wire N__97722;
    wire N__97721;
    wire N__97720;
    wire N__97719;
    wire N__97718;
    wire N__97717;
    wire N__97716;
    wire N__97715;
    wire N__97714;
    wire N__97713;
    wire N__97712;
    wire N__97711;
    wire N__97710;
    wire N__97709;
    wire N__97708;
    wire N__97707;
    wire N__97706;
    wire N__97705;
    wire N__97704;
    wire N__97703;
    wire N__97702;
    wire N__97701;
    wire N__97700;
    wire N__97699;
    wire N__97698;
    wire N__97697;
    wire N__97696;
    wire N__97695;
    wire N__97694;
    wire N__97693;
    wire N__97692;
    wire N__97691;
    wire N__97690;
    wire N__97689;
    wire N__97688;
    wire N__97687;
    wire N__97686;
    wire N__97685;
    wire N__97684;
    wire N__97683;
    wire N__97682;
    wire N__97681;
    wire N__97680;
    wire N__97679;
    wire N__97678;
    wire N__97677;
    wire N__97676;
    wire N__97675;
    wire N__97674;
    wire N__97673;
    wire N__97672;
    wire N__97671;
    wire N__97670;
    wire N__97669;
    wire N__97668;
    wire N__97667;
    wire N__97666;
    wire N__97665;
    wire N__97664;
    wire N__97663;
    wire N__97662;
    wire N__97661;
    wire N__97660;
    wire N__97659;
    wire N__97658;
    wire N__97657;
    wire N__97656;
    wire N__97655;
    wire N__97654;
    wire N__97653;
    wire N__97652;
    wire N__97651;
    wire N__97650;
    wire N__97649;
    wire N__97648;
    wire N__97647;
    wire N__97646;
    wire N__97645;
    wire N__97644;
    wire N__97643;
    wire N__97642;
    wire N__97641;
    wire N__97640;
    wire N__97639;
    wire N__97638;
    wire N__97637;
    wire N__97636;
    wire N__97635;
    wire N__97634;
    wire N__97633;
    wire N__97632;
    wire N__97631;
    wire N__97630;
    wire N__97629;
    wire N__97628;
    wire N__97627;
    wire N__97626;
    wire N__97625;
    wire N__97624;
    wire N__97623;
    wire N__97622;
    wire N__97621;
    wire N__97620;
    wire N__97619;
    wire N__97618;
    wire N__97617;
    wire N__97616;
    wire N__97615;
    wire N__97614;
    wire N__97613;
    wire N__97612;
    wire N__97611;
    wire N__97610;
    wire N__97609;
    wire N__97608;
    wire N__97607;
    wire N__97606;
    wire N__97605;
    wire N__97604;
    wire N__97603;
    wire N__97602;
    wire N__97601;
    wire N__97600;
    wire N__97599;
    wire N__97598;
    wire N__97597;
    wire N__97596;
    wire N__97595;
    wire N__97594;
    wire N__97593;
    wire N__97592;
    wire N__97591;
    wire N__97590;
    wire N__97589;
    wire N__97588;
    wire N__97587;
    wire N__97586;
    wire N__97585;
    wire N__97584;
    wire N__97583;
    wire N__97582;
    wire N__97581;
    wire N__97580;
    wire N__97579;
    wire N__97578;
    wire N__97577;
    wire N__97576;
    wire N__97575;
    wire N__97574;
    wire N__97573;
    wire N__97572;
    wire N__97571;
    wire N__97570;
    wire N__97569;
    wire N__97568;
    wire N__97567;
    wire N__97566;
    wire N__97565;
    wire N__97564;
    wire N__97563;
    wire N__97562;
    wire N__97561;
    wire N__97560;
    wire N__97559;
    wire N__97558;
    wire N__97557;
    wire N__97556;
    wire N__97555;
    wire N__97554;
    wire N__97553;
    wire N__97552;
    wire N__97551;
    wire N__97550;
    wire N__97549;
    wire N__97548;
    wire N__97547;
    wire N__97546;
    wire N__97545;
    wire N__97544;
    wire N__97543;
    wire N__97542;
    wire N__97541;
    wire N__97540;
    wire N__97539;
    wire N__97538;
    wire N__97537;
    wire N__97002;
    wire N__96999;
    wire N__96998;
    wire N__96997;
    wire N__96996;
    wire N__96995;
    wire N__96992;
    wire N__96989;
    wire N__96988;
    wire N__96985;
    wire N__96982;
    wire N__96979;
    wire N__96976;
    wire N__96973;
    wire N__96970;
    wire N__96969;
    wire N__96966;
    wire N__96961;
    wire N__96958;
    wire N__96953;
    wire N__96950;
    wire N__96949;
    wire N__96948;
    wire N__96945;
    wire N__96936;
    wire N__96933;
    wire N__96930;
    wire N__96929;
    wire N__96924;
    wire N__96921;
    wire N__96918;
    wire N__96915;
    wire N__96914;
    wire N__96911;
    wire N__96908;
    wire N__96905;
    wire N__96902;
    wire N__96899;
    wire N__96894;
    wire N__96887;
    wire N__96882;
    wire N__96881;
    wire N__96878;
    wire N__96875;
    wire N__96870;
    wire N__96867;
    wire N__96864;
    wire N__96863;
    wire N__96860;
    wire N__96857;
    wire N__96854;
    wire N__96851;
    wire N__96848;
    wire N__96843;
    wire N__96840;
    wire N__96837;
    wire N__96834;
    wire N__96833;
    wire N__96830;
    wire N__96827;
    wire N__96822;
    wire N__96819;
    wire N__96818;
    wire N__96815;
    wire N__96812;
    wire N__96811;
    wire N__96810;
    wire N__96809;
    wire N__96806;
    wire N__96803;
    wire N__96800;
    wire N__96797;
    wire N__96794;
    wire N__96783;
    wire N__96780;
    wire N__96777;
    wire N__96776;
    wire N__96773;
    wire N__96770;
    wire N__96765;
    wire N__96762;
    wire N__96759;
    wire N__96758;
    wire N__96755;
    wire N__96752;
    wire N__96749;
    wire N__96746;
    wire N__96741;
    wire N__96738;
    wire N__96735;
    wire N__96734;
    wire N__96733;
    wire N__96730;
    wire N__96729;
    wire N__96726;
    wire N__96725;
    wire N__96722;
    wire N__96719;
    wire N__96716;
    wire N__96713;
    wire N__96708;
    wire N__96699;
    wire N__96698;
    wire N__96695;
    wire N__96692;
    wire N__96689;
    wire N__96688;
    wire N__96683;
    wire N__96680;
    wire N__96675;
    wire N__96674;
    wire N__96671;
    wire N__96668;
    wire N__96663;
    wire N__96660;
    wire N__96657;
    wire N__96654;
    wire N__96651;
    wire N__96648;
    wire N__96645;
    wire N__96642;
    wire N__96639;
    wire N__96638;
    wire N__96635;
    wire N__96634;
    wire N__96631;
    wire N__96630;
    wire N__96627;
    wire N__96626;
    wire N__96623;
    wire N__96620;
    wire N__96617;
    wire N__96614;
    wire N__96611;
    wire N__96608;
    wire N__96605;
    wire N__96602;
    wire N__96601;
    wire N__96596;
    wire N__96593;
    wire N__96588;
    wire N__96585;
    wire N__96582;
    wire N__96577;
    wire N__96570;
    wire N__96567;
    wire N__96564;
    wire N__96561;
    wire N__96558;
    wire N__96555;
    wire N__96552;
    wire N__96549;
    wire N__96546;
    wire N__96543;
    wire N__96540;
    wire N__96537;
    wire N__96534;
    wire N__96531;
    wire N__96530;
    wire N__96527;
    wire N__96522;
    wire N__96519;
    wire N__96516;
    wire N__96513;
    wire N__96512;
    wire N__96511;
    wire N__96510;
    wire N__96507;
    wire N__96502;
    wire N__96499;
    wire N__96496;
    wire N__96493;
    wire N__96492;
    wire N__96491;
    wire N__96488;
    wire N__96485;
    wire N__96482;
    wire N__96479;
    wire N__96476;
    wire N__96473;
    wire N__96466;
    wire N__96459;
    wire N__96458;
    wire N__96455;
    wire N__96452;
    wire N__96451;
    wire N__96448;
    wire N__96445;
    wire N__96442;
    wire N__96437;
    wire N__96434;
    wire N__96431;
    wire N__96426;
    wire N__96423;
    wire N__96420;
    wire N__96419;
    wire N__96418;
    wire N__96417;
    wire N__96416;
    wire N__96411;
    wire N__96408;
    wire N__96405;
    wire N__96402;
    wire N__96397;
    wire N__96390;
    wire N__96387;
    wire N__96386;
    wire N__96385;
    wire N__96378;
    wire N__96375;
    wire N__96372;
    wire N__96371;
    wire N__96368;
    wire N__96365;
    wire N__96362;
    wire N__96357;
    wire N__96356;
    wire N__96351;
    wire N__96350;
    wire N__96349;
    wire N__96346;
    wire N__96343;
    wire N__96340;
    wire N__96333;
    wire N__96332;
    wire N__96329;
    wire N__96328;
    wire N__96325;
    wire N__96322;
    wire N__96319;
    wire N__96312;
    wire N__96309;
    wire N__96306;
    wire N__96303;
    wire N__96300;
    wire N__96299;
    wire N__96298;
    wire N__96297;
    wire N__96296;
    wire N__96293;
    wire N__96288;
    wire N__96285;
    wire N__96282;
    wire N__96279;
    wire N__96274;
    wire N__96271;
    wire N__96270;
    wire N__96265;
    wire N__96262;
    wire N__96259;
    wire N__96256;
    wire N__96249;
    wire N__96246;
    wire N__96243;
    wire N__96242;
    wire N__96241;
    wire N__96240;
    wire N__96239;
    wire N__96236;
    wire N__96227;
    wire N__96222;
    wire N__96219;
    wire N__96218;
    wire N__96217;
    wire N__96214;
    wire N__96209;
    wire N__96204;
    wire N__96201;
    wire N__96198;
    wire N__96195;
    wire N__96192;
    wire N__96189;
    wire N__96186;
    wire N__96183;
    wire N__96182;
    wire N__96181;
    wire N__96180;
    wire N__96179;
    wire N__96178;
    wire N__96177;
    wire N__96176;
    wire N__96175;
    wire N__96174;
    wire N__96171;
    wire N__96170;
    wire N__96169;
    wire N__96168;
    wire N__96167;
    wire N__96164;
    wire N__96161;
    wire N__96160;
    wire N__96159;
    wire N__96156;
    wire N__96155;
    wire N__96152;
    wire N__96149;
    wire N__96146;
    wire N__96145;
    wire N__96142;
    wire N__96139;
    wire N__96136;
    wire N__96135;
    wire N__96132;
    wire N__96127;
    wire N__96124;
    wire N__96123;
    wire N__96122;
    wire N__96121;
    wire N__96120;
    wire N__96119;
    wire N__96118;
    wire N__96115;
    wire N__96114;
    wire N__96113;
    wire N__96112;
    wire N__96111;
    wire N__96110;
    wire N__96109;
    wire N__96108;
    wire N__96107;
    wire N__96104;
    wire N__96101;
    wire N__96096;
    wire N__96093;
    wire N__96090;
    wire N__96087;
    wire N__96084;
    wire N__96081;
    wire N__96078;
    wire N__96075;
    wire N__96072;
    wire N__96069;
    wire N__96068;
    wire N__96067;
    wire N__96064;
    wire N__96059;
    wire N__96056;
    wire N__96055;
    wire N__96052;
    wire N__96049;
    wire N__96044;
    wire N__96039;
    wire N__96036;
    wire N__96033;
    wire N__96030;
    wire N__96027;
    wire N__96022;
    wire N__96021;
    wire N__96020;
    wire N__96017;
    wire N__96016;
    wire N__96015;
    wire N__96014;
    wire N__96011;
    wire N__96008;
    wire N__95999;
    wire N__95990;
    wire N__95989;
    wire N__95986;
    wire N__95979;
    wire N__95976;
    wire N__95973;
    wire N__95970;
    wire N__95967;
    wire N__95966;
    wire N__95963;
    wire N__95958;
    wire N__95951;
    wire N__95940;
    wire N__95935;
    wire N__95930;
    wire N__95927;
    wire N__95924;
    wire N__95919;
    wire N__95914;
    wire N__95913;
    wire N__95912;
    wire N__95909;
    wire N__95904;
    wire N__95899;
    wire N__95896;
    wire N__95893;
    wire N__95890;
    wire N__95883;
    wire N__95880;
    wire N__95867;
    wire N__95864;
    wire N__95861;
    wire N__95856;
    wire N__95845;
    wire N__95840;
    wire N__95829;
    wire N__95826;
    wire N__95823;
    wire N__95820;
    wire N__95817;
    wire N__95814;
    wire N__95811;
    wire N__95808;
    wire N__95805;
    wire N__95802;
    wire N__95799;
    wire N__95796;
    wire N__95795;
    wire N__95792;
    wire N__95791;
    wire N__95790;
    wire N__95789;
    wire N__95786;
    wire N__95783;
    wire N__95780;
    wire N__95777;
    wire N__95776;
    wire N__95773;
    wire N__95772;
    wire N__95769;
    wire N__95766;
    wire N__95763;
    wire N__95762;
    wire N__95759;
    wire N__95756;
    wire N__95753;
    wire N__95750;
    wire N__95747;
    wire N__95742;
    wire N__95741;
    wire N__95738;
    wire N__95735;
    wire N__95734;
    wire N__95733;
    wire N__95732;
    wire N__95729;
    wire N__95720;
    wire N__95717;
    wire N__95714;
    wire N__95711;
    wire N__95708;
    wire N__95705;
    wire N__95702;
    wire N__95699;
    wire N__95694;
    wire N__95689;
    wire N__95676;
    wire N__95673;
    wire N__95670;
    wire N__95667;
    wire N__95666;
    wire N__95663;
    wire N__95660;
    wire N__95657;
    wire N__95652;
    wire N__95649;
    wire N__95646;
    wire N__95643;
    wire N__95642;
    wire N__95639;
    wire N__95636;
    wire N__95633;
    wire N__95630;
    wire N__95625;
    wire N__95622;
    wire N__95621;
    wire N__95620;
    wire N__95617;
    wire N__95614;
    wire N__95611;
    wire N__95608;
    wire N__95601;
    wire N__95598;
    wire N__95595;
    wire N__95592;
    wire N__95589;
    wire N__95586;
    wire N__95583;
    wire N__95580;
    wire N__95577;
    wire N__95576;
    wire N__95573;
    wire N__95570;
    wire N__95565;
    wire N__95562;
    wire N__95559;
    wire N__95556;
    wire N__95553;
    wire N__95550;
    wire N__95547;
    wire N__95544;
    wire N__95543;
    wire N__95538;
    wire N__95535;
    wire N__95532;
    wire N__95529;
    wire N__95528;
    wire N__95527;
    wire N__95524;
    wire N__95521;
    wire N__95518;
    wire N__95511;
    wire N__95508;
    wire N__95507;
    wire N__95506;
    wire N__95503;
    wire N__95500;
    wire N__95497;
    wire N__95490;
    wire N__95487;
    wire N__95486;
    wire N__95483;
    wire N__95480;
    wire N__95475;
    wire N__95474;
    wire N__95473;
    wire N__95470;
    wire N__95467;
    wire N__95464;
    wire N__95457;
    wire N__95454;
    wire N__95453;
    wire N__95452;
    wire N__95449;
    wire N__95446;
    wire N__95443;
    wire N__95436;
    wire N__95433;
    wire N__95432;
    wire N__95431;
    wire N__95428;
    wire N__95425;
    wire N__95422;
    wire N__95415;
    wire N__95412;
    wire N__95411;
    wire N__95410;
    wire N__95407;
    wire N__95404;
    wire N__95401;
    wire N__95394;
    wire N__95391;
    wire N__95390;
    wire N__95389;
    wire N__95386;
    wire N__95383;
    wire N__95380;
    wire N__95373;
    wire N__95370;
    wire N__95367;
    wire N__95366;
    wire N__95365;
    wire N__95362;
    wire N__95359;
    wire N__95356;
    wire N__95349;
    wire N__95346;
    wire N__95345;
    wire N__95344;
    wire N__95341;
    wire N__95338;
    wire N__95335;
    wire N__95332;
    wire N__95325;
    wire N__95322;
    wire N__95321;
    wire N__95320;
    wire N__95317;
    wire N__95314;
    wire N__95311;
    wire N__95308;
    wire N__95307;
    wire N__95304;
    wire N__95299;
    wire N__95296;
    wire N__95293;
    wire N__95290;
    wire N__95283;
    wire N__95280;
    wire N__95277;
    wire N__95274;
    wire N__95271;
    wire N__95268;
    wire N__95265;
    wire N__95262;
    wire N__95259;
    wire N__95256;
    wire N__95253;
    wire N__95250;
    wire N__95247;
    wire N__95246;
    wire N__95243;
    wire N__95240;
    wire N__95239;
    wire N__95236;
    wire N__95233;
    wire N__95230;
    wire N__95223;
    wire N__95222;
    wire N__95221;
    wire N__95218;
    wire N__95215;
    wire N__95212;
    wire N__95209;
    wire N__95206;
    wire N__95203;
    wire N__95202;
    wire N__95199;
    wire N__95196;
    wire N__95193;
    wire N__95190;
    wire N__95185;
    wire N__95182;
    wire N__95175;
    wire N__95174;
    wire N__95171;
    wire N__95168;
    wire N__95163;
    wire N__95160;
    wire N__95157;
    wire N__95154;
    wire N__95151;
    wire N__95148;
    wire N__95145;
    wire N__95142;
    wire N__95141;
    wire N__95140;
    wire N__95137;
    wire N__95132;
    wire N__95127;
    wire N__95124;
    wire N__95123;
    wire N__95122;
    wire N__95119;
    wire N__95114;
    wire N__95109;
    wire N__95106;
    wire N__95103;
    wire N__95100;
    wire N__95097;
    wire N__95094;
    wire N__95091;
    wire N__95090;
    wire N__95089;
    wire N__95086;
    wire N__95081;
    wire N__95076;
    wire N__95073;
    wire N__95070;
    wire N__95069;
    wire N__95066;
    wire N__95065;
    wire N__95060;
    wire N__95057;
    wire N__95052;
    wire N__95051;
    wire N__95046;
    wire N__95043;
    wire N__95040;
    wire N__95037;
    wire N__95034;
    wire N__95033;
    wire N__95030;
    wire N__95027;
    wire N__95022;
    wire N__95019;
    wire N__95016;
    wire N__95013;
    wire N__95010;
    wire N__95009;
    wire N__95008;
    wire N__95007;
    wire N__95004;
    wire N__94999;
    wire N__94996;
    wire N__94993;
    wire N__94990;
    wire N__94987;
    wire N__94984;
    wire N__94983;
    wire N__94982;
    wire N__94979;
    wire N__94974;
    wire N__94969;
    wire N__94962;
    wire N__94959;
    wire N__94956;
    wire N__94955;
    wire N__94952;
    wire N__94949;
    wire N__94946;
    wire N__94941;
    wire N__94938;
    wire N__94935;
    wire N__94932;
    wire N__94929;
    wire N__94928;
    wire N__94925;
    wire N__94924;
    wire N__94921;
    wire N__94918;
    wire N__94915;
    wire N__94910;
    wire N__94909;
    wire N__94904;
    wire N__94901;
    wire N__94898;
    wire N__94893;
    wire N__94890;
    wire N__94889;
    wire N__94886;
    wire N__94883;
    wire N__94882;
    wire N__94877;
    wire N__94874;
    wire N__94871;
    wire N__94866;
    wire N__94863;
    wire N__94862;
    wire N__94859;
    wire N__94856;
    wire N__94855;
    wire N__94852;
    wire N__94849;
    wire N__94846;
    wire N__94843;
    wire N__94836;
    wire N__94835;
    wire N__94834;
    wire N__94833;
    wire N__94832;
    wire N__94831;
    wire N__94826;
    wire N__94825;
    wire N__94822;
    wire N__94821;
    wire N__94818;
    wire N__94817;
    wire N__94816;
    wire N__94815;
    wire N__94814;
    wire N__94811;
    wire N__94808;
    wire N__94805;
    wire N__94804;
    wire N__94803;
    wire N__94802;
    wire N__94801;
    wire N__94800;
    wire N__94797;
    wire N__94796;
    wire N__94793;
    wire N__94790;
    wire N__94787;
    wire N__94786;
    wire N__94785;
    wire N__94784;
    wire N__94783;
    wire N__94782;
    wire N__94781;
    wire N__94780;
    wire N__94775;
    wire N__94770;
    wire N__94763;
    wire N__94754;
    wire N__94751;
    wire N__94750;
    wire N__94749;
    wire N__94748;
    wire N__94747;
    wire N__94744;
    wire N__94741;
    wire N__94738;
    wire N__94735;
    wire N__94732;
    wire N__94727;
    wire N__94724;
    wire N__94715;
    wire N__94706;
    wire N__94703;
    wire N__94700;
    wire N__94699;
    wire N__94694;
    wire N__94691;
    wire N__94690;
    wire N__94689;
    wire N__94684;
    wire N__94681;
    wire N__94678;
    wire N__94675;
    wire N__94666;
    wire N__94663;
    wire N__94660;
    wire N__94657;
    wire N__94654;
    wire N__94651;
    wire N__94648;
    wire N__94645;
    wire N__94640;
    wire N__94633;
    wire N__94630;
    wire N__94627;
    wire N__94624;
    wire N__94621;
    wire N__94618;
    wire N__94609;
    wire N__94604;
    wire N__94601;
    wire N__94592;
    wire N__94587;
    wire N__94584;
    wire N__94581;
    wire N__94578;
    wire N__94577;
    wire N__94576;
    wire N__94575;
    wire N__94574;
    wire N__94573;
    wire N__94572;
    wire N__94569;
    wire N__94564;
    wire N__94561;
    wire N__94556;
    wire N__94551;
    wire N__94542;
    wire N__94539;
    wire N__94536;
    wire N__94535;
    wire N__94534;
    wire N__94533;
    wire N__94528;
    wire N__94527;
    wire N__94524;
    wire N__94521;
    wire N__94518;
    wire N__94515;
    wire N__94514;
    wire N__94513;
    wire N__94510;
    wire N__94507;
    wire N__94504;
    wire N__94501;
    wire N__94498;
    wire N__94495;
    wire N__94490;
    wire N__94485;
    wire N__94482;
    wire N__94473;
    wire N__94472;
    wire N__94469;
    wire N__94464;
    wire N__94463;
    wire N__94460;
    wire N__94457;
    wire N__94454;
    wire N__94449;
    wire N__94446;
    wire N__94443;
    wire N__94440;
    wire N__94437;
    wire N__94434;
    wire N__94431;
    wire N__94428;
    wire N__94425;
    wire N__94422;
    wire N__94421;
    wire N__94420;
    wire N__94417;
    wire N__94414;
    wire N__94411;
    wire N__94408;
    wire N__94405;
    wire N__94402;
    wire N__94399;
    wire N__94396;
    wire N__94389;
    wire N__94388;
    wire N__94385;
    wire N__94382;
    wire N__94379;
    wire N__94374;
    wire N__94371;
    wire N__94370;
    wire N__94367;
    wire N__94364;
    wire N__94363;
    wire N__94362;
    wire N__94359;
    wire N__94356;
    wire N__94351;
    wire N__94348;
    wire N__94341;
    wire N__94338;
    wire N__94335;
    wire N__94332;
    wire N__94329;
    wire N__94326;
    wire N__94325;
    wire N__94324;
    wire N__94323;
    wire N__94318;
    wire N__94315;
    wire N__94312;
    wire N__94311;
    wire N__94310;
    wire N__94307;
    wire N__94304;
    wire N__94301;
    wire N__94296;
    wire N__94295;
    wire N__94292;
    wire N__94287;
    wire N__94284;
    wire N__94281;
    wire N__94278;
    wire N__94273;
    wire N__94266;
    wire N__94263;
    wire N__94262;
    wire N__94259;
    wire N__94256;
    wire N__94253;
    wire N__94250;
    wire N__94245;
    wire N__94242;
    wire N__94239;
    wire N__94236;
    wire N__94235;
    wire N__94232;
    wire N__94229;
    wire N__94224;
    wire N__94221;
    wire N__94218;
    wire N__94215;
    wire N__94212;
    wire N__94209;
    wire N__94206;
    wire N__94203;
    wire N__94200;
    wire N__94197;
    wire N__94194;
    wire N__94191;
    wire N__94190;
    wire N__94187;
    wire N__94184;
    wire N__94181;
    wire N__94178;
    wire N__94177;
    wire N__94174;
    wire N__94171;
    wire N__94168;
    wire N__94165;
    wire N__94158;
    wire N__94155;
    wire N__94152;
    wire N__94151;
    wire N__94148;
    wire N__94145;
    wire N__94144;
    wire N__94141;
    wire N__94138;
    wire N__94135;
    wire N__94132;
    wire N__94125;
    wire N__94122;
    wire N__94119;
    wire N__94116;
    wire N__94113;
    wire N__94112;
    wire N__94109;
    wire N__94106;
    wire N__94103;
    wire N__94100;
    wire N__94095;
    wire N__94094;
    wire N__94091;
    wire N__94088;
    wire N__94083;
    wire N__94080;
    wire N__94077;
    wire N__94076;
    wire N__94073;
    wire N__94070;
    wire N__94067;
    wire N__94064;
    wire N__94059;
    wire N__94056;
    wire N__94053;
    wire N__94050;
    wire N__94047;
    wire N__94044;
    wire N__94041;
    wire N__94038;
    wire N__94035;
    wire N__94034;
    wire N__94031;
    wire N__94028;
    wire N__94023;
    wire N__94022;
    wire N__94021;
    wire N__94016;
    wire N__94015;
    wire N__94012;
    wire N__94009;
    wire N__94004;
    wire N__93999;
    wire N__93996;
    wire N__93993;
    wire N__93992;
    wire N__93989;
    wire N__93988;
    wire N__93985;
    wire N__93982;
    wire N__93977;
    wire N__93972;
    wire N__93969;
    wire N__93966;
    wire N__93963;
    wire N__93960;
    wire N__93957;
    wire N__93956;
    wire N__93953;
    wire N__93950;
    wire N__93945;
    wire N__93944;
    wire N__93941;
    wire N__93938;
    wire N__93933;
    wire N__93932;
    wire N__93929;
    wire N__93926;
    wire N__93921;
    wire N__93920;
    wire N__93917;
    wire N__93914;
    wire N__93909;
    wire N__93906;
    wire N__93903;
    wire N__93900;
    wire N__93897;
    wire N__93894;
    wire N__93891;
    wire N__93888;
    wire N__93885;
    wire N__93882;
    wire N__93879;
    wire N__93876;
    wire N__93873;
    wire N__93870;
    wire N__93867;
    wire N__93864;
    wire N__93861;
    wire N__93858;
    wire N__93855;
    wire N__93852;
    wire N__93849;
    wire N__93846;
    wire N__93843;
    wire N__93840;
    wire N__93837;
    wire N__93834;
    wire N__93831;
    wire N__93830;
    wire N__93827;
    wire N__93824;
    wire N__93821;
    wire N__93818;
    wire N__93815;
    wire N__93810;
    wire N__93807;
    wire N__93804;
    wire N__93803;
    wire N__93800;
    wire N__93797;
    wire N__93794;
    wire N__93791;
    wire N__93788;
    wire N__93783;
    wire N__93782;
    wire N__93779;
    wire N__93776;
    wire N__93775;
    wire N__93770;
    wire N__93767;
    wire N__93762;
    wire N__93759;
    wire N__93756;
    wire N__93755;
    wire N__93752;
    wire N__93749;
    wire N__93748;
    wire N__93743;
    wire N__93740;
    wire N__93735;
    wire N__93732;
    wire N__93729;
    wire N__93728;
    wire N__93725;
    wire N__93722;
    wire N__93721;
    wire N__93716;
    wire N__93713;
    wire N__93708;
    wire N__93705;
    wire N__93702;
    wire N__93701;
    wire N__93700;
    wire N__93699;
    wire N__93698;
    wire N__93697;
    wire N__93694;
    wire N__93691;
    wire N__93688;
    wire N__93685;
    wire N__93682;
    wire N__93679;
    wire N__93674;
    wire N__93665;
    wire N__93660;
    wire N__93657;
    wire N__93656;
    wire N__93653;
    wire N__93650;
    wire N__93649;
    wire N__93646;
    wire N__93643;
    wire N__93640;
    wire N__93635;
    wire N__93632;
    wire N__93627;
    wire N__93624;
    wire N__93621;
    wire N__93620;
    wire N__93619;
    wire N__93616;
    wire N__93613;
    wire N__93610;
    wire N__93603;
    wire N__93600;
    wire N__93597;
    wire N__93594;
    wire N__93591;
    wire N__93590;
    wire N__93589;
    wire N__93586;
    wire N__93583;
    wire N__93580;
    wire N__93573;
    wire N__93570;
    wire N__93567;
    wire N__93564;
    wire N__93563;
    wire N__93562;
    wire N__93559;
    wire N__93556;
    wire N__93553;
    wire N__93552;
    wire N__93551;
    wire N__93548;
    wire N__93543;
    wire N__93540;
    wire N__93537;
    wire N__93532;
    wire N__93527;
    wire N__93522;
    wire N__93519;
    wire N__93516;
    wire N__93513;
    wire N__93510;
    wire N__93507;
    wire N__93504;
    wire N__93503;
    wire N__93502;
    wire N__93499;
    wire N__93496;
    wire N__93493;
    wire N__93486;
    wire N__93485;
    wire N__93482;
    wire N__93479;
    wire N__93476;
    wire N__93471;
    wire N__93470;
    wire N__93467;
    wire N__93464;
    wire N__93463;
    wire N__93458;
    wire N__93455;
    wire N__93452;
    wire N__93449;
    wire N__93444;
    wire N__93441;
    wire N__93440;
    wire N__93439;
    wire N__93436;
    wire N__93433;
    wire N__93430;
    wire N__93425;
    wire N__93422;
    wire N__93419;
    wire N__93416;
    wire N__93411;
    wire N__93408;
    wire N__93407;
    wire N__93404;
    wire N__93401;
    wire N__93400;
    wire N__93395;
    wire N__93392;
    wire N__93387;
    wire N__93384;
    wire N__93381;
    wire N__93380;
    wire N__93379;
    wire N__93376;
    wire N__93373;
    wire N__93370;
    wire N__93369;
    wire N__93364;
    wire N__93361;
    wire N__93358;
    wire N__93355;
    wire N__93352;
    wire N__93345;
    wire N__93342;
    wire N__93341;
    wire N__93340;
    wire N__93337;
    wire N__93334;
    wire N__93331;
    wire N__93330;
    wire N__93325;
    wire N__93322;
    wire N__93319;
    wire N__93316;
    wire N__93313;
    wire N__93306;
    wire N__93305;
    wire N__93304;
    wire N__93303;
    wire N__93302;
    wire N__93301;
    wire N__93298;
    wire N__93295;
    wire N__93292;
    wire N__93289;
    wire N__93286;
    wire N__93283;
    wire N__93278;
    wire N__93269;
    wire N__93264;
    wire N__93261;
    wire N__93258;
    wire N__93255;
    wire N__93252;
    wire N__93249;
    wire N__93246;
    wire N__93243;
    wire N__93240;
    wire N__93237;
    wire N__93234;
    wire N__93231;
    wire N__93228;
    wire N__93227;
    wire N__93226;
    wire N__93225;
    wire N__93224;
    wire N__93223;
    wire N__93220;
    wire N__93219;
    wire N__93216;
    wire N__93209;
    wire N__93206;
    wire N__93203;
    wire N__93202;
    wire N__93199;
    wire N__93198;
    wire N__93195;
    wire N__93192;
    wire N__93189;
    wire N__93186;
    wire N__93185;
    wire N__93182;
    wire N__93179;
    wire N__93176;
    wire N__93171;
    wire N__93166;
    wire N__93163;
    wire N__93160;
    wire N__93155;
    wire N__93152;
    wire N__93149;
    wire N__93146;
    wire N__93143;
    wire N__93134;
    wire N__93133;
    wire N__93130;
    wire N__93127;
    wire N__93124;
    wire N__93117;
    wire N__93114;
    wire N__93111;
    wire N__93108;
    wire N__93105;
    wire N__93104;
    wire N__93103;
    wire N__93100;
    wire N__93097;
    wire N__93094;
    wire N__93093;
    wire N__93088;
    wire N__93085;
    wire N__93082;
    wire N__93079;
    wire N__93076;
    wire N__93069;
    wire N__93066;
    wire N__93065;
    wire N__93064;
    wire N__93061;
    wire N__93058;
    wire N__93055;
    wire N__93054;
    wire N__93047;
    wire N__93044;
    wire N__93041;
    wire N__93036;
    wire N__93033;
    wire N__93030;
    wire N__93027;
    wire N__93024;
    wire N__93023;
    wire N__93022;
    wire N__93019;
    wire N__93016;
    wire N__93013;
    wire N__93012;
    wire N__93007;
    wire N__93004;
    wire N__93001;
    wire N__92998;
    wire N__92995;
    wire N__92988;
    wire N__92985;
    wire N__92984;
    wire N__92983;
    wire N__92980;
    wire N__92977;
    wire N__92974;
    wire N__92973;
    wire N__92966;
    wire N__92963;
    wire N__92960;
    wire N__92955;
    wire N__92952;
    wire N__92951;
    wire N__92950;
    wire N__92947;
    wire N__92944;
    wire N__92941;
    wire N__92938;
    wire N__92937;
    wire N__92930;
    wire N__92927;
    wire N__92924;
    wire N__92919;
    wire N__92916;
    wire N__92915;
    wire N__92914;
    wire N__92911;
    wire N__92908;
    wire N__92905;
    wire N__92904;
    wire N__92903;
    wire N__92902;
    wire N__92901;
    wire N__92900;
    wire N__92899;
    wire N__92898;
    wire N__92897;
    wire N__92896;
    wire N__92895;
    wire N__92894;
    wire N__92887;
    wire N__92884;
    wire N__92881;
    wire N__92878;
    wire N__92877;
    wire N__92876;
    wire N__92875;
    wire N__92874;
    wire N__92873;
    wire N__92872;
    wire N__92871;
    wire N__92870;
    wire N__92867;
    wire N__92866;
    wire N__92865;
    wire N__92864;
    wire N__92861;
    wire N__92858;
    wire N__92855;
    wire N__92852;
    wire N__92849;
    wire N__92846;
    wire N__92845;
    wire N__92844;
    wire N__92843;
    wire N__92842;
    wire N__92841;
    wire N__92840;
    wire N__92839;
    wire N__92838;
    wire N__92837;
    wire N__92834;
    wire N__92831;
    wire N__92826;
    wire N__92823;
    wire N__92820;
    wire N__92817;
    wire N__92814;
    wire N__92811;
    wire N__92808;
    wire N__92805;
    wire N__92802;
    wire N__92799;
    wire N__92796;
    wire N__92793;
    wire N__92790;
    wire N__92787;
    wire N__92778;
    wire N__92775;
    wire N__92772;
    wire N__92769;
    wire N__92766;
    wire N__92763;
    wire N__92760;
    wire N__92757;
    wire N__92754;
    wire N__92751;
    wire N__92750;
    wire N__92747;
    wire N__92744;
    wire N__92735;
    wire N__92724;
    wire N__92707;
    wire N__92702;
    wire N__92687;
    wire N__92684;
    wire N__92681;
    wire N__92680;
    wire N__92679;
    wire N__92678;
    wire N__92675;
    wire N__92670;
    wire N__92661;
    wire N__92658;
    wire N__92655;
    wire N__92650;
    wire N__92647;
    wire N__92642;
    wire N__92637;
    wire N__92634;
    wire N__92625;
    wire N__92622;
    wire N__92619;
    wire N__92618;
    wire N__92617;
    wire N__92616;
    wire N__92615;
    wire N__92614;
    wire N__92613;
    wire N__92610;
    wire N__92607;
    wire N__92604;
    wire N__92601;
    wire N__92600;
    wire N__92599;
    wire N__92596;
    wire N__92591;
    wire N__92586;
    wire N__92583;
    wire N__92580;
    wire N__92577;
    wire N__92574;
    wire N__92571;
    wire N__92564;
    wire N__92561;
    wire N__92558;
    wire N__92555;
    wire N__92550;
    wire N__92547;
    wire N__92544;
    wire N__92541;
    wire N__92538;
    wire N__92533;
    wire N__92530;
    wire N__92525;
    wire N__92524;
    wire N__92523;
    wire N__92518;
    wire N__92513;
    wire N__92510;
    wire N__92505;
    wire N__92502;
    wire N__92499;
    wire N__92496;
    wire N__92493;
    wire N__92490;
    wire N__92489;
    wire N__92486;
    wire N__92483;
    wire N__92482;
    wire N__92479;
    wire N__92476;
    wire N__92473;
    wire N__92470;
    wire N__92463;
    wire N__92460;
    wire N__92457;
    wire N__92454;
    wire N__92451;
    wire N__92448;
    wire N__92445;
    wire N__92442;
    wire N__92439;
    wire N__92436;
    wire N__92433;
    wire N__92430;
    wire N__92427;
    wire N__92424;
    wire N__92423;
    wire N__92420;
    wire N__92417;
    wire N__92416;
    wire N__92411;
    wire N__92408;
    wire N__92405;
    wire N__92400;
    wire N__92397;
    wire N__92394;
    wire N__92391;
    wire N__92390;
    wire N__92389;
    wire N__92386;
    wire N__92383;
    wire N__92380;
    wire N__92377;
    wire N__92370;
    wire N__92367;
    wire N__92364;
    wire N__92361;
    wire N__92358;
    wire N__92355;
    wire N__92354;
    wire N__92353;
    wire N__92350;
    wire N__92347;
    wire N__92344;
    wire N__92341;
    wire N__92334;
    wire N__92331;
    wire N__92328;
    wire N__92325;
    wire N__92322;
    wire N__92319;
    wire N__92318;
    wire N__92317;
    wire N__92314;
    wire N__92311;
    wire N__92308;
    wire N__92305;
    wire N__92298;
    wire N__92295;
    wire N__92292;
    wire N__92289;
    wire N__92286;
    wire N__92283;
    wire N__92280;
    wire N__92277;
    wire N__92274;
    wire N__92273;
    wire N__92272;
    wire N__92269;
    wire N__92266;
    wire N__92263;
    wire N__92256;
    wire N__92253;
    wire N__92250;
    wire N__92247;
    wire N__92244;
    wire N__92241;
    wire N__92240;
    wire N__92239;
    wire N__92236;
    wire N__92233;
    wire N__92230;
    wire N__92227;
    wire N__92220;
    wire N__92217;
    wire N__92214;
    wire N__92211;
    wire N__92208;
    wire N__92205;
    wire N__92202;
    wire N__92199;
    wire N__92196;
    wire N__92195;
    wire N__92194;
    wire N__92191;
    wire N__92186;
    wire N__92181;
    wire N__92178;
    wire N__92175;
    wire N__92172;
    wire N__92169;
    wire N__92166;
    wire N__92163;
    wire N__92162;
    wire N__92157;
    wire N__92156;
    wire N__92153;
    wire N__92150;
    wire N__92147;
    wire N__92142;
    wire N__92139;
    wire N__92136;
    wire N__92133;
    wire N__92130;
    wire N__92127;
    wire N__92124;
    wire N__92121;
    wire N__92120;
    wire N__92119;
    wire N__92116;
    wire N__92113;
    wire N__92110;
    wire N__92107;
    wire N__92100;
    wire N__92097;
    wire N__92094;
    wire N__92093;
    wire N__92090;
    wire N__92087;
    wire N__92084;
    wire N__92081;
    wire N__92080;
    wire N__92075;
    wire N__92072;
    wire N__92069;
    wire N__92064;
    wire N__92061;
    wire N__92058;
    wire N__92055;
    wire N__92052;
    wire N__92049;
    wire N__92048;
    wire N__92045;
    wire N__92042;
    wire N__92041;
    wire N__92038;
    wire N__92035;
    wire N__92032;
    wire N__92029;
    wire N__92022;
    wire N__92019;
    wire N__92016;
    wire N__92013;
    wire N__92010;
    wire N__92009;
    wire N__92006;
    wire N__92003;
    wire N__92000;
    wire N__91999;
    wire N__91994;
    wire N__91991;
    wire N__91988;
    wire N__91983;
    wire N__91980;
    wire N__91977;
    wire N__91974;
    wire N__91971;
    wire N__91968;
    wire N__91967;
    wire N__91964;
    wire N__91961;
    wire N__91960;
    wire N__91955;
    wire N__91952;
    wire N__91949;
    wire N__91944;
    wire N__91941;
    wire N__91938;
    wire N__91935;
    wire N__91932;
    wire N__91929;
    wire N__91928;
    wire N__91925;
    wire N__91922;
    wire N__91917;
    wire N__91914;
    wire N__91913;
    wire N__91910;
    wire N__91907;
    wire N__91902;
    wire N__91899;
    wire N__91896;
    wire N__91893;
    wire N__91890;
    wire N__91887;
    wire N__91886;
    wire N__91883;
    wire N__91880;
    wire N__91879;
    wire N__91874;
    wire N__91871;
    wire N__91868;
    wire N__91863;
    wire N__91860;
    wire N__91857;
    wire N__91854;
    wire N__91851;
    wire N__91848;
    wire N__91845;
    wire N__91842;
    wire N__91841;
    wire N__91838;
    wire N__91835;
    wire N__91832;
    wire N__91829;
    wire N__91826;
    wire N__91823;
    wire N__91822;
    wire N__91819;
    wire N__91816;
    wire N__91813;
    wire N__91810;
    wire N__91803;
    wire N__91800;
    wire N__91797;
    wire N__91794;
    wire N__91791;
    wire N__91788;
    wire N__91785;
    wire N__91784;
    wire N__91779;
    wire N__91778;
    wire N__91775;
    wire N__91772;
    wire N__91769;
    wire N__91764;
    wire N__91761;
    wire N__91758;
    wire N__91755;
    wire N__91752;
    wire N__91749;
    wire N__91746;
    wire N__91743;
    wire N__91740;
    wire N__91737;
    wire N__91736;
    wire N__91735;
    wire N__91732;
    wire N__91729;
    wire N__91726;
    wire N__91723;
    wire N__91716;
    wire N__91713;
    wire N__91710;
    wire N__91709;
    wire N__91706;
    wire N__91703;
    wire N__91700;
    wire N__91697;
    wire N__91694;
    wire N__91693;
    wire N__91690;
    wire N__91687;
    wire N__91684;
    wire N__91681;
    wire N__91674;
    wire N__91671;
    wire N__91668;
    wire N__91665;
    wire N__91662;
    wire N__91659;
    wire N__91656;
    wire N__91653;
    wire N__91650;
    wire N__91649;
    wire N__91648;
    wire N__91645;
    wire N__91640;
    wire N__91639;
    wire N__91638;
    wire N__91635;
    wire N__91632;
    wire N__91629;
    wire N__91628;
    wire N__91625;
    wire N__91622;
    wire N__91619;
    wire N__91616;
    wire N__91613;
    wire N__91610;
    wire N__91607;
    wire N__91602;
    wire N__91599;
    wire N__91592;
    wire N__91591;
    wire N__91586;
    wire N__91583;
    wire N__91578;
    wire N__91575;
    wire N__91572;
    wire N__91569;
    wire N__91566;
    wire N__91563;
    wire N__91560;
    wire N__91557;
    wire N__91556;
    wire N__91555;
    wire N__91554;
    wire N__91551;
    wire N__91546;
    wire N__91543;
    wire N__91540;
    wire N__91537;
    wire N__91534;
    wire N__91529;
    wire N__91528;
    wire N__91523;
    wire N__91520;
    wire N__91519;
    wire N__91514;
    wire N__91511;
    wire N__91508;
    wire N__91505;
    wire N__91502;
    wire N__91501;
    wire N__91498;
    wire N__91495;
    wire N__91492;
    wire N__91485;
    wire N__91482;
    wire N__91479;
    wire N__91476;
    wire N__91473;
    wire N__91470;
    wire N__91469;
    wire N__91468;
    wire N__91467;
    wire N__91464;
    wire N__91457;
    wire N__91456;
    wire N__91453;
    wire N__91452;
    wire N__91449;
    wire N__91446;
    wire N__91443;
    wire N__91440;
    wire N__91439;
    wire N__91436;
    wire N__91433;
    wire N__91428;
    wire N__91425;
    wire N__91422;
    wire N__91419;
    wire N__91416;
    wire N__91409;
    wire N__91406;
    wire N__91405;
    wire N__91404;
    wire N__91399;
    wire N__91396;
    wire N__91393;
    wire N__91390;
    wire N__91383;
    wire N__91380;
    wire N__91377;
    wire N__91374;
    wire N__91371;
    wire N__91368;
    wire N__91367;
    wire N__91366;
    wire N__91365;
    wire N__91362;
    wire N__91359;
    wire N__91356;
    wire N__91353;
    wire N__91352;
    wire N__91349;
    wire N__91346;
    wire N__91339;
    wire N__91336;
    wire N__91333;
    wire N__91330;
    wire N__91329;
    wire N__91322;
    wire N__91321;
    wire N__91318;
    wire N__91315;
    wire N__91312;
    wire N__91309;
    wire N__91302;
    wire N__91299;
    wire N__91298;
    wire N__91295;
    wire N__91294;
    wire N__91291;
    wire N__91288;
    wire N__91285;
    wire N__91278;
    wire N__91275;
    wire N__91272;
    wire N__91269;
    wire N__91266;
    wire N__91263;
    wire N__91260;
    wire N__91259;
    wire N__91258;
    wire N__91255;
    wire N__91252;
    wire N__91251;
    wire N__91250;
    wire N__91247;
    wire N__91246;
    wire N__91241;
    wire N__91240;
    wire N__91239;
    wire N__91236;
    wire N__91231;
    wire N__91228;
    wire N__91225;
    wire N__91222;
    wire N__91221;
    wire N__91218;
    wire N__91215;
    wire N__91210;
    wire N__91209;
    wire N__91206;
    wire N__91203;
    wire N__91202;
    wire N__91199;
    wire N__91192;
    wire N__91189;
    wire N__91184;
    wire N__91181;
    wire N__91178;
    wire N__91175;
    wire N__91172;
    wire N__91169;
    wire N__91166;
    wire N__91159;
    wire N__91156;
    wire N__91155;
    wire N__91150;
    wire N__91147;
    wire N__91144;
    wire N__91137;
    wire N__91134;
    wire N__91131;
    wire N__91128;
    wire N__91125;
    wire N__91122;
    wire N__91119;
    wire N__91116;
    wire N__91115;
    wire N__91112;
    wire N__91111;
    wire N__91110;
    wire N__91107;
    wire N__91104;
    wire N__91103;
    wire N__91102;
    wire N__91101;
    wire N__91098;
    wire N__91097;
    wire N__91094;
    wire N__91089;
    wire N__91082;
    wire N__91079;
    wire N__91078;
    wire N__91075;
    wire N__91072;
    wire N__91071;
    wire N__91066;
    wire N__91063;
    wire N__91060;
    wire N__91057;
    wire N__91054;
    wire N__91051;
    wire N__91048;
    wire N__91045;
    wire N__91042;
    wire N__91039;
    wire N__91036;
    wire N__91033;
    wire N__91032;
    wire N__91029;
    wire N__91026;
    wire N__91023;
    wire N__91018;
    wire N__91015;
    wire N__91012;
    wire N__91009;
    wire N__91006;
    wire N__91003;
    wire N__91000;
    wire N__90997;
    wire N__90994;
    wire N__90991;
    wire N__90982;
    wire N__90981;
    wire N__90978;
    wire N__90973;
    wire N__90970;
    wire N__90963;
    wire N__90960;
    wire N__90957;
    wire N__90954;
    wire N__90951;
    wire N__90948;
    wire N__90945;
    wire N__90942;
    wire N__90941;
    wire N__90940;
    wire N__90937;
    wire N__90934;
    wire N__90931;
    wire N__90930;
    wire N__90929;
    wire N__90922;
    wire N__90917;
    wire N__90912;
    wire N__90909;
    wire N__90906;
    wire N__90903;
    wire N__90900;
    wire N__90897;
    wire N__90894;
    wire N__90891;
    wire N__90888;
    wire N__90885;
    wire N__90884;
    wire N__90881;
    wire N__90878;
    wire N__90877;
    wire N__90874;
    wire N__90873;
    wire N__90872;
    wire N__90871;
    wire N__90870;
    wire N__90867;
    wire N__90864;
    wire N__90861;
    wire N__90858;
    wire N__90855;
    wire N__90852;
    wire N__90849;
    wire N__90846;
    wire N__90843;
    wire N__90840;
    wire N__90835;
    wire N__90832;
    wire N__90829;
    wire N__90826;
    wire N__90819;
    wire N__90814;
    wire N__90807;
    wire N__90804;
    wire N__90801;
    wire N__90798;
    wire N__90795;
    wire N__90794;
    wire N__90793;
    wire N__90790;
    wire N__90789;
    wire N__90786;
    wire N__90785;
    wire N__90782;
    wire N__90779;
    wire N__90778;
    wire N__90775;
    wire N__90774;
    wire N__90771;
    wire N__90768;
    wire N__90767;
    wire N__90764;
    wire N__90761;
    wire N__90760;
    wire N__90759;
    wire N__90758;
    wire N__90755;
    wire N__90752;
    wire N__90749;
    wire N__90746;
    wire N__90743;
    wire N__90740;
    wire N__90735;
    wire N__90732;
    wire N__90729;
    wire N__90728;
    wire N__90725;
    wire N__90724;
    wire N__90721;
    wire N__90718;
    wire N__90711;
    wire N__90702;
    wire N__90699;
    wire N__90696;
    wire N__90695;
    wire N__90694;
    wire N__90693;
    wire N__90692;
    wire N__90689;
    wire N__90686;
    wire N__90683;
    wire N__90678;
    wire N__90675;
    wire N__90672;
    wire N__90669;
    wire N__90666;
    wire N__90663;
    wire N__90660;
    wire N__90657;
    wire N__90650;
    wire N__90643;
    wire N__90630;
    wire N__90627;
    wire N__90624;
    wire N__90621;
    wire N__90618;
    wire N__90615;
    wire N__90612;
    wire N__90609;
    wire N__90606;
    wire N__90603;
    wire N__90602;
    wire N__90599;
    wire N__90596;
    wire N__90591;
    wire N__90588;
    wire N__90585;
    wire N__90582;
    wire N__90579;
    wire N__90578;
    wire N__90575;
    wire N__90574;
    wire N__90573;
    wire N__90570;
    wire N__90567;
    wire N__90562;
    wire N__90559;
    wire N__90554;
    wire N__90551;
    wire N__90548;
    wire N__90543;
    wire N__90540;
    wire N__90537;
    wire N__90534;
    wire N__90531;
    wire N__90528;
    wire N__90525;
    wire N__90522;
    wire N__90519;
    wire N__90516;
    wire N__90513;
    wire N__90510;
    wire N__90507;
    wire N__90504;
    wire N__90501;
    wire N__90498;
    wire N__90497;
    wire N__90494;
    wire N__90493;
    wire N__90490;
    wire N__90487;
    wire N__90484;
    wire N__90481;
    wire N__90476;
    wire N__90473;
    wire N__90470;
    wire N__90467;
    wire N__90464;
    wire N__90461;
    wire N__90458;
    wire N__90453;
    wire N__90450;
    wire N__90449;
    wire N__90448;
    wire N__90445;
    wire N__90442;
    wire N__90439;
    wire N__90434;
    wire N__90429;
    wire N__90426;
    wire N__90423;
    wire N__90420;
    wire N__90417;
    wire N__90414;
    wire N__90411;
    wire N__90408;
    wire N__90405;
    wire N__90402;
    wire N__90399;
    wire N__90396;
    wire N__90395;
    wire N__90394;
    wire N__90393;
    wire N__90392;
    wire N__90391;
    wire N__90388;
    wire N__90387;
    wire N__90386;
    wire N__90385;
    wire N__90382;
    wire N__90381;
    wire N__90380;
    wire N__90379;
    wire N__90378;
    wire N__90377;
    wire N__90376;
    wire N__90375;
    wire N__90374;
    wire N__90373;
    wire N__90372;
    wire N__90371;
    wire N__90370;
    wire N__90367;
    wire N__90364;
    wire N__90361;
    wire N__90358;
    wire N__90355;
    wire N__90348;
    wire N__90345;
    wire N__90344;
    wire N__90343;
    wire N__90340;
    wire N__90339;
    wire N__90336;
    wire N__90335;
    wire N__90332;
    wire N__90329;
    wire N__90326;
    wire N__90323;
    wire N__90322;
    wire N__90321;
    wire N__90320;
    wire N__90319;
    wire N__90318;
    wire N__90317;
    wire N__90316;
    wire N__90315;
    wire N__90314;
    wire N__90311;
    wire N__90304;
    wire N__90301;
    wire N__90298;
    wire N__90295;
    wire N__90292;
    wire N__90289;
    wire N__90286;
    wire N__90279;
    wire N__90276;
    wire N__90273;
    wire N__90270;
    wire N__90267;
    wire N__90264;
    wire N__90259;
    wire N__90254;
    wire N__90251;
    wire N__90244;
    wire N__90239;
    wire N__90232;
    wire N__90231;
    wire N__90228;
    wire N__90225;
    wire N__90222;
    wire N__90219;
    wire N__90212;
    wire N__90209;
    wire N__90208;
    wire N__90207;
    wire N__90206;
    wire N__90201;
    wire N__90194;
    wire N__90193;
    wire N__90192;
    wire N__90183;
    wire N__90180;
    wire N__90173;
    wire N__90170;
    wire N__90167;
    wire N__90156;
    wire N__90149;
    wire N__90144;
    wire N__90141;
    wire N__90138;
    wire N__90133;
    wire N__90128;
    wire N__90123;
    wire N__90118;
    wire N__90105;
    wire N__90104;
    wire N__90103;
    wire N__90102;
    wire N__90101;
    wire N__90100;
    wire N__90097;
    wire N__90096;
    wire N__90095;
    wire N__90094;
    wire N__90093;
    wire N__90090;
    wire N__90087;
    wire N__90086;
    wire N__90085;
    wire N__90084;
    wire N__90079;
    wire N__90076;
    wire N__90075;
    wire N__90074;
    wire N__90071;
    wire N__90068;
    wire N__90065;
    wire N__90064;
    wire N__90055;
    wire N__90052;
    wire N__90051;
    wire N__90048;
    wire N__90047;
    wire N__90046;
    wire N__90045;
    wire N__90044;
    wire N__90041;
    wire N__90040;
    wire N__90039;
    wire N__90034;
    wire N__90031;
    wire N__90028;
    wire N__90027;
    wire N__90024;
    wire N__90019;
    wire N__90018;
    wire N__90017;
    wire N__90014;
    wire N__90009;
    wire N__90006;
    wire N__90005;
    wire N__90004;
    wire N__90001;
    wire N__89998;
    wire N__89995;
    wire N__89992;
    wire N__89989;
    wire N__89986;
    wire N__89983;
    wire N__89980;
    wire N__89975;
    wire N__89974;
    wire N__89971;
    wire N__89968;
    wire N__89963;
    wire N__89960;
    wire N__89957;
    wire N__89950;
    wire N__89949;
    wire N__89946;
    wire N__89943;
    wire N__89936;
    wire N__89933;
    wire N__89928;
    wire N__89921;
    wire N__89918;
    wire N__89911;
    wire N__89904;
    wire N__89901;
    wire N__89892;
    wire N__89885;
    wire N__89880;
    wire N__89871;
    wire N__89868;
    wire N__89867;
    wire N__89864;
    wire N__89861;
    wire N__89858;
    wire N__89855;
    wire N__89852;
    wire N__89847;
    wire N__89844;
    wire N__89841;
    wire N__89840;
    wire N__89837;
    wire N__89834;
    wire N__89831;
    wire N__89826;
    wire N__89825;
    wire N__89824;
    wire N__89823;
    wire N__89820;
    wire N__89819;
    wire N__89812;
    wire N__89809;
    wire N__89808;
    wire N__89807;
    wire N__89804;
    wire N__89799;
    wire N__89798;
    wire N__89797;
    wire N__89796;
    wire N__89795;
    wire N__89794;
    wire N__89791;
    wire N__89788;
    wire N__89785;
    wire N__89784;
    wire N__89781;
    wire N__89778;
    wire N__89775;
    wire N__89774;
    wire N__89773;
    wire N__89772;
    wire N__89771;
    wire N__89768;
    wire N__89765;
    wire N__89762;
    wire N__89761;
    wire N__89760;
    wire N__89759;
    wire N__89758;
    wire N__89753;
    wire N__89752;
    wire N__89749;
    wire N__89746;
    wire N__89739;
    wire N__89736;
    wire N__89735;
    wire N__89730;
    wire N__89727;
    wire N__89724;
    wire N__89721;
    wire N__89718;
    wire N__89713;
    wire N__89712;
    wire N__89707;
    wire N__89704;
    wire N__89701;
    wire N__89696;
    wire N__89693;
    wire N__89690;
    wire N__89687;
    wire N__89682;
    wire N__89679;
    wire N__89672;
    wire N__89669;
    wire N__89666;
    wire N__89663;
    wire N__89660;
    wire N__89657;
    wire N__89652;
    wire N__89645;
    wire N__89640;
    wire N__89637;
    wire N__89634;
    wire N__89629;
    wire N__89626;
    wire N__89623;
    wire N__89620;
    wire N__89617;
    wire N__89614;
    wire N__89611;
    wire N__89608;
    wire N__89605;
    wire N__89596;
    wire N__89589;
    wire N__89586;
    wire N__89583;
    wire N__89580;
    wire N__89579;
    wire N__89578;
    wire N__89577;
    wire N__89576;
    wire N__89575;
    wire N__89574;
    wire N__89573;
    wire N__89572;
    wire N__89571;
    wire N__89570;
    wire N__89569;
    wire N__89568;
    wire N__89567;
    wire N__89566;
    wire N__89565;
    wire N__89564;
    wire N__89561;
    wire N__89558;
    wire N__89555;
    wire N__89552;
    wire N__89549;
    wire N__89546;
    wire N__89543;
    wire N__89540;
    wire N__89537;
    wire N__89534;
    wire N__89531;
    wire N__89528;
    wire N__89525;
    wire N__89522;
    wire N__89519;
    wire N__89516;
    wire N__89513;
    wire N__89506;
    wire N__89497;
    wire N__89488;
    wire N__89483;
    wire N__89474;
    wire N__89467;
    wire N__89464;
    wire N__89457;
    wire N__89454;
    wire N__89453;
    wire N__89452;
    wire N__89451;
    wire N__89450;
    wire N__89449;
    wire N__89446;
    wire N__89443;
    wire N__89440;
    wire N__89437;
    wire N__89434;
    wire N__89431;
    wire N__89426;
    wire N__89417;
    wire N__89412;
    wire N__89409;
    wire N__89406;
    wire N__89403;
    wire N__89402;
    wire N__89399;
    wire N__89396;
    wire N__89395;
    wire N__89394;
    wire N__89391;
    wire N__89388;
    wire N__89385;
    wire N__89382;
    wire N__89379;
    wire N__89374;
    wire N__89367;
    wire N__89366;
    wire N__89365;
    wire N__89362;
    wire N__89359;
    wire N__89356;
    wire N__89351;
    wire N__89348;
    wire N__89343;
    wire N__89342;
    wire N__89339;
    wire N__89338;
    wire N__89335;
    wire N__89332;
    wire N__89329;
    wire N__89326;
    wire N__89319;
    wire N__89318;
    wire N__89317;
    wire N__89314;
    wire N__89311;
    wire N__89308;
    wire N__89303;
    wire N__89300;
    wire N__89295;
    wire N__89292;
    wire N__89291;
    wire N__89290;
    wire N__89287;
    wire N__89284;
    wire N__89281;
    wire N__89276;
    wire N__89273;
    wire N__89268;
    wire N__89267;
    wire N__89264;
    wire N__89263;
    wire N__89260;
    wire N__89257;
    wire N__89254;
    wire N__89251;
    wire N__89244;
    wire N__89241;
    wire N__89238;
    wire N__89235;
    wire N__89232;
    wire N__89231;
    wire N__89230;
    wire N__89227;
    wire N__89224;
    wire N__89221;
    wire N__89216;
    wire N__89213;
    wire N__89208;
    wire N__89205;
    wire N__89202;
    wire N__89199;
    wire N__89198;
    wire N__89195;
    wire N__89192;
    wire N__89189;
    wire N__89184;
    wire N__89181;
    wire N__89180;
    wire N__89177;
    wire N__89174;
    wire N__89171;
    wire N__89166;
    wire N__89163;
    wire N__89160;
    wire N__89157;
    wire N__89154;
    wire N__89151;
    wire N__89148;
    wire N__89145;
    wire N__89144;
    wire N__89143;
    wire N__89140;
    wire N__89137;
    wire N__89134;
    wire N__89131;
    wire N__89124;
    wire N__89121;
    wire N__89118;
    wire N__89115;
    wire N__89112;
    wire N__89111;
    wire N__89110;
    wire N__89107;
    wire N__89104;
    wire N__89101;
    wire N__89094;
    wire N__89091;
    wire N__89088;
    wire N__89085;
    wire N__89082;
    wire N__89081;
    wire N__89080;
    wire N__89077;
    wire N__89074;
    wire N__89071;
    wire N__89064;
    wire N__89061;
    wire N__89058;
    wire N__89055;
    wire N__89052;
    wire N__89049;
    wire N__89046;
    wire N__89043;
    wire N__89040;
    wire N__89037;
    wire N__89034;
    wire N__89031;
    wire N__89028;
    wire N__89025;
    wire N__89022;
    wire N__89019;
    wire N__89018;
    wire N__89017;
    wire N__89014;
    wire N__89011;
    wire N__89008;
    wire N__89001;
    wire N__89000;
    wire N__88999;
    wire N__88996;
    wire N__88993;
    wire N__88990;
    wire N__88983;
    wire N__88982;
    wire N__88981;
    wire N__88978;
    wire N__88975;
    wire N__88972;
    wire N__88969;
    wire N__88962;
    wire N__88959;
    wire N__88958;
    wire N__88957;
    wire N__88954;
    wire N__88951;
    wire N__88948;
    wire N__88945;
    wire N__88938;
    wire N__88935;
    wire N__88932;
    wire N__88929;
    wire N__88926;
    wire N__88923;
    wire N__88920;
    wire N__88917;
    wire N__88914;
    wire N__88911;
    wire N__88910;
    wire N__88907;
    wire N__88906;
    wire N__88903;
    wire N__88900;
    wire N__88897;
    wire N__88890;
    wire N__88887;
    wire N__88884;
    wire N__88881;
    wire N__88878;
    wire N__88875;
    wire N__88874;
    wire N__88873;
    wire N__88870;
    wire N__88867;
    wire N__88864;
    wire N__88861;
    wire N__88854;
    wire N__88851;
    wire N__88848;
    wire N__88845;
    wire N__88842;
    wire N__88839;
    wire N__88838;
    wire N__88837;
    wire N__88834;
    wire N__88831;
    wire N__88828;
    wire N__88821;
    wire N__88818;
    wire N__88815;
    wire N__88812;
    wire N__88809;
    wire N__88806;
    wire N__88805;
    wire N__88804;
    wire N__88801;
    wire N__88798;
    wire N__88795;
    wire N__88788;
    wire N__88785;
    wire N__88782;
    wire N__88779;
    wire N__88776;
    wire N__88775;
    wire N__88774;
    wire N__88771;
    wire N__88768;
    wire N__88765;
    wire N__88762;
    wire N__88755;
    wire N__88752;
    wire N__88749;
    wire N__88746;
    wire N__88743;
    wire N__88742;
    wire N__88741;
    wire N__88738;
    wire N__88735;
    wire N__88732;
    wire N__88725;
    wire N__88722;
    wire N__88719;
    wire N__88716;
    wire N__88715;
    wire N__88714;
    wire N__88711;
    wire N__88708;
    wire N__88705;
    wire N__88698;
    wire N__88695;
    wire N__88694;
    wire N__88691;
    wire N__88688;
    wire N__88687;
    wire N__88682;
    wire N__88679;
    wire N__88674;
    wire N__88671;
    wire N__88670;
    wire N__88669;
    wire N__88666;
    wire N__88663;
    wire N__88660;
    wire N__88653;
    wire N__88650;
    wire N__88649;
    wire N__88648;
    wire N__88645;
    wire N__88642;
    wire N__88639;
    wire N__88632;
    wire N__88629;
    wire N__88626;
    wire N__88623;
    wire N__88620;
    wire N__88617;
    wire N__88614;
    wire N__88611;
    wire N__88608;
    wire N__88607;
    wire N__88606;
    wire N__88603;
    wire N__88600;
    wire N__88597;
    wire N__88594;
    wire N__88587;
    wire N__88584;
    wire N__88581;
    wire N__88578;
    wire N__88575;
    wire N__88572;
    wire N__88569;
    wire N__88568;
    wire N__88567;
    wire N__88564;
    wire N__88561;
    wire N__88558;
    wire N__88551;
    wire N__88548;
    wire N__88547;
    wire N__88546;
    wire N__88543;
    wire N__88540;
    wire N__88537;
    wire N__88530;
    wire N__88529;
    wire N__88528;
    wire N__88527;
    wire N__88526;
    wire N__88525;
    wire N__88522;
    wire N__88519;
    wire N__88516;
    wire N__88513;
    wire N__88510;
    wire N__88507;
    wire N__88502;
    wire N__88493;
    wire N__88488;
    wire N__88485;
    wire N__88482;
    wire N__88479;
    wire N__88478;
    wire N__88477;
    wire N__88476;
    wire N__88473;
    wire N__88470;
    wire N__88467;
    wire N__88464;
    wire N__88461;
    wire N__88452;
    wire N__88449;
    wire N__88446;
    wire N__88443;
    wire N__88442;
    wire N__88441;
    wire N__88440;
    wire N__88437;
    wire N__88434;
    wire N__88433;
    wire N__88432;
    wire N__88429;
    wire N__88426;
    wire N__88421;
    wire N__88418;
    wire N__88415;
    wire N__88414;
    wire N__88409;
    wire N__88406;
    wire N__88399;
    wire N__88392;
    wire N__88391;
    wire N__88390;
    wire N__88387;
    wire N__88384;
    wire N__88381;
    wire N__88380;
    wire N__88375;
    wire N__88372;
    wire N__88369;
    wire N__88366;
    wire N__88363;
    wire N__88356;
    wire N__88353;
    wire N__88352;
    wire N__88351;
    wire N__88348;
    wire N__88345;
    wire N__88342;
    wire N__88339;
    wire N__88332;
    wire N__88329;
    wire N__88328;
    wire N__88327;
    wire N__88324;
    wire N__88321;
    wire N__88318;
    wire N__88311;
    wire N__88308;
    wire N__88307;
    wire N__88306;
    wire N__88303;
    wire N__88300;
    wire N__88297;
    wire N__88292;
    wire N__88289;
    wire N__88286;
    wire N__88283;
    wire N__88278;
    wire N__88275;
    wire N__88274;
    wire N__88273;
    wire N__88270;
    wire N__88267;
    wire N__88264;
    wire N__88259;
    wire N__88256;
    wire N__88253;
    wire N__88250;
    wire N__88245;
    wire N__88242;
    wire N__88241;
    wire N__88240;
    wire N__88237;
    wire N__88234;
    wire N__88231;
    wire N__88228;
    wire N__88223;
    wire N__88220;
    wire N__88215;
    wire N__88212;
    wire N__88209;
    wire N__88208;
    wire N__88207;
    wire N__88204;
    wire N__88201;
    wire N__88198;
    wire N__88195;
    wire N__88190;
    wire N__88187;
    wire N__88182;
    wire N__88179;
    wire N__88178;
    wire N__88177;
    wire N__88174;
    wire N__88171;
    wire N__88168;
    wire N__88165;
    wire N__88158;
    wire N__88155;
    wire N__88152;
    wire N__88149;
    wire N__88148;
    wire N__88147;
    wire N__88144;
    wire N__88141;
    wire N__88138;
    wire N__88135;
    wire N__88128;
    wire N__88125;
    wire N__88124;
    wire N__88123;
    wire N__88122;
    wire N__88119;
    wire N__88116;
    wire N__88113;
    wire N__88110;
    wire N__88101;
    wire N__88100;
    wire N__88097;
    wire N__88094;
    wire N__88093;
    wire N__88088;
    wire N__88085;
    wire N__88082;
    wire N__88079;
    wire N__88074;
    wire N__88073;
    wire N__88070;
    wire N__88067;
    wire N__88062;
    wire N__88061;
    wire N__88058;
    wire N__88055;
    wire N__88050;
    wire N__88047;
    wire N__88044;
    wire N__88041;
    wire N__88038;
    wire N__88035;
    wire N__88034;
    wire N__88031;
    wire N__88028;
    wire N__88027;
    wire N__88022;
    wire N__88019;
    wire N__88016;
    wire N__88013;
    wire N__88008;
    wire N__88005;
    wire N__88004;
    wire N__88001;
    wire N__87998;
    wire N__87997;
    wire N__87992;
    wire N__87989;
    wire N__87986;
    wire N__87983;
    wire N__87978;
    wire N__87975;
    wire N__87974;
    wire N__87971;
    wire N__87968;
    wire N__87967;
    wire N__87962;
    wire N__87959;
    wire N__87956;
    wire N__87953;
    wire N__87948;
    wire N__87947;
    wire N__87946;
    wire N__87945;
    wire N__87944;
    wire N__87941;
    wire N__87938;
    wire N__87937;
    wire N__87936;
    wire N__87935;
    wire N__87932;
    wire N__87929;
    wire N__87926;
    wire N__87921;
    wire N__87918;
    wire N__87915;
    wire N__87912;
    wire N__87911;
    wire N__87904;
    wire N__87901;
    wire N__87892;
    wire N__87885;
    wire N__87882;
    wire N__87881;
    wire N__87880;
    wire N__87879;
    wire N__87878;
    wire N__87877;
    wire N__87874;
    wire N__87871;
    wire N__87868;
    wire N__87865;
    wire N__87862;
    wire N__87859;
    wire N__87854;
    wire N__87845;
    wire N__87840;
    wire N__87837;
    wire N__87834;
    wire N__87833;
    wire N__87832;
    wire N__87829;
    wire N__87826;
    wire N__87823;
    wire N__87820;
    wire N__87813;
    wire N__87810;
    wire N__87807;
    wire N__87806;
    wire N__87805;
    wire N__87802;
    wire N__87799;
    wire N__87796;
    wire N__87793;
    wire N__87788;
    wire N__87785;
    wire N__87780;
    wire N__87777;
    wire N__87776;
    wire N__87775;
    wire N__87772;
    wire N__87769;
    wire N__87766;
    wire N__87763;
    wire N__87758;
    wire N__87755;
    wire N__87750;
    wire N__87747;
    wire N__87746;
    wire N__87745;
    wire N__87742;
    wire N__87739;
    wire N__87736;
    wire N__87733;
    wire N__87728;
    wire N__87725;
    wire N__87720;
    wire N__87717;
    wire N__87716;
    wire N__87713;
    wire N__87710;
    wire N__87705;
    wire N__87704;
    wire N__87701;
    wire N__87698;
    wire N__87693;
    wire N__87692;
    wire N__87689;
    wire N__87686;
    wire N__87681;
    wire N__87680;
    wire N__87677;
    wire N__87674;
    wire N__87669;
    wire N__87666;
    wire N__87665;
    wire N__87662;
    wire N__87659;
    wire N__87654;
    wire N__87653;
    wire N__87650;
    wire N__87647;
    wire N__87642;
    wire N__87641;
    wire N__87638;
    wire N__87635;
    wire N__87630;
    wire N__87629;
    wire N__87626;
    wire N__87623;
    wire N__87618;
    wire N__87615;
    wire N__87614;
    wire N__87611;
    wire N__87608;
    wire N__87603;
    wire N__87602;
    wire N__87599;
    wire N__87596;
    wire N__87591;
    wire N__87590;
    wire N__87587;
    wire N__87584;
    wire N__87579;
    wire N__87578;
    wire N__87575;
    wire N__87572;
    wire N__87567;
    wire N__87564;
    wire N__87563;
    wire N__87560;
    wire N__87557;
    wire N__87552;
    wire N__87551;
    wire N__87548;
    wire N__87545;
    wire N__87540;
    wire N__87539;
    wire N__87536;
    wire N__87533;
    wire N__87532;
    wire N__87527;
    wire N__87524;
    wire N__87521;
    wire N__87518;
    wire N__87513;
    wire N__87510;
    wire N__87509;
    wire N__87508;
    wire N__87505;
    wire N__87502;
    wire N__87499;
    wire N__87494;
    wire N__87491;
    wire N__87488;
    wire N__87485;
    wire N__87480;
    wire N__87479;
    wire N__87476;
    wire N__87473;
    wire N__87472;
    wire N__87467;
    wire N__87464;
    wire N__87461;
    wire N__87458;
    wire N__87453;
    wire N__87450;
    wire N__87449;
    wire N__87446;
    wire N__87443;
    wire N__87442;
    wire N__87437;
    wire N__87434;
    wire N__87431;
    wire N__87428;
    wire N__87423;
    wire N__87422;
    wire N__87419;
    wire N__87416;
    wire N__87415;
    wire N__87410;
    wire N__87407;
    wire N__87404;
    wire N__87401;
    wire N__87396;
    wire N__87393;
    wire N__87392;
    wire N__87389;
    wire N__87386;
    wire N__87385;
    wire N__87382;
    wire N__87379;
    wire N__87376;
    wire N__87371;
    wire N__87368;
    wire N__87363;
    wire N__87362;
    wire N__87359;
    wire N__87356;
    wire N__87355;
    wire N__87350;
    wire N__87347;
    wire N__87344;
    wire N__87341;
    wire N__87336;
    wire N__87333;
    wire N__87332;
    wire N__87329;
    wire N__87326;
    wire N__87325;
    wire N__87320;
    wire N__87317;
    wire N__87314;
    wire N__87311;
    wire N__87306;
    wire N__87305;
    wire N__87304;
    wire N__87303;
    wire N__87302;
    wire N__87301;
    wire N__87300;
    wire N__87299;
    wire N__87298;
    wire N__87297;
    wire N__87296;
    wire N__87295;
    wire N__87294;
    wire N__87291;
    wire N__87290;
    wire N__87287;
    wire N__87284;
    wire N__87281;
    wire N__87278;
    wire N__87275;
    wire N__87274;
    wire N__87271;
    wire N__87270;
    wire N__87267;
    wire N__87264;
    wire N__87263;
    wire N__87260;
    wire N__87259;
    wire N__87256;
    wire N__87253;
    wire N__87248;
    wire N__87245;
    wire N__87242;
    wire N__87241;
    wire N__87240;
    wire N__87239;
    wire N__87234;
    wire N__87231;
    wire N__87228;
    wire N__87225;
    wire N__87222;
    wire N__87221;
    wire N__87220;
    wire N__87215;
    wire N__87212;
    wire N__87209;
    wire N__87206;
    wire N__87203;
    wire N__87200;
    wire N__87199;
    wire N__87198;
    wire N__87193;
    wire N__87188;
    wire N__87187;
    wire N__87184;
    wire N__87179;
    wire N__87176;
    wire N__87173;
    wire N__87170;
    wire N__87169;
    wire N__87168;
    wire N__87163;
    wire N__87160;
    wire N__87157;
    wire N__87154;
    wire N__87149;
    wire N__87148;
    wire N__87143;
    wire N__87140;
    wire N__87139;
    wire N__87136;
    wire N__87133;
    wire N__87130;
    wire N__87127;
    wire N__87126;
    wire N__87123;
    wire N__87118;
    wire N__87115;
    wire N__87112;
    wire N__87109;
    wire N__87106;
    wire N__87105;
    wire N__87102;
    wire N__87099;
    wire N__87094;
    wire N__87091;
    wire N__87088;
    wire N__87085;
    wire N__87080;
    wire N__87077;
    wire N__87074;
    wire N__87071;
    wire N__87066;
    wire N__87063;
    wire N__87060;
    wire N__87057;
    wire N__87054;
    wire N__87051;
    wire N__87048;
    wire N__87041;
    wire N__87036;
    wire N__87033;
    wire N__87028;
    wire N__87025;
    wire N__87018;
    wire N__87015;
    wire N__87012;
    wire N__87007;
    wire N__87004;
    wire N__86999;
    wire N__86996;
    wire N__86993;
    wire N__86988;
    wire N__86981;
    wire N__86970;
    wire N__86965;
    wire N__86960;
    wire N__86955;
    wire N__86954;
    wire N__86951;
    wire N__86948;
    wire N__86947;
    wire N__86946;
    wire N__86941;
    wire N__86938;
    wire N__86935;
    wire N__86930;
    wire N__86925;
    wire N__86922;
    wire N__86919;
    wire N__86916;
    wire N__86913;
    wire N__86912;
    wire N__86909;
    wire N__86906;
    wire N__86905;
    wire N__86900;
    wire N__86899;
    wire N__86896;
    wire N__86893;
    wire N__86890;
    wire N__86883;
    wire N__86882;
    wire N__86879;
    wire N__86876;
    wire N__86873;
    wire N__86870;
    wire N__86869;
    wire N__86866;
    wire N__86863;
    wire N__86860;
    wire N__86853;
    wire N__86850;
    wire N__86849;
    wire N__86846;
    wire N__86843;
    wire N__86838;
    wire N__86837;
    wire N__86834;
    wire N__86831;
    wire N__86826;
    wire N__86825;
    wire N__86822;
    wire N__86819;
    wire N__86814;
    wire N__86813;
    wire N__86810;
    wire N__86807;
    wire N__86802;
    wire N__86799;
    wire N__86798;
    wire N__86795;
    wire N__86792;
    wire N__86787;
    wire N__86786;
    wire N__86783;
    wire N__86780;
    wire N__86775;
    wire N__86774;
    wire N__86771;
    wire N__86768;
    wire N__86763;
    wire N__86762;
    wire N__86759;
    wire N__86756;
    wire N__86751;
    wire N__86748;
    wire N__86747;
    wire N__86744;
    wire N__86741;
    wire N__86736;
    wire N__86735;
    wire N__86732;
    wire N__86729;
    wire N__86724;
    wire N__86723;
    wire N__86720;
    wire N__86717;
    wire N__86712;
    wire N__86711;
    wire N__86708;
    wire N__86705;
    wire N__86700;
    wire N__86697;
    wire N__86696;
    wire N__86693;
    wire N__86690;
    wire N__86685;
    wire N__86684;
    wire N__86681;
    wire N__86678;
    wire N__86673;
    wire N__86672;
    wire N__86669;
    wire N__86666;
    wire N__86661;
    wire N__86660;
    wire N__86657;
    wire N__86654;
    wire N__86649;
    wire N__86646;
    wire N__86645;
    wire N__86642;
    wire N__86639;
    wire N__86638;
    wire N__86637;
    wire N__86636;
    wire N__86631;
    wire N__86628;
    wire N__86623;
    wire N__86620;
    wire N__86617;
    wire N__86610;
    wire N__86609;
    wire N__86608;
    wire N__86607;
    wire N__86606;
    wire N__86601;
    wire N__86600;
    wire N__86599;
    wire N__86596;
    wire N__86593;
    wire N__86590;
    wire N__86587;
    wire N__86584;
    wire N__86583;
    wire N__86580;
    wire N__86577;
    wire N__86570;
    wire N__86567;
    wire N__86564;
    wire N__86561;
    wire N__86558;
    wire N__86553;
    wire N__86544;
    wire N__86541;
    wire N__86540;
    wire N__86535;
    wire N__86532;
    wire N__86529;
    wire N__86526;
    wire N__86525;
    wire N__86522;
    wire N__86519;
    wire N__86516;
    wire N__86515;
    wire N__86512;
    wire N__86509;
    wire N__86506;
    wire N__86499;
    wire N__86496;
    wire N__86495;
    wire N__86492;
    wire N__86491;
    wire N__86490;
    wire N__86489;
    wire N__86486;
    wire N__86483;
    wire N__86480;
    wire N__86477;
    wire N__86474;
    wire N__86473;
    wire N__86470;
    wire N__86461;
    wire N__86458;
    wire N__86453;
    wire N__86448;
    wire N__86445;
    wire N__86444;
    wire N__86443;
    wire N__86440;
    wire N__86435;
    wire N__86430;
    wire N__86427;
    wire N__86426;
    wire N__86423;
    wire N__86420;
    wire N__86419;
    wire N__86416;
    wire N__86413;
    wire N__86412;
    wire N__86411;
    wire N__86408;
    wire N__86407;
    wire N__86404;
    wire N__86401;
    wire N__86398;
    wire N__86395;
    wire N__86392;
    wire N__86389;
    wire N__86386;
    wire N__86379;
    wire N__86376;
    wire N__86367;
    wire N__86364;
    wire N__86363;
    wire N__86360;
    wire N__86357;
    wire N__86354;
    wire N__86353;
    wire N__86352;
    wire N__86349;
    wire N__86348;
    wire N__86345;
    wire N__86342;
    wire N__86339;
    wire N__86336;
    wire N__86333;
    wire N__86330;
    wire N__86327;
    wire N__86324;
    wire N__86321;
    wire N__86310;
    wire N__86309;
    wire N__86308;
    wire N__86305;
    wire N__86300;
    wire N__86295;
    wire N__86292;
    wire N__86289;
    wire N__86286;
    wire N__86283;
    wire N__86280;
    wire N__86277;
    wire N__86274;
    wire N__86273;
    wire N__86272;
    wire N__86271;
    wire N__86268;
    wire N__86265;
    wire N__86262;
    wire N__86259;
    wire N__86258;
    wire N__86255;
    wire N__86252;
    wire N__86247;
    wire N__86244;
    wire N__86241;
    wire N__86238;
    wire N__86235;
    wire N__86226;
    wire N__86225;
    wire N__86222;
    wire N__86219;
    wire N__86214;
    wire N__86211;
    wire N__86208;
    wire N__86205;
    wire N__86202;
    wire N__86199;
    wire N__86198;
    wire N__86195;
    wire N__86192;
    wire N__86187;
    wire N__86186;
    wire N__86185;
    wire N__86184;
    wire N__86183;
    wire N__86182;
    wire N__86181;
    wire N__86178;
    wire N__86175;
    wire N__86170;
    wire N__86165;
    wire N__86162;
    wire N__86159;
    wire N__86156;
    wire N__86151;
    wire N__86142;
    wire N__86141;
    wire N__86140;
    wire N__86139;
    wire N__86138;
    wire N__86137;
    wire N__86132;
    wire N__86129;
    wire N__86126;
    wire N__86121;
    wire N__86120;
    wire N__86119;
    wire N__86118;
    wire N__86117;
    wire N__86116;
    wire N__86115;
    wire N__86114;
    wire N__86113;
    wire N__86112;
    wire N__86111;
    wire N__86110;
    wire N__86109;
    wire N__86108;
    wire N__86107;
    wire N__86106;
    wire N__86105;
    wire N__86104;
    wire N__86103;
    wire N__86094;
    wire N__86087;
    wire N__86082;
    wire N__86081;
    wire N__86080;
    wire N__86077;
    wire N__86074;
    wire N__86071;
    wire N__86064;
    wire N__86061;
    wire N__86056;
    wire N__86047;
    wire N__86046;
    wire N__86045;
    wire N__86044;
    wire N__86043;
    wire N__86042;
    wire N__86041;
    wire N__86038;
    wire N__86033;
    wire N__86030;
    wire N__86027;
    wire N__86022;
    wire N__86013;
    wire N__86010;
    wire N__86007;
    wire N__86002;
    wire N__85997;
    wire N__85994;
    wire N__85989;
    wire N__85986;
    wire N__85983;
    wire N__85972;
    wire N__85967;
    wire N__85964;
    wire N__85959;
    wire N__85954;
    wire N__85951;
    wire N__85946;
    wire N__85941;
    wire N__85938;
    wire N__85935;
    wire N__85932;
    wire N__85929;
    wire N__85926;
    wire N__85923;
    wire N__85922;
    wire N__85921;
    wire N__85920;
    wire N__85917;
    wire N__85914;
    wire N__85911;
    wire N__85908;
    wire N__85905;
    wire N__85902;
    wire N__85901;
    wire N__85900;
    wire N__85897;
    wire N__85896;
    wire N__85893;
    wire N__85888;
    wire N__85885;
    wire N__85882;
    wire N__85879;
    wire N__85876;
    wire N__85871;
    wire N__85868;
    wire N__85857;
    wire N__85854;
    wire N__85851;
    wire N__85848;
    wire N__85845;
    wire N__85844;
    wire N__85841;
    wire N__85840;
    wire N__85837;
    wire N__85834;
    wire N__85831;
    wire N__85830;
    wire N__85827;
    wire N__85824;
    wire N__85821;
    wire N__85818;
    wire N__85817;
    wire N__85814;
    wire N__85807;
    wire N__85804;
    wire N__85801;
    wire N__85798;
    wire N__85791;
    wire N__85788;
    wire N__85787;
    wire N__85784;
    wire N__85783;
    wire N__85782;
    wire N__85781;
    wire N__85778;
    wire N__85777;
    wire N__85774;
    wire N__85769;
    wire N__85766;
    wire N__85763;
    wire N__85760;
    wire N__85757;
    wire N__85754;
    wire N__85743;
    wire N__85740;
    wire N__85739;
    wire N__85736;
    wire N__85735;
    wire N__85732;
    wire N__85729;
    wire N__85726;
    wire N__85723;
    wire N__85720;
    wire N__85717;
    wire N__85716;
    wire N__85713;
    wire N__85708;
    wire N__85705;
    wire N__85700;
    wire N__85695;
    wire N__85692;
    wire N__85689;
    wire N__85688;
    wire N__85685;
    wire N__85684;
    wire N__85683;
    wire N__85680;
    wire N__85677;
    wire N__85676;
    wire N__85675;
    wire N__85674;
    wire N__85671;
    wire N__85668;
    wire N__85665;
    wire N__85662;
    wire N__85657;
    wire N__85654;
    wire N__85649;
    wire N__85646;
    wire N__85641;
    wire N__85632;
    wire N__85631;
    wire N__85630;
    wire N__85627;
    wire N__85626;
    wire N__85625;
    wire N__85622;
    wire N__85619;
    wire N__85616;
    wire N__85613;
    wire N__85610;
    wire N__85607;
    wire N__85604;
    wire N__85603;
    wire N__85600;
    wire N__85597;
    wire N__85594;
    wire N__85593;
    wire N__85590;
    wire N__85587;
    wire N__85584;
    wire N__85581;
    wire N__85576;
    wire N__85573;
    wire N__85570;
    wire N__85567;
    wire N__85564;
    wire N__85559;
    wire N__85548;
    wire N__85545;
    wire N__85542;
    wire N__85541;
    wire N__85538;
    wire N__85537;
    wire N__85534;
    wire N__85531;
    wire N__85528;
    wire N__85525;
    wire N__85522;
    wire N__85515;
    wire N__85512;
    wire N__85511;
    wire N__85510;
    wire N__85507;
    wire N__85506;
    wire N__85501;
    wire N__85500;
    wire N__85497;
    wire N__85494;
    wire N__85491;
    wire N__85490;
    wire N__85487;
    wire N__85484;
    wire N__85481;
    wire N__85478;
    wire N__85475;
    wire N__85464;
    wire N__85463;
    wire N__85460;
    wire N__85459;
    wire N__85456;
    wire N__85455;
    wire N__85452;
    wire N__85451;
    wire N__85448;
    wire N__85445;
    wire N__85442;
    wire N__85441;
    wire N__85438;
    wire N__85435;
    wire N__85432;
    wire N__85427;
    wire N__85424;
    wire N__85421;
    wire N__85418;
    wire N__85415;
    wire N__85412;
    wire N__85401;
    wire N__85398;
    wire N__85395;
    wire N__85392;
    wire N__85391;
    wire N__85388;
    wire N__85385;
    wire N__85380;
    wire N__85379;
    wire N__85378;
    wire N__85375;
    wire N__85374;
    wire N__85371;
    wire N__85368;
    wire N__85365;
    wire N__85362;
    wire N__85361;
    wire N__85358;
    wire N__85355;
    wire N__85352;
    wire N__85349;
    wire N__85346;
    wire N__85341;
    wire N__85338;
    wire N__85335;
    wire N__85326;
    wire N__85323;
    wire N__85322;
    wire N__85321;
    wire N__85318;
    wire N__85315;
    wire N__85312;
    wire N__85305;
    wire N__85302;
    wire N__85299;
    wire N__85296;
    wire N__85293;
    wire N__85290;
    wire N__85287;
    wire N__85284;
    wire N__85283;
    wire N__85282;
    wire N__85281;
    wire N__85280;
    wire N__85279;
    wire N__85278;
    wire N__85277;
    wire N__85276;
    wire N__85275;
    wire N__85274;
    wire N__85273;
    wire N__85270;
    wire N__85263;
    wire N__85256;
    wire N__85253;
    wire N__85252;
    wire N__85251;
    wire N__85250;
    wire N__85247;
    wire N__85246;
    wire N__85245;
    wire N__85242;
    wire N__85239;
    wire N__85236;
    wire N__85235;
    wire N__85234;
    wire N__85233;
    wire N__85232;
    wire N__85231;
    wire N__85230;
    wire N__85229;
    wire N__85228;
    wire N__85227;
    wire N__85220;
    wire N__85217;
    wire N__85216;
    wire N__85215;
    wire N__85214;
    wire N__85213;
    wire N__85212;
    wire N__85211;
    wire N__85210;
    wire N__85209;
    wire N__85206;
    wire N__85205;
    wire N__85204;
    wire N__85203;
    wire N__85200;
    wire N__85199;
    wire N__85198;
    wire N__85197;
    wire N__85194;
    wire N__85191;
    wire N__85184;
    wire N__85179;
    wire N__85178;
    wire N__85177;
    wire N__85176;
    wire N__85175;
    wire N__85174;
    wire N__85173;
    wire N__85172;
    wire N__85171;
    wire N__85166;
    wire N__85165;
    wire N__85164;
    wire N__85163;
    wire N__85162;
    wire N__85161;
    wire N__85160;
    wire N__85159;
    wire N__85158;
    wire N__85155;
    wire N__85152;
    wire N__85151;
    wire N__85150;
    wire N__85147;
    wire N__85146;
    wire N__85143;
    wire N__85142;
    wire N__85141;
    wire N__85136;
    wire N__85133;
    wire N__85128;
    wire N__85117;
    wire N__85108;
    wire N__85101;
    wire N__85100;
    wire N__85097;
    wire N__85096;
    wire N__85093;
    wire N__85088;
    wire N__85085;
    wire N__85082;
    wire N__85077;
    wire N__85076;
    wire N__85073;
    wire N__85072;
    wire N__85071;
    wire N__85070;
    wire N__85069;
    wire N__85068;
    wire N__85067;
    wire N__85066;
    wire N__85063;
    wire N__85060;
    wire N__85057;
    wire N__85056;
    wire N__85053;
    wire N__85052;
    wire N__85045;
    wire N__85042;
    wire N__85041;
    wire N__85040;
    wire N__85037;
    wire N__85034;
    wire N__85033;
    wire N__85030;
    wire N__85029;
    wire N__85028;
    wire N__85021;
    wire N__85012;
    wire N__85007;
    wire N__85004;
    wire N__85001;
    wire N__84998;
    wire N__84993;
    wire N__84990;
    wire N__84985;
    wire N__84980;
    wire N__84977;
    wire N__84974;
    wire N__84971;
    wire N__84968;
    wire N__84965;
    wire N__84958;
    wire N__84955;
    wire N__84950;
    wire N__84945;
    wire N__84940;
    wire N__84931;
    wire N__84928;
    wire N__84921;
    wire N__84918;
    wire N__84913;
    wire N__84906;
    wire N__84903;
    wire N__84898;
    wire N__84893;
    wire N__84890;
    wire N__84881;
    wire N__84878;
    wire N__84869;
    wire N__84864;
    wire N__84861;
    wire N__84850;
    wire N__84845;
    wire N__84838;
    wire N__84833;
    wire N__84824;
    wire N__84823;
    wire N__84822;
    wire N__84819;
    wire N__84816;
    wire N__84811;
    wire N__84806;
    wire N__84803;
    wire N__84794;
    wire N__84789;
    wire N__84774;
    wire N__84773;
    wire N__84770;
    wire N__84769;
    wire N__84766;
    wire N__84761;
    wire N__84760;
    wire N__84759;
    wire N__84756;
    wire N__84753;
    wire N__84750;
    wire N__84747;
    wire N__84746;
    wire N__84743;
    wire N__84738;
    wire N__84735;
    wire N__84732;
    wire N__84727;
    wire N__84724;
    wire N__84717;
    wire N__84716;
    wire N__84715;
    wire N__84714;
    wire N__84713;
    wire N__84712;
    wire N__84711;
    wire N__84710;
    wire N__84709;
    wire N__84708;
    wire N__84707;
    wire N__84706;
    wire N__84705;
    wire N__84704;
    wire N__84703;
    wire N__84702;
    wire N__84701;
    wire N__84700;
    wire N__84699;
    wire N__84698;
    wire N__84697;
    wire N__84696;
    wire N__84695;
    wire N__84694;
    wire N__84693;
    wire N__84692;
    wire N__84691;
    wire N__84690;
    wire N__84689;
    wire N__84688;
    wire N__84687;
    wire N__84686;
    wire N__84685;
    wire N__84684;
    wire N__84683;
    wire N__84682;
    wire N__84681;
    wire N__84680;
    wire N__84679;
    wire N__84678;
    wire N__84677;
    wire N__84674;
    wire N__84671;
    wire N__84670;
    wire N__84669;
    wire N__84662;
    wire N__84655;
    wire N__84652;
    wire N__84647;
    wire N__84640;
    wire N__84639;
    wire N__84638;
    wire N__84637;
    wire N__84634;
    wire N__84629;
    wire N__84628;
    wire N__84627;
    wire N__84626;
    wire N__84625;
    wire N__84624;
    wire N__84623;
    wire N__84620;
    wire N__84619;
    wire N__84618;
    wire N__84617;
    wire N__84616;
    wire N__84615;
    wire N__84614;
    wire N__84611;
    wire N__84606;
    wire N__84605;
    wire N__84604;
    wire N__84597;
    wire N__84590;
    wire N__84581;
    wire N__84574;
    wire N__84571;
    wire N__84562;
    wire N__84561;
    wire N__84560;
    wire N__84559;
    wire N__84558;
    wire N__84555;
    wire N__84554;
    wire N__84543;
    wire N__84538;
    wire N__84535;
    wire N__84530;
    wire N__84525;
    wire N__84522;
    wire N__84519;
    wire N__84516;
    wire N__84509;
    wire N__84506;
    wire N__84501;
    wire N__84498;
    wire N__84497;
    wire N__84488;
    wire N__84483;
    wire N__84480;
    wire N__84477;
    wire N__84476;
    wire N__84475;
    wire N__84470;
    wire N__84465;
    wire N__84462;
    wire N__84455;
    wire N__84454;
    wire N__84451;
    wire N__84448;
    wire N__84445;
    wire N__84442;
    wire N__84439;
    wire N__84436;
    wire N__84427;
    wire N__84426;
    wire N__84425;
    wire N__84424;
    wire N__84423;
    wire N__84422;
    wire N__84417;
    wire N__84414;
    wire N__84411;
    wire N__84402;
    wire N__84399;
    wire N__84390;
    wire N__84385;
    wire N__84380;
    wire N__84375;
    wire N__84372;
    wire N__84369;
    wire N__84364;
    wire N__84359;
    wire N__84354;
    wire N__84353;
    wire N__84352;
    wire N__84351;
    wire N__84350;
    wire N__84347;
    wire N__84342;
    wire N__84337;
    wire N__84328;
    wire N__84323;
    wire N__84316;
    wire N__84307;
    wire N__84304;
    wire N__84299;
    wire N__84294;
    wire N__84273;
    wire N__84270;
    wire N__84269;
    wire N__84266;
    wire N__84263;
    wire N__84260;
    wire N__84255;
    wire N__84254;
    wire N__84251;
    wire N__84248;
    wire N__84247;
    wire N__84246;
    wire N__84245;
    wire N__84244;
    wire N__84243;
    wire N__84242;
    wire N__84241;
    wire N__84240;
    wire N__84237;
    wire N__84236;
    wire N__84235;
    wire N__84234;
    wire N__84233;
    wire N__84232;
    wire N__84231;
    wire N__84230;
    wire N__84227;
    wire N__84222;
    wire N__84221;
    wire N__84218;
    wire N__84217;
    wire N__84214;
    wire N__84207;
    wire N__84204;
    wire N__84203;
    wire N__84200;
    wire N__84197;
    wire N__84190;
    wire N__84187;
    wire N__84184;
    wire N__84181;
    wire N__84180;
    wire N__84175;
    wire N__84172;
    wire N__84171;
    wire N__84168;
    wire N__84165;
    wire N__84162;
    wire N__84157;
    wire N__84154;
    wire N__84147;
    wire N__84146;
    wire N__84143;
    wire N__84142;
    wire N__84139;
    wire N__84136;
    wire N__84133;
    wire N__84128;
    wire N__84125;
    wire N__84122;
    wire N__84121;
    wire N__84118;
    wire N__84117;
    wire N__84116;
    wire N__84111;
    wire N__84106;
    wire N__84103;
    wire N__84100;
    wire N__84097;
    wire N__84092;
    wire N__84089;
    wire N__84084;
    wire N__84081;
    wire N__84078;
    wire N__84075;
    wire N__84072;
    wire N__84071;
    wire N__84068;
    wire N__84057;
    wire N__84050;
    wire N__84047;
    wire N__84044;
    wire N__84039;
    wire N__84036;
    wire N__84033;
    wire N__84032;
    wire N__84031;
    wire N__84030;
    wire N__84029;
    wire N__84026;
    wire N__84023;
    wire N__84018;
    wire N__84013;
    wire N__84010;
    wire N__84007;
    wire N__84004;
    wire N__84001;
    wire N__83998;
    wire N__83979;
    wire N__83978;
    wire N__83977;
    wire N__83976;
    wire N__83975;
    wire N__83974;
    wire N__83973;
    wire N__83972;
    wire N__83971;
    wire N__83970;
    wire N__83969;
    wire N__83968;
    wire N__83967;
    wire N__83966;
    wire N__83965;
    wire N__83964;
    wire N__83963;
    wire N__83962;
    wire N__83961;
    wire N__83960;
    wire N__83959;
    wire N__83958;
    wire N__83957;
    wire N__83956;
    wire N__83955;
    wire N__83954;
    wire N__83953;
    wire N__83944;
    wire N__83943;
    wire N__83942;
    wire N__83941;
    wire N__83938;
    wire N__83937;
    wire N__83936;
    wire N__83933;
    wire N__83928;
    wire N__83921;
    wire N__83920;
    wire N__83919;
    wire N__83918;
    wire N__83915;
    wire N__83914;
    wire N__83913;
    wire N__83912;
    wire N__83911;
    wire N__83910;
    wire N__83909;
    wire N__83906;
    wire N__83899;
    wire N__83894;
    wire N__83893;
    wire N__83892;
    wire N__83891;
    wire N__83888;
    wire N__83885;
    wire N__83882;
    wire N__83877;
    wire N__83872;
    wire N__83869;
    wire N__83868;
    wire N__83867;
    wire N__83864;
    wire N__83863;
    wire N__83860;
    wire N__83855;
    wire N__83852;
    wire N__83849;
    wire N__83844;
    wire N__83841;
    wire N__83836;
    wire N__83829;
    wire N__83826;
    wire N__83823;
    wire N__83820;
    wire N__83813;
    wire N__83812;
    wire N__83811;
    wire N__83810;
    wire N__83809;
    wire N__83808;
    wire N__83807;
    wire N__83804;
    wire N__83797;
    wire N__83794;
    wire N__83789;
    wire N__83786;
    wire N__83781;
    wire N__83776;
    wire N__83773;
    wire N__83770;
    wire N__83767;
    wire N__83764;
    wire N__83761;
    wire N__83756;
    wire N__83751;
    wire N__83744;
    wire N__83733;
    wire N__83732;
    wire N__83729;
    wire N__83724;
    wire N__83717;
    wire N__83712;
    wire N__83707;
    wire N__83700;
    wire N__83699;
    wire N__83698;
    wire N__83695;
    wire N__83692;
    wire N__83689;
    wire N__83676;
    wire N__83673;
    wire N__83670;
    wire N__83665;
    wire N__83662;
    wire N__83657;
    wire N__83654;
    wire N__83651;
    wire N__83646;
    wire N__83641;
    wire N__83630;
    wire N__83619;
    wire N__83618;
    wire N__83617;
    wire N__83616;
    wire N__83613;
    wire N__83610;
    wire N__83605;
    wire N__83602;
    wire N__83599;
    wire N__83596;
    wire N__83595;
    wire N__83594;
    wire N__83591;
    wire N__83586;
    wire N__83583;
    wire N__83580;
    wire N__83577;
    wire N__83574;
    wire N__83571;
    wire N__83568;
    wire N__83565;
    wire N__83562;
    wire N__83553;
    wire N__83550;
    wire N__83547;
    wire N__83544;
    wire N__83541;
    wire N__83538;
    wire N__83535;
    wire N__83534;
    wire N__83533;
    wire N__83530;
    wire N__83529;
    wire N__83526;
    wire N__83523;
    wire N__83522;
    wire N__83519;
    wire N__83516;
    wire N__83513;
    wire N__83510;
    wire N__83507;
    wire N__83504;
    wire N__83501;
    wire N__83498;
    wire N__83495;
    wire N__83484;
    wire N__83483;
    wire N__83482;
    wire N__83481;
    wire N__83478;
    wire N__83477;
    wire N__83474;
    wire N__83471;
    wire N__83468;
    wire N__83467;
    wire N__83466;
    wire N__83463;
    wire N__83460;
    wire N__83455;
    wire N__83452;
    wire N__83449;
    wire N__83446;
    wire N__83443;
    wire N__83438;
    wire N__83433;
    wire N__83424;
    wire N__83423;
    wire N__83422;
    wire N__83421;
    wire N__83418;
    wire N__83415;
    wire N__83412;
    wire N__83409;
    wire N__83404;
    wire N__83401;
    wire N__83398;
    wire N__83395;
    wire N__83392;
    wire N__83385;
    wire N__83382;
    wire N__83379;
    wire N__83376;
    wire N__83373;
    wire N__83370;
    wire N__83367;
    wire N__83364;
    wire N__83361;
    wire N__83358;
    wire N__83355;
    wire N__83352;
    wire N__83349;
    wire N__83346;
    wire N__83343;
    wire N__83342;
    wire N__83339;
    wire N__83336;
    wire N__83331;
    wire N__83330;
    wire N__83327;
    wire N__83324;
    wire N__83321;
    wire N__83320;
    wire N__83317;
    wire N__83316;
    wire N__83313;
    wire N__83310;
    wire N__83309;
    wire N__83306;
    wire N__83303;
    wire N__83300;
    wire N__83297;
    wire N__83294;
    wire N__83291;
    wire N__83280;
    wire N__83279;
    wire N__83276;
    wire N__83273;
    wire N__83272;
    wire N__83271;
    wire N__83268;
    wire N__83267;
    wire N__83264;
    wire N__83261;
    wire N__83258;
    wire N__83255;
    wire N__83252;
    wire N__83249;
    wire N__83244;
    wire N__83241;
    wire N__83232;
    wire N__83229;
    wire N__83228;
    wire N__83225;
    wire N__83224;
    wire N__83221;
    wire N__83220;
    wire N__83217;
    wire N__83214;
    wire N__83211;
    wire N__83208;
    wire N__83205;
    wire N__83202;
    wire N__83199;
    wire N__83190;
    wire N__83187;
    wire N__83186;
    wire N__83183;
    wire N__83180;
    wire N__83179;
    wire N__83178;
    wire N__83175;
    wire N__83170;
    wire N__83169;
    wire N__83166;
    wire N__83161;
    wire N__83158;
    wire N__83151;
    wire N__83148;
    wire N__83147;
    wire N__83142;
    wire N__83139;
    wire N__83138;
    wire N__83137;
    wire N__83132;
    wire N__83129;
    wire N__83128;
    wire N__83127;
    wire N__83124;
    wire N__83121;
    wire N__83118;
    wire N__83117;
    wire N__83114;
    wire N__83111;
    wire N__83106;
    wire N__83103;
    wire N__83100;
    wire N__83097;
    wire N__83094;
    wire N__83085;
    wire N__83082;
    wire N__83081;
    wire N__83078;
    wire N__83075;
    wire N__83070;
    wire N__83067;
    wire N__83064;
    wire N__83061;
    wire N__83060;
    wire N__83059;
    wire N__83058;
    wire N__83055;
    wire N__83054;
    wire N__83051;
    wire N__83048;
    wire N__83045;
    wire N__83042;
    wire N__83041;
    wire N__83038;
    wire N__83035;
    wire N__83032;
    wire N__83027;
    wire N__83024;
    wire N__83013;
    wire N__83012;
    wire N__83009;
    wire N__83006;
    wire N__83001;
    wire N__83000;
    wire N__82997;
    wire N__82994;
    wire N__82989;
    wire N__82986;
    wire N__82985;
    wire N__82982;
    wire N__82979;
    wire N__82978;
    wire N__82973;
    wire N__82970;
    wire N__82967;
    wire N__82964;
    wire N__82959;
    wire N__82956;
    wire N__82955;
    wire N__82952;
    wire N__82949;
    wire N__82944;
    wire N__82943;
    wire N__82940;
    wire N__82937;
    wire N__82932;
    wire N__82929;
    wire N__82928;
    wire N__82925;
    wire N__82922;
    wire N__82917;
    wire N__82916;
    wire N__82913;
    wire N__82910;
    wire N__82905;
    wire N__82902;
    wire N__82901;
    wire N__82898;
    wire N__82895;
    wire N__82890;
    wire N__82889;
    wire N__82886;
    wire N__82883;
    wire N__82878;
    wire N__82875;
    wire N__82874;
    wire N__82871;
    wire N__82868;
    wire N__82863;
    wire N__82862;
    wire N__82859;
    wire N__82856;
    wire N__82851;
    wire N__82850;
    wire N__82849;
    wire N__82848;
    wire N__82847;
    wire N__82846;
    wire N__82845;
    wire N__82844;
    wire N__82843;
    wire N__82842;
    wire N__82841;
    wire N__82840;
    wire N__82839;
    wire N__82838;
    wire N__82837;
    wire N__82836;
    wire N__82833;
    wire N__82830;
    wire N__82827;
    wire N__82824;
    wire N__82821;
    wire N__82818;
    wire N__82815;
    wire N__82812;
    wire N__82809;
    wire N__82806;
    wire N__82803;
    wire N__82800;
    wire N__82797;
    wire N__82794;
    wire N__82791;
    wire N__82788;
    wire N__82781;
    wire N__82774;
    wire N__82765;
    wire N__82756;
    wire N__82751;
    wire N__82740;
    wire N__82737;
    wire N__82734;
    wire N__82731;
    wire N__82728;
    wire N__82727;
    wire N__82724;
    wire N__82721;
    wire N__82720;
    wire N__82715;
    wire N__82712;
    wire N__82707;
    wire N__82704;
    wire N__82701;
    wire N__82700;
    wire N__82697;
    wire N__82694;
    wire N__82693;
    wire N__82688;
    wire N__82685;
    wire N__82680;
    wire N__82677;
    wire N__82674;
    wire N__82673;
    wire N__82670;
    wire N__82667;
    wire N__82666;
    wire N__82661;
    wire N__82658;
    wire N__82655;
    wire N__82652;
    wire N__82647;
    wire N__82644;
    wire N__82643;
    wire N__82640;
    wire N__82637;
    wire N__82632;
    wire N__82631;
    wire N__82628;
    wire N__82625;
    wire N__82620;
    wire N__82617;
    wire N__82616;
    wire N__82613;
    wire N__82610;
    wire N__82609;
    wire N__82604;
    wire N__82601;
    wire N__82598;
    wire N__82595;
    wire N__82590;
    wire N__82587;
    wire N__82586;
    wire N__82583;
    wire N__82580;
    wire N__82575;
    wire N__82574;
    wire N__82571;
    wire N__82568;
    wire N__82563;
    wire N__82560;
    wire N__82559;
    wire N__82556;
    wire N__82553;
    wire N__82552;
    wire N__82547;
    wire N__82544;
    wire N__82541;
    wire N__82538;
    wire N__82533;
    wire N__82530;
    wire N__82529;
    wire N__82526;
    wire N__82523;
    wire N__82522;
    wire N__82517;
    wire N__82514;
    wire N__82511;
    wire N__82508;
    wire N__82503;
    wire N__82500;
    wire N__82499;
    wire N__82496;
    wire N__82493;
    wire N__82488;
    wire N__82487;
    wire N__82484;
    wire N__82481;
    wire N__82476;
    wire N__82473;
    wire N__82472;
    wire N__82469;
    wire N__82466;
    wire N__82463;
    wire N__82458;
    wire N__82457;
    wire N__82454;
    wire N__82451;
    wire N__82448;
    wire N__82443;
    wire N__82440;
    wire N__82439;
    wire N__82436;
    wire N__82433;
    wire N__82430;
    wire N__82425;
    wire N__82422;
    wire N__82419;
    wire N__82418;
    wire N__82417;
    wire N__82414;
    wire N__82411;
    wire N__82410;
    wire N__82407;
    wire N__82402;
    wire N__82399;
    wire N__82396;
    wire N__82393;
    wire N__82388;
    wire N__82383;
    wire N__82380;
    wire N__82379;
    wire N__82376;
    wire N__82373;
    wire N__82368;
    wire N__82367;
    wire N__82364;
    wire N__82361;
    wire N__82356;
    wire N__82353;
    wire N__82352;
    wire N__82349;
    wire N__82346;
    wire N__82345;
    wire N__82340;
    wire N__82337;
    wire N__82334;
    wire N__82331;
    wire N__82326;
    wire N__82323;
    wire N__82322;
    wire N__82319;
    wire N__82316;
    wire N__82311;
    wire N__82310;
    wire N__82307;
    wire N__82304;
    wire N__82299;
    wire N__82296;
    wire N__82295;
    wire N__82292;
    wire N__82289;
    wire N__82284;
    wire N__82283;
    wire N__82280;
    wire N__82277;
    wire N__82272;
    wire N__82269;
    wire N__82268;
    wire N__82265;
    wire N__82262;
    wire N__82257;
    wire N__82256;
    wire N__82253;
    wire N__82250;
    wire N__82245;
    wire N__82242;
    wire N__82241;
    wire N__82238;
    wire N__82235;
    wire N__82234;
    wire N__82229;
    wire N__82226;
    wire N__82223;
    wire N__82220;
    wire N__82215;
    wire N__82214;
    wire N__82213;
    wire N__82212;
    wire N__82211;
    wire N__82210;
    wire N__82207;
    wire N__82204;
    wire N__82201;
    wire N__82198;
    wire N__82195;
    wire N__82192;
    wire N__82187;
    wire N__82178;
    wire N__82173;
    wire N__82170;
    wire N__82167;
    wire N__82164;
    wire N__82161;
    wire N__82158;
    wire N__82155;
    wire N__82152;
    wire N__82149;
    wire N__82146;
    wire N__82143;
    wire N__82140;
    wire N__82137;
    wire N__82134;
    wire N__82131;
    wire N__82128;
    wire N__82125;
    wire N__82122;
    wire N__82119;
    wire N__82116;
    wire N__82113;
    wire N__82112;
    wire N__82109;
    wire N__82106;
    wire N__82103;
    wire N__82098;
    wire N__82095;
    wire N__82092;
    wire N__82091;
    wire N__82088;
    wire N__82085;
    wire N__82082;
    wire N__82077;
    wire N__82074;
    wire N__82071;
    wire N__82068;
    wire N__82065;
    wire N__82062;
    wire N__82059;
    wire N__82056;
    wire N__82053;
    wire N__82050;
    wire N__82047;
    wire N__82044;
    wire N__82041;
    wire N__82038;
    wire N__82035;
    wire N__82032;
    wire N__82029;
    wire N__82026;
    wire N__82023;
    wire N__82020;
    wire N__82017;
    wire N__82014;
    wire N__82011;
    wire N__82008;
    wire N__82007;
    wire N__82004;
    wire N__82001;
    wire N__82000;
    wire N__81999;
    wire N__81994;
    wire N__81991;
    wire N__81988;
    wire N__81985;
    wire N__81982;
    wire N__81975;
    wire N__81972;
    wire N__81971;
    wire N__81970;
    wire N__81967;
    wire N__81964;
    wire N__81961;
    wire N__81960;
    wire N__81957;
    wire N__81954;
    wire N__81951;
    wire N__81948;
    wire N__81943;
    wire N__81940;
    wire N__81933;
    wire N__81930;
    wire N__81929;
    wire N__81928;
    wire N__81925;
    wire N__81922;
    wire N__81919;
    wire N__81916;
    wire N__81913;
    wire N__81910;
    wire N__81909;
    wire N__81906;
    wire N__81903;
    wire N__81900;
    wire N__81897;
    wire N__81892;
    wire N__81889;
    wire N__81882;
    wire N__81879;
    wire N__81878;
    wire N__81877;
    wire N__81874;
    wire N__81871;
    wire N__81868;
    wire N__81861;
    wire N__81860;
    wire N__81857;
    wire N__81854;
    wire N__81851;
    wire N__81846;
    wire N__81843;
    wire N__81842;
    wire N__81841;
    wire N__81838;
    wire N__81835;
    wire N__81832;
    wire N__81831;
    wire N__81826;
    wire N__81823;
    wire N__81820;
    wire N__81817;
    wire N__81814;
    wire N__81807;
    wire N__81804;
    wire N__81803;
    wire N__81800;
    wire N__81797;
    wire N__81796;
    wire N__81791;
    wire N__81788;
    wire N__81787;
    wire N__81784;
    wire N__81781;
    wire N__81778;
    wire N__81775;
    wire N__81772;
    wire N__81765;
    wire N__81762;
    wire N__81759;
    wire N__81756;
    wire N__81753;
    wire N__81750;
    wire N__81749;
    wire N__81746;
    wire N__81743;
    wire N__81738;
    wire N__81735;
    wire N__81732;
    wire N__81729;
    wire N__81726;
    wire N__81723;
    wire N__81722;
    wire N__81719;
    wire N__81716;
    wire N__81711;
    wire N__81708;
    wire N__81705;
    wire N__81702;
    wire N__81699;
    wire N__81698;
    wire N__81695;
    wire N__81692;
    wire N__81687;
    wire N__81684;
    wire N__81681;
    wire N__81678;
    wire N__81677;
    wire N__81676;
    wire N__81673;
    wire N__81670;
    wire N__81667;
    wire N__81660;
    wire N__81657;
    wire N__81654;
    wire N__81651;
    wire N__81650;
    wire N__81649;
    wire N__81646;
    wire N__81643;
    wire N__81640;
    wire N__81633;
    wire N__81632;
    wire N__81631;
    wire N__81630;
    wire N__81629;
    wire N__81628;
    wire N__81627;
    wire N__81626;
    wire N__81625;
    wire N__81624;
    wire N__81621;
    wire N__81618;
    wire N__81615;
    wire N__81612;
    wire N__81609;
    wire N__81606;
    wire N__81603;
    wire N__81600;
    wire N__81597;
    wire N__81594;
    wire N__81589;
    wire N__81580;
    wire N__81571;
    wire N__81568;
    wire N__81567;
    wire N__81562;
    wire N__81559;
    wire N__81556;
    wire N__81549;
    wire N__81548;
    wire N__81547;
    wire N__81544;
    wire N__81541;
    wire N__81538;
    wire N__81533;
    wire N__81530;
    wire N__81525;
    wire N__81522;
    wire N__81521;
    wire N__81520;
    wire N__81517;
    wire N__81514;
    wire N__81511;
    wire N__81506;
    wire N__81503;
    wire N__81500;
    wire N__81497;
    wire N__81492;
    wire N__81491;
    wire N__81490;
    wire N__81487;
    wire N__81484;
    wire N__81481;
    wire N__81478;
    wire N__81475;
    wire N__81470;
    wire N__81467;
    wire N__81462;
    wire N__81459;
    wire N__81458;
    wire N__81455;
    wire N__81454;
    wire N__81451;
    wire N__81448;
    wire N__81445;
    wire N__81442;
    wire N__81437;
    wire N__81434;
    wire N__81429;
    wire N__81426;
    wire N__81423;
    wire N__81420;
    wire N__81417;
    wire N__81414;
    wire N__81411;
    wire N__81410;
    wire N__81409;
    wire N__81408;
    wire N__81407;
    wire N__81406;
    wire N__81405;
    wire N__81404;
    wire N__81403;
    wire N__81400;
    wire N__81397;
    wire N__81394;
    wire N__81391;
    wire N__81388;
    wire N__81385;
    wire N__81382;
    wire N__81379;
    wire N__81376;
    wire N__81369;
    wire N__81360;
    wire N__81355;
    wire N__81348;
    wire N__81345;
    wire N__81344;
    wire N__81343;
    wire N__81342;
    wire N__81341;
    wire N__81340;
    wire N__81337;
    wire N__81334;
    wire N__81331;
    wire N__81328;
    wire N__81325;
    wire N__81322;
    wire N__81317;
    wire N__81308;
    wire N__81303;
    wire N__81300;
    wire N__81297;
    wire N__81294;
    wire N__81293;
    wire N__81290;
    wire N__81287;
    wire N__81284;
    wire N__81279;
    wire N__81276;
    wire N__81275;
    wire N__81272;
    wire N__81271;
    wire N__81270;
    wire N__81267;
    wire N__81264;
    wire N__81261;
    wire N__81260;
    wire N__81257;
    wire N__81254;
    wire N__81249;
    wire N__81248;
    wire N__81247;
    wire N__81246;
    wire N__81245;
    wire N__81244;
    wire N__81243;
    wire N__81242;
    wire N__81241;
    wire N__81240;
    wire N__81237;
    wire N__81234;
    wire N__81229;
    wire N__81226;
    wire N__81225;
    wire N__81224;
    wire N__81223;
    wire N__81222;
    wire N__81221;
    wire N__81220;
    wire N__81217;
    wire N__81214;
    wire N__81213;
    wire N__81210;
    wire N__81207;
    wire N__81204;
    wire N__81203;
    wire N__81202;
    wire N__81201;
    wire N__81196;
    wire N__81191;
    wire N__81184;
    wire N__81181;
    wire N__81178;
    wire N__81175;
    wire N__81174;
    wire N__81173;
    wire N__81172;
    wire N__81169;
    wire N__81166;
    wire N__81163;
    wire N__81160;
    wire N__81157;
    wire N__81154;
    wire N__81151;
    wire N__81148;
    wire N__81145;
    wire N__81142;
    wire N__81139;
    wire N__81136;
    wire N__81133;
    wire N__81126;
    wire N__81123;
    wire N__81120;
    wire N__81117;
    wire N__81116;
    wire N__81113;
    wire N__81110;
    wire N__81105;
    wire N__81104;
    wire N__81103;
    wire N__81100;
    wire N__81097;
    wire N__81094;
    wire N__81089;
    wire N__81084;
    wire N__81081;
    wire N__81076;
    wire N__81073;
    wire N__81066;
    wire N__81063;
    wire N__81060;
    wire N__81055;
    wire N__81052;
    wire N__81047;
    wire N__81036;
    wire N__81027;
    wire N__81026;
    wire N__81025;
    wire N__81022;
    wire N__81015;
    wire N__81012;
    wire N__81007;
    wire N__81004;
    wire N__81001;
    wire N__80998;
    wire N__80995;
    wire N__80990;
    wire N__80979;
    wire N__80978;
    wire N__80977;
    wire N__80976;
    wire N__80975;
    wire N__80974;
    wire N__80971;
    wire N__80970;
    wire N__80969;
    wire N__80968;
    wire N__80963;
    wire N__80960;
    wire N__80957;
    wire N__80956;
    wire N__80955;
    wire N__80954;
    wire N__80953;
    wire N__80950;
    wire N__80943;
    wire N__80940;
    wire N__80937;
    wire N__80934;
    wire N__80933;
    wire N__80932;
    wire N__80931;
    wire N__80930;
    wire N__80927;
    wire N__80926;
    wire N__80925;
    wire N__80924;
    wire N__80923;
    wire N__80922;
    wire N__80921;
    wire N__80918;
    wire N__80915;
    wire N__80912;
    wire N__80911;
    wire N__80910;
    wire N__80907;
    wire N__80906;
    wire N__80903;
    wire N__80900;
    wire N__80895;
    wire N__80892;
    wire N__80889;
    wire N__80884;
    wire N__80881;
    wire N__80878;
    wire N__80877;
    wire N__80876;
    wire N__80873;
    wire N__80870;
    wire N__80867;
    wire N__80866;
    wire N__80865;
    wire N__80862;
    wire N__80857;
    wire N__80850;
    wire N__80845;
    wire N__80842;
    wire N__80839;
    wire N__80836;
    wire N__80825;
    wire N__80822;
    wire N__80819;
    wire N__80814;
    wire N__80809;
    wire N__80808;
    wire N__80807;
    wire N__80804;
    wire N__80799;
    wire N__80796;
    wire N__80793;
    wire N__80790;
    wire N__80785;
    wire N__80782;
    wire N__80777;
    wire N__80772;
    wire N__80767;
    wire N__80764;
    wire N__80761;
    wire N__80758;
    wire N__80749;
    wire N__80746;
    wire N__80741;
    wire N__80736;
    wire N__80721;
    wire N__80720;
    wire N__80719;
    wire N__80718;
    wire N__80713;
    wire N__80712;
    wire N__80711;
    wire N__80710;
    wire N__80709;
    wire N__80708;
    wire N__80705;
    wire N__80702;
    wire N__80701;
    wire N__80700;
    wire N__80697;
    wire N__80694;
    wire N__80693;
    wire N__80690;
    wire N__80689;
    wire N__80688;
    wire N__80685;
    wire N__80684;
    wire N__80681;
    wire N__80680;
    wire N__80677;
    wire N__80676;
    wire N__80671;
    wire N__80668;
    wire N__80665;
    wire N__80664;
    wire N__80663;
    wire N__80658;
    wire N__80655;
    wire N__80652;
    wire N__80647;
    wire N__80644;
    wire N__80641;
    wire N__80640;
    wire N__80637;
    wire N__80634;
    wire N__80633;
    wire N__80630;
    wire N__80627;
    wire N__80624;
    wire N__80619;
    wire N__80618;
    wire N__80617;
    wire N__80612;
    wire N__80607;
    wire N__80602;
    wire N__80601;
    wire N__80596;
    wire N__80593;
    wire N__80592;
    wire N__80587;
    wire N__80584;
    wire N__80575;
    wire N__80572;
    wire N__80569;
    wire N__80564;
    wire N__80561;
    wire N__80558;
    wire N__80555;
    wire N__80554;
    wire N__80553;
    wire N__80548;
    wire N__80547;
    wire N__80544;
    wire N__80541;
    wire N__80538;
    wire N__80537;
    wire N__80534;
    wire N__80531;
    wire N__80526;
    wire N__80523;
    wire N__80520;
    wire N__80519;
    wire N__80514;
    wire N__80511;
    wire N__80508;
    wire N__80505;
    wire N__80500;
    wire N__80499;
    wire N__80498;
    wire N__80495;
    wire N__80492;
    wire N__80487;
    wire N__80482;
    wire N__80479;
    wire N__80476;
    wire N__80473;
    wire N__80466;
    wire N__80463;
    wire N__80460;
    wire N__80457;
    wire N__80452;
    wire N__80449;
    wire N__80440;
    wire N__80427;
    wire N__80424;
    wire N__80423;
    wire N__80422;
    wire N__80419;
    wire N__80416;
    wire N__80413;
    wire N__80412;
    wire N__80411;
    wire N__80410;
    wire N__80409;
    wire N__80408;
    wire N__80407;
    wire N__80406;
    wire N__80403;
    wire N__80398;
    wire N__80397;
    wire N__80396;
    wire N__80395;
    wire N__80392;
    wire N__80387;
    wire N__80386;
    wire N__80385;
    wire N__80382;
    wire N__80375;
    wire N__80370;
    wire N__80367;
    wire N__80366;
    wire N__80363;
    wire N__80362;
    wire N__80361;
    wire N__80358;
    wire N__80355;
    wire N__80352;
    wire N__80349;
    wire N__80344;
    wire N__80337;
    wire N__80336;
    wire N__80333;
    wire N__80332;
    wire N__80331;
    wire N__80328;
    wire N__80325;
    wire N__80322;
    wire N__80321;
    wire N__80320;
    wire N__80319;
    wire N__80316;
    wire N__80313;
    wire N__80308;
    wire N__80303;
    wire N__80300;
    wire N__80299;
    wire N__80298;
    wire N__80295;
    wire N__80292;
    wire N__80289;
    wire N__80286;
    wire N__80283;
    wire N__80280;
    wire N__80277;
    wire N__80274;
    wire N__80273;
    wire N__80270;
    wire N__80269;
    wire N__80268;
    wire N__80267;
    wire N__80266;
    wire N__80265;
    wire N__80258;
    wire N__80253;
    wire N__80250;
    wire N__80247;
    wire N__80242;
    wire N__80235;
    wire N__80232;
    wire N__80227;
    wire N__80222;
    wire N__80217;
    wire N__80212;
    wire N__80209;
    wire N__80206;
    wire N__80203;
    wire N__80200;
    wire N__80197;
    wire N__80192;
    wire N__80187;
    wire N__80182;
    wire N__80175;
    wire N__80172;
    wire N__80165;
    wire N__80162;
    wire N__80155;
    wire N__80152;
    wire N__80145;
    wire N__80144;
    wire N__80141;
    wire N__80138;
    wire N__80137;
    wire N__80136;
    wire N__80135;
    wire N__80132;
    wire N__80129;
    wire N__80128;
    wire N__80127;
    wire N__80124;
    wire N__80123;
    wire N__80122;
    wire N__80121;
    wire N__80120;
    wire N__80119;
    wire N__80116;
    wire N__80113;
    wire N__80112;
    wire N__80111;
    wire N__80106;
    wire N__80103;
    wire N__80102;
    wire N__80101;
    wire N__80100;
    wire N__80099;
    wire N__80098;
    wire N__80093;
    wire N__80088;
    wire N__80083;
    wire N__80082;
    wire N__80079;
    wire N__80074;
    wire N__80071;
    wire N__80068;
    wire N__80063;
    wire N__80058;
    wire N__80057;
    wire N__80054;
    wire N__80053;
    wire N__80052;
    wire N__80051;
    wire N__80048;
    wire N__80045;
    wire N__80042;
    wire N__80039;
    wire N__80036;
    wire N__80033;
    wire N__80028;
    wire N__80023;
    wire N__80018;
    wire N__80017;
    wire N__80016;
    wire N__80013;
    wire N__80010;
    wire N__80009;
    wire N__80008;
    wire N__80005;
    wire N__80002;
    wire N__79999;
    wire N__79998;
    wire N__79997;
    wire N__79994;
    wire N__79989;
    wire N__79984;
    wire N__79981;
    wire N__79978;
    wire N__79973;
    wire N__79970;
    wire N__79967;
    wire N__79962;
    wire N__79961;
    wire N__79960;
    wire N__79957;
    wire N__79954;
    wire N__79951;
    wire N__79948;
    wire N__79945;
    wire N__79942;
    wire N__79939;
    wire N__79932;
    wire N__79925;
    wire N__79918;
    wire N__79913;
    wire N__79906;
    wire N__79901;
    wire N__79890;
    wire N__79881;
    wire N__79880;
    wire N__79879;
    wire N__79878;
    wire N__79875;
    wire N__79872;
    wire N__79871;
    wire N__79870;
    wire N__79869;
    wire N__79868;
    wire N__79867;
    wire N__79866;
    wire N__79865;
    wire N__79864;
    wire N__79863;
    wire N__79862;
    wire N__79861;
    wire N__79860;
    wire N__79859;
    wire N__79856;
    wire N__79855;
    wire N__79854;
    wire N__79851;
    wire N__79850;
    wire N__79849;
    wire N__79848;
    wire N__79847;
    wire N__79846;
    wire N__79845;
    wire N__79844;
    wire N__79843;
    wire N__79842;
    wire N__79839;
    wire N__79838;
    wire N__79835;
    wire N__79834;
    wire N__79833;
    wire N__79830;
    wire N__79823;
    wire N__79822;
    wire N__79821;
    wire N__79820;
    wire N__79819;
    wire N__79818;
    wire N__79817;
    wire N__79816;
    wire N__79809;
    wire N__79808;
    wire N__79807;
    wire N__79794;
    wire N__79791;
    wire N__79786;
    wire N__79783;
    wire N__79776;
    wire N__79773;
    wire N__79770;
    wire N__79767;
    wire N__79764;
    wire N__79759;
    wire N__79756;
    wire N__79753;
    wire N__79750;
    wire N__79747;
    wire N__79744;
    wire N__79739;
    wire N__79734;
    wire N__79727;
    wire N__79722;
    wire N__79719;
    wire N__79714;
    wire N__79711;
    wire N__79702;
    wire N__79697;
    wire N__79692;
    wire N__79687;
    wire N__79684;
    wire N__79667;
    wire N__79664;
    wire N__79659;
    wire N__79654;
    wire N__79649;
    wire N__79646;
    wire N__79641;
    wire N__79632;
    wire N__79629;
    wire N__79628;
    wire N__79627;
    wire N__79624;
    wire N__79623;
    wire N__79620;
    wire N__79617;
    wire N__79614;
    wire N__79611;
    wire N__79608;
    wire N__79605;
    wire N__79600;
    wire N__79593;
    wire N__79590;
    wire N__79589;
    wire N__79586;
    wire N__79583;
    wire N__79578;
    wire N__79577;
    wire N__79576;
    wire N__79573;
    wire N__79570;
    wire N__79567;
    wire N__79564;
    wire N__79563;
    wire N__79560;
    wire N__79555;
    wire N__79552;
    wire N__79545;
    wire N__79544;
    wire N__79541;
    wire N__79538;
    wire N__79535;
    wire N__79532;
    wire N__79529;
    wire N__79526;
    wire N__79525;
    wire N__79522;
    wire N__79519;
    wire N__79516;
    wire N__79509;
    wire N__79508;
    wire N__79505;
    wire N__79502;
    wire N__79497;
    wire N__79494;
    wire N__79491;
    wire N__79488;
    wire N__79485;
    wire N__79484;
    wire N__79481;
    wire N__79478;
    wire N__79477;
    wire N__79476;
    wire N__79475;
    wire N__79470;
    wire N__79469;
    wire N__79464;
    wire N__79463;
    wire N__79460;
    wire N__79457;
    wire N__79454;
    wire N__79453;
    wire N__79452;
    wire N__79449;
    wire N__79446;
    wire N__79439;
    wire N__79434;
    wire N__79431;
    wire N__79422;
    wire N__79421;
    wire N__79420;
    wire N__79415;
    wire N__79412;
    wire N__79407;
    wire N__79404;
    wire N__79401;
    wire N__79398;
    wire N__79395;
    wire N__79394;
    wire N__79391;
    wire N__79388;
    wire N__79383;
    wire N__79380;
    wire N__79377;
    wire N__79374;
    wire N__79371;
    wire N__79368;
    wire N__79365;
    wire N__79362;
    wire N__79361;
    wire N__79360;
    wire N__79357;
    wire N__79354;
    wire N__79351;
    wire N__79344;
    wire N__79343;
    wire N__79342;
    wire N__79339;
    wire N__79336;
    wire N__79333;
    wire N__79326;
    wire N__79325;
    wire N__79324;
    wire N__79321;
    wire N__79318;
    wire N__79315;
    wire N__79312;
    wire N__79305;
    wire N__79304;
    wire N__79303;
    wire N__79300;
    wire N__79297;
    wire N__79294;
    wire N__79287;
    wire N__79286;
    wire N__79285;
    wire N__79282;
    wire N__79279;
    wire N__79276;
    wire N__79269;
    wire N__79266;
    wire N__79265;
    wire N__79264;
    wire N__79261;
    wire N__79258;
    wire N__79255;
    wire N__79248;
    wire N__79245;
    wire N__79244;
    wire N__79243;
    wire N__79240;
    wire N__79237;
    wire N__79234;
    wire N__79233;
    wire N__79230;
    wire N__79227;
    wire N__79226;
    wire N__79223;
    wire N__79222;
    wire N__79221;
    wire N__79218;
    wire N__79213;
    wire N__79210;
    wire N__79207;
    wire N__79202;
    wire N__79191;
    wire N__79190;
    wire N__79187;
    wire N__79184;
    wire N__79181;
    wire N__79180;
    wire N__79179;
    wire N__79176;
    wire N__79173;
    wire N__79170;
    wire N__79167;
    wire N__79162;
    wire N__79155;
    wire N__79154;
    wire N__79153;
    wire N__79152;
    wire N__79149;
    wire N__79148;
    wire N__79147;
    wire N__79146;
    wire N__79141;
    wire N__79138;
    wire N__79133;
    wire N__79130;
    wire N__79127;
    wire N__79124;
    wire N__79121;
    wire N__79118;
    wire N__79117;
    wire N__79114;
    wire N__79111;
    wire N__79108;
    wire N__79103;
    wire N__79100;
    wire N__79097;
    wire N__79092;
    wire N__79089;
    wire N__79080;
    wire N__79077;
    wire N__79074;
    wire N__79071;
    wire N__79070;
    wire N__79069;
    wire N__79066;
    wire N__79065;
    wire N__79064;
    wire N__79061;
    wire N__79060;
    wire N__79057;
    wire N__79054;
    wire N__79051;
    wire N__79048;
    wire N__79045;
    wire N__79042;
    wire N__79039;
    wire N__79036;
    wire N__79031;
    wire N__79030;
    wire N__79027;
    wire N__79018;
    wire N__79015;
    wire N__79012;
    wire N__79009;
    wire N__79002;
    wire N__78999;
    wire N__78996;
    wire N__78995;
    wire N__78992;
    wire N__78991;
    wire N__78990;
    wire N__78989;
    wire N__78988;
    wire N__78987;
    wire N__78986;
    wire N__78983;
    wire N__78982;
    wire N__78981;
    wire N__78980;
    wire N__78979;
    wire N__78978;
    wire N__78971;
    wire N__78966;
    wire N__78965;
    wire N__78964;
    wire N__78963;
    wire N__78962;
    wire N__78961;
    wire N__78958;
    wire N__78955;
    wire N__78952;
    wire N__78949;
    wire N__78948;
    wire N__78947;
    wire N__78946;
    wire N__78943;
    wire N__78940;
    wire N__78937;
    wire N__78934;
    wire N__78931;
    wire N__78928;
    wire N__78925;
    wire N__78922;
    wire N__78917;
    wire N__78916;
    wire N__78915;
    wire N__78914;
    wire N__78913;
    wire N__78910;
    wire N__78909;
    wire N__78908;
    wire N__78907;
    wire N__78900;
    wire N__78897;
    wire N__78894;
    wire N__78889;
    wire N__78886;
    wire N__78881;
    wire N__78874;
    wire N__78871;
    wire N__78866;
    wire N__78861;
    wire N__78858;
    wire N__78853;
    wire N__78852;
    wire N__78851;
    wire N__78848;
    wire N__78845;
    wire N__78842;
    wire N__78839;
    wire N__78834;
    wire N__78831;
    wire N__78828;
    wire N__78825;
    wire N__78822;
    wire N__78815;
    wire N__78812;
    wire N__78809;
    wire N__78808;
    wire N__78805;
    wire N__78802;
    wire N__78801;
    wire N__78798;
    wire N__78793;
    wire N__78788;
    wire N__78785;
    wire N__78778;
    wire N__78775;
    wire N__78770;
    wire N__78767;
    wire N__78764;
    wire N__78759;
    wire N__78752;
    wire N__78747;
    wire N__78742;
    wire N__78729;
    wire N__78726;
    wire N__78725;
    wire N__78724;
    wire N__78719;
    wire N__78716;
    wire N__78715;
    wire N__78710;
    wire N__78707;
    wire N__78706;
    wire N__78703;
    wire N__78698;
    wire N__78693;
    wire N__78690;
    wire N__78689;
    wire N__78686;
    wire N__78685;
    wire N__78682;
    wire N__78679;
    wire N__78676;
    wire N__78673;
    wire N__78670;
    wire N__78667;
    wire N__78664;
    wire N__78657;
    wire N__78656;
    wire N__78655;
    wire N__78654;
    wire N__78651;
    wire N__78642;
    wire N__78641;
    wire N__78640;
    wire N__78639;
    wire N__78638;
    wire N__78635;
    wire N__78632;
    wire N__78629;
    wire N__78628;
    wire N__78625;
    wire N__78622;
    wire N__78621;
    wire N__78620;
    wire N__78619;
    wire N__78612;
    wire N__78609;
    wire N__78604;
    wire N__78601;
    wire N__78596;
    wire N__78595;
    wire N__78594;
    wire N__78585;
    wire N__78582;
    wire N__78581;
    wire N__78576;
    wire N__78575;
    wire N__78574;
    wire N__78573;
    wire N__78572;
    wire N__78567;
    wire N__78564;
    wire N__78561;
    wire N__78560;
    wire N__78559;
    wire N__78558;
    wire N__78557;
    wire N__78556;
    wire N__78553;
    wire N__78550;
    wire N__78545;
    wire N__78540;
    wire N__78537;
    wire N__78536;
    wire N__78533;
    wire N__78528;
    wire N__78525;
    wire N__78522;
    wire N__78517;
    wire N__78516;
    wire N__78515;
    wire N__78512;
    wire N__78507;
    wire N__78506;
    wire N__78505;
    wire N__78504;
    wire N__78503;
    wire N__78500;
    wire N__78497;
    wire N__78494;
    wire N__78491;
    wire N__78486;
    wire N__78481;
    wire N__78478;
    wire N__78475;
    wire N__78470;
    wire N__78465;
    wire N__78458;
    wire N__78453;
    wire N__78448;
    wire N__78445;
    wire N__78432;
    wire N__78431;
    wire N__78430;
    wire N__78429;
    wire N__78426;
    wire N__78425;
    wire N__78424;
    wire N__78423;
    wire N__78422;
    wire N__78421;
    wire N__78418;
    wire N__78415;
    wire N__78410;
    wire N__78405;
    wire N__78400;
    wire N__78397;
    wire N__78394;
    wire N__78391;
    wire N__78388;
    wire N__78383;
    wire N__78380;
    wire N__78377;
    wire N__78370;
    wire N__78365;
    wire N__78360;
    wire N__78357;
    wire N__78356;
    wire N__78351;
    wire N__78350;
    wire N__78349;
    wire N__78346;
    wire N__78341;
    wire N__78336;
    wire N__78335;
    wire N__78334;
    wire N__78333;
    wire N__78332;
    wire N__78331;
    wire N__78328;
    wire N__78327;
    wire N__78326;
    wire N__78325;
    wire N__78322;
    wire N__78321;
    wire N__78320;
    wire N__78315;
    wire N__78312;
    wire N__78309;
    wire N__78306;
    wire N__78303;
    wire N__78300;
    wire N__78297;
    wire N__78296;
    wire N__78293;
    wire N__78290;
    wire N__78289;
    wire N__78288;
    wire N__78287;
    wire N__78286;
    wire N__78285;
    wire N__78282;
    wire N__78279;
    wire N__78276;
    wire N__78271;
    wire N__78270;
    wire N__78267;
    wire N__78264;
    wire N__78261;
    wire N__78260;
    wire N__78259;
    wire N__78256;
    wire N__78255;
    wire N__78252;
    wire N__78249;
    wire N__78246;
    wire N__78241;
    wire N__78240;
    wire N__78235;
    wire N__78232;
    wire N__78225;
    wire N__78222;
    wire N__78221;
    wire N__78220;
    wire N__78219;
    wire N__78216;
    wire N__78211;
    wire N__78210;
    wire N__78209;
    wire N__78208;
    wire N__78207;
    wire N__78204;
    wire N__78201;
    wire N__78198;
    wire N__78195;
    wire N__78190;
    wire N__78187;
    wire N__78184;
    wire N__78181;
    wire N__78176;
    wire N__78171;
    wire N__78168;
    wire N__78167;
    wire N__78166;
    wire N__78163;
    wire N__78160;
    wire N__78155;
    wire N__78152;
    wire N__78145;
    wire N__78140;
    wire N__78139;
    wire N__78136;
    wire N__78131;
    wire N__78124;
    wire N__78119;
    wire N__78116;
    wire N__78111;
    wire N__78104;
    wire N__78097;
    wire N__78094;
    wire N__78091;
    wire N__78088;
    wire N__78083;
    wire N__78076;
    wire N__78073;
    wire N__78060;
    wire N__78057;
    wire N__78054;
    wire N__78051;
    wire N__78048;
    wire N__78045;
    wire N__78042;
    wire N__78039;
    wire N__78038;
    wire N__78037;
    wire N__78036;
    wire N__78035;
    wire N__78032;
    wire N__78029;
    wire N__78026;
    wire N__78025;
    wire N__78024;
    wire N__78021;
    wire N__78020;
    wire N__78017;
    wire N__78012;
    wire N__78009;
    wire N__78004;
    wire N__78001;
    wire N__77998;
    wire N__77995;
    wire N__77992;
    wire N__77985;
    wire N__77976;
    wire N__77973;
    wire N__77970;
    wire N__77967;
    wire N__77964;
    wire N__77961;
    wire N__77958;
    wire N__77955;
    wire N__77952;
    wire N__77949;
    wire N__77948;
    wire N__77947;
    wire N__77944;
    wire N__77943;
    wire N__77940;
    wire N__77937;
    wire N__77936;
    wire N__77933;
    wire N__77930;
    wire N__77925;
    wire N__77922;
    wire N__77919;
    wire N__77916;
    wire N__77913;
    wire N__77904;
    wire N__77903;
    wire N__77902;
    wire N__77901;
    wire N__77896;
    wire N__77893;
    wire N__77890;
    wire N__77883;
    wire N__77880;
    wire N__77877;
    wire N__77874;
    wire N__77873;
    wire N__77870;
    wire N__77867;
    wire N__77866;
    wire N__77863;
    wire N__77860;
    wire N__77857;
    wire N__77856;
    wire N__77853;
    wire N__77850;
    wire N__77847;
    wire N__77844;
    wire N__77841;
    wire N__77838;
    wire N__77835;
    wire N__77826;
    wire N__77825;
    wire N__77822;
    wire N__77821;
    wire N__77820;
    wire N__77819;
    wire N__77816;
    wire N__77813;
    wire N__77810;
    wire N__77807;
    wire N__77804;
    wire N__77801;
    wire N__77798;
    wire N__77795;
    wire N__77792;
    wire N__77781;
    wire N__77778;
    wire N__77775;
    wire N__77772;
    wire N__77769;
    wire N__77766;
    wire N__77763;
    wire N__77760;
    wire N__77759;
    wire N__77756;
    wire N__77753;
    wire N__77750;
    wire N__77747;
    wire N__77744;
    wire N__77741;
    wire N__77736;
    wire N__77733;
    wire N__77732;
    wire N__77731;
    wire N__77728;
    wire N__77723;
    wire N__77718;
    wire N__77715;
    wire N__77712;
    wire N__77711;
    wire N__77706;
    wire N__77703;
    wire N__77700;
    wire N__77699;
    wire N__77696;
    wire N__77693;
    wire N__77692;
    wire N__77691;
    wire N__77688;
    wire N__77685;
    wire N__77682;
    wire N__77679;
    wire N__77678;
    wire N__77677;
    wire N__77676;
    wire N__77673;
    wire N__77670;
    wire N__77667;
    wire N__77664;
    wire N__77659;
    wire N__77656;
    wire N__77651;
    wire N__77648;
    wire N__77645;
    wire N__77642;
    wire N__77631;
    wire N__77630;
    wire N__77629;
    wire N__77628;
    wire N__77627;
    wire N__77626;
    wire N__77623;
    wire N__77620;
    wire N__77619;
    wire N__77618;
    wire N__77613;
    wire N__77610;
    wire N__77607;
    wire N__77604;
    wire N__77601;
    wire N__77596;
    wire N__77593;
    wire N__77588;
    wire N__77585;
    wire N__77582;
    wire N__77579;
    wire N__77576;
    wire N__77573;
    wire N__77568;
    wire N__77559;
    wire N__77558;
    wire N__77555;
    wire N__77554;
    wire N__77553;
    wire N__77550;
    wire N__77547;
    wire N__77544;
    wire N__77543;
    wire N__77542;
    wire N__77539;
    wire N__77536;
    wire N__77533;
    wire N__77530;
    wire N__77525;
    wire N__77522;
    wire N__77519;
    wire N__77508;
    wire N__77505;
    wire N__77504;
    wire N__77501;
    wire N__77500;
    wire N__77499;
    wire N__77496;
    wire N__77493;
    wire N__77490;
    wire N__77489;
    wire N__77486;
    wire N__77483;
    wire N__77478;
    wire N__77475;
    wire N__77472;
    wire N__77467;
    wire N__77460;
    wire N__77457;
    wire N__77454;
    wire N__77453;
    wire N__77450;
    wire N__77447;
    wire N__77444;
    wire N__77441;
    wire N__77436;
    wire N__77435;
    wire N__77432;
    wire N__77429;
    wire N__77428;
    wire N__77427;
    wire N__77424;
    wire N__77421;
    wire N__77416;
    wire N__77409;
    wire N__77408;
    wire N__77405;
    wire N__77402;
    wire N__77399;
    wire N__77394;
    wire N__77391;
    wire N__77390;
    wire N__77389;
    wire N__77382;
    wire N__77379;
    wire N__77376;
    wire N__77373;
    wire N__77370;
    wire N__77367;
    wire N__77366;
    wire N__77363;
    wire N__77360;
    wire N__77357;
    wire N__77352;
    wire N__77351;
    wire N__77348;
    wire N__77345;
    wire N__77344;
    wire N__77343;
    wire N__77340;
    wire N__77337;
    wire N__77336;
    wire N__77333;
    wire N__77330;
    wire N__77325;
    wire N__77322;
    wire N__77313;
    wire N__77312;
    wire N__77307;
    wire N__77304;
    wire N__77301;
    wire N__77298;
    wire N__77295;
    wire N__77294;
    wire N__77291;
    wire N__77288;
    wire N__77287;
    wire N__77286;
    wire N__77285;
    wire N__77282;
    wire N__77281;
    wire N__77278;
    wire N__77273;
    wire N__77272;
    wire N__77269;
    wire N__77266;
    wire N__77263;
    wire N__77260;
    wire N__77257;
    wire N__77254;
    wire N__77241;
    wire N__77238;
    wire N__77235;
    wire N__77232;
    wire N__77229;
    wire N__77226;
    wire N__77223;
    wire N__77220;
    wire N__77217;
    wire N__77214;
    wire N__77211;
    wire N__77210;
    wire N__77207;
    wire N__77204;
    wire N__77203;
    wire N__77202;
    wire N__77197;
    wire N__77194;
    wire N__77191;
    wire N__77186;
    wire N__77185;
    wire N__77184;
    wire N__77181;
    wire N__77178;
    wire N__77175;
    wire N__77172;
    wire N__77169;
    wire N__77166;
    wire N__77157;
    wire N__77154;
    wire N__77151;
    wire N__77148;
    wire N__77145;
    wire N__77142;
    wire N__77141;
    wire N__77138;
    wire N__77135;
    wire N__77132;
    wire N__77129;
    wire N__77128;
    wire N__77125;
    wire N__77122;
    wire N__77121;
    wire N__77118;
    wire N__77113;
    wire N__77110;
    wire N__77103;
    wire N__77100;
    wire N__77097;
    wire N__77096;
    wire N__77095;
    wire N__77094;
    wire N__77091;
    wire N__77084;
    wire N__77083;
    wire N__77082;
    wire N__77081;
    wire N__77076;
    wire N__77073;
    wire N__77068;
    wire N__77065;
    wire N__77058;
    wire N__77055;
    wire N__77052;
    wire N__77049;
    wire N__77048;
    wire N__77047;
    wire N__77046;
    wire N__77043;
    wire N__77036;
    wire N__77031;
    wire N__77030;
    wire N__77027;
    wire N__77026;
    wire N__77025;
    wire N__77022;
    wire N__77021;
    wire N__77020;
    wire N__77017;
    wire N__77014;
    wire N__77011;
    wire N__77004;
    wire N__76995;
    wire N__76994;
    wire N__76993;
    wire N__76992;
    wire N__76991;
    wire N__76990;
    wire N__76985;
    wire N__76982;
    wire N__76981;
    wire N__76980;
    wire N__76979;
    wire N__76976;
    wire N__76971;
    wire N__76968;
    wire N__76965;
    wire N__76958;
    wire N__76955;
    wire N__76952;
    wire N__76945;
    wire N__76942;
    wire N__76937;
    wire N__76932;
    wire N__76929;
    wire N__76926;
    wire N__76923;
    wire N__76920;
    wire N__76917;
    wire N__76914;
    wire N__76911;
    wire N__76910;
    wire N__76907;
    wire N__76906;
    wire N__76905;
    wire N__76904;
    wire N__76901;
    wire N__76898;
    wire N__76895;
    wire N__76890;
    wire N__76889;
    wire N__76886;
    wire N__76881;
    wire N__76878;
    wire N__76875;
    wire N__76870;
    wire N__76867;
    wire N__76860;
    wire N__76857;
    wire N__76856;
    wire N__76855;
    wire N__76852;
    wire N__76847;
    wire N__76846;
    wire N__76843;
    wire N__76840;
    wire N__76839;
    wire N__76836;
    wire N__76831;
    wire N__76828;
    wire N__76825;
    wire N__76822;
    wire N__76815;
    wire N__76812;
    wire N__76809;
    wire N__76808;
    wire N__76807;
    wire N__76804;
    wire N__76801;
    wire N__76798;
    wire N__76795;
    wire N__76792;
    wire N__76791;
    wire N__76790;
    wire N__76789;
    wire N__76788;
    wire N__76785;
    wire N__76782;
    wire N__76779;
    wire N__76776;
    wire N__76773;
    wire N__76768;
    wire N__76765;
    wire N__76752;
    wire N__76751;
    wire N__76750;
    wire N__76747;
    wire N__76746;
    wire N__76743;
    wire N__76740;
    wire N__76739;
    wire N__76738;
    wire N__76735;
    wire N__76732;
    wire N__76729;
    wire N__76726;
    wire N__76723;
    wire N__76720;
    wire N__76717;
    wire N__76714;
    wire N__76713;
    wire N__76710;
    wire N__76707;
    wire N__76702;
    wire N__76697;
    wire N__76694;
    wire N__76691;
    wire N__76684;
    wire N__76677;
    wire N__76674;
    wire N__76673;
    wire N__76670;
    wire N__76667;
    wire N__76662;
    wire N__76659;
    wire N__76656;
    wire N__76653;
    wire N__76652;
    wire N__76651;
    wire N__76648;
    wire N__76645;
    wire N__76644;
    wire N__76641;
    wire N__76636;
    wire N__76635;
    wire N__76632;
    wire N__76629;
    wire N__76626;
    wire N__76623;
    wire N__76614;
    wire N__76611;
    wire N__76608;
    wire N__76605;
    wire N__76602;
    wire N__76599;
    wire N__76596;
    wire N__76593;
    wire N__76590;
    wire N__76589;
    wire N__76586;
    wire N__76585;
    wire N__76584;
    wire N__76583;
    wire N__76580;
    wire N__76579;
    wire N__76576;
    wire N__76573;
    wire N__76572;
    wire N__76569;
    wire N__76566;
    wire N__76565;
    wire N__76564;
    wire N__76563;
    wire N__76562;
    wire N__76561;
    wire N__76558;
    wire N__76555;
    wire N__76552;
    wire N__76549;
    wire N__76546;
    wire N__76545;
    wire N__76544;
    wire N__76543;
    wire N__76542;
    wire N__76541;
    wire N__76540;
    wire N__76537;
    wire N__76532;
    wire N__76529;
    wire N__76524;
    wire N__76523;
    wire N__76522;
    wire N__76521;
    wire N__76520;
    wire N__76517;
    wire N__76508;
    wire N__76505;
    wire N__76500;
    wire N__76497;
    wire N__76490;
    wire N__76483;
    wire N__76482;
    wire N__76481;
    wire N__76480;
    wire N__76479;
    wire N__76478;
    wire N__76477;
    wire N__76476;
    wire N__76475;
    wire N__76474;
    wire N__76473;
    wire N__76470;
    wire N__76467;
    wire N__76462;
    wire N__76459;
    wire N__76452;
    wire N__76447;
    wire N__76442;
    wire N__76439;
    wire N__76436;
    wire N__76433;
    wire N__76430;
    wire N__76423;
    wire N__76420;
    wire N__76415;
    wire N__76410;
    wire N__76405;
    wire N__76402;
    wire N__76397;
    wire N__76380;
    wire N__76375;
    wire N__76372;
    wire N__76369;
    wire N__76366;
    wire N__76363;
    wire N__76356;
    wire N__76353;
    wire N__76352;
    wire N__76349;
    wire N__76346;
    wire N__76341;
    wire N__76338;
    wire N__76335;
    wire N__76334;
    wire N__76331;
    wire N__76328;
    wire N__76325;
    wire N__76322;
    wire N__76319;
    wire N__76314;
    wire N__76311;
    wire N__76308;
    wire N__76305;
    wire N__76302;
    wire N__76301;
    wire N__76298;
    wire N__76295;
    wire N__76290;
    wire N__76287;
    wire N__76284;
    wire N__76281;
    wire N__76278;
    wire N__76275;
    wire N__76272;
    wire N__76269;
    wire N__76266;
    wire N__76263;
    wire N__76262;
    wire N__76261;
    wire N__76258;
    wire N__76255;
    wire N__76252;
    wire N__76247;
    wire N__76244;
    wire N__76239;
    wire N__76236;
    wire N__76235;
    wire N__76232;
    wire N__76229;
    wire N__76224;
    wire N__76221;
    wire N__76218;
    wire N__76215;
    wire N__76214;
    wire N__76211;
    wire N__76208;
    wire N__76205;
    wire N__76202;
    wire N__76197;
    wire N__76194;
    wire N__76191;
    wire N__76190;
    wire N__76187;
    wire N__76184;
    wire N__76181;
    wire N__76176;
    wire N__76175;
    wire N__76172;
    wire N__76169;
    wire N__76166;
    wire N__76161;
    wire N__76158;
    wire N__76155;
    wire N__76152;
    wire N__76149;
    wire N__76146;
    wire N__76145;
    wire N__76144;
    wire N__76143;
    wire N__76142;
    wire N__76139;
    wire N__76134;
    wire N__76131;
    wire N__76128;
    wire N__76123;
    wire N__76122;
    wire N__76119;
    wire N__76116;
    wire N__76113;
    wire N__76110;
    wire N__76101;
    wire N__76100;
    wire N__76097;
    wire N__76096;
    wire N__76091;
    wire N__76090;
    wire N__76087;
    wire N__76084;
    wire N__76083;
    wire N__76082;
    wire N__76079;
    wire N__76076;
    wire N__76073;
    wire N__76068;
    wire N__76059;
    wire N__76058;
    wire N__76055;
    wire N__76054;
    wire N__76051;
    wire N__76050;
    wire N__76047;
    wire N__76044;
    wire N__76043;
    wire N__76040;
    wire N__76037;
    wire N__76034;
    wire N__76031;
    wire N__76028;
    wire N__76025;
    wire N__76014;
    wire N__76011;
    wire N__76008;
    wire N__76005;
    wire N__76002;
    wire N__75999;
    wire N__75996;
    wire N__75993;
    wire N__75990;
    wire N__75987;
    wire N__75984;
    wire N__75981;
    wire N__75978;
    wire N__75975;
    wire N__75972;
    wire N__75969;
    wire N__75966;
    wire N__75963;
    wire N__75960;
    wire N__75957;
    wire N__75954;
    wire N__75951;
    wire N__75948;
    wire N__75945;
    wire N__75944;
    wire N__75943;
    wire N__75940;
    wire N__75937;
    wire N__75934;
    wire N__75931;
    wire N__75930;
    wire N__75927;
    wire N__75924;
    wire N__75923;
    wire N__75922;
    wire N__75919;
    wire N__75916;
    wire N__75913;
    wire N__75910;
    wire N__75905;
    wire N__75902;
    wire N__75895;
    wire N__75892;
    wire N__75885;
    wire N__75882;
    wire N__75879;
    wire N__75876;
    wire N__75875;
    wire N__75874;
    wire N__75873;
    wire N__75870;
    wire N__75867;
    wire N__75864;
    wire N__75863;
    wire N__75860;
    wire N__75857;
    wire N__75854;
    wire N__75851;
    wire N__75848;
    wire N__75837;
    wire N__75836;
    wire N__75833;
    wire N__75830;
    wire N__75827;
    wire N__75826;
    wire N__75825;
    wire N__75824;
    wire N__75819;
    wire N__75816;
    wire N__75813;
    wire N__75810;
    wire N__75807;
    wire N__75804;
    wire N__75795;
    wire N__75794;
    wire N__75793;
    wire N__75792;
    wire N__75791;
    wire N__75790;
    wire N__75787;
    wire N__75784;
    wire N__75781;
    wire N__75778;
    wire N__75775;
    wire N__75772;
    wire N__75767;
    wire N__75758;
    wire N__75753;
    wire N__75750;
    wire N__75747;
    wire N__75746;
    wire N__75745;
    wire N__75744;
    wire N__75741;
    wire N__75738;
    wire N__75737;
    wire N__75736;
    wire N__75735;
    wire N__75732;
    wire N__75729;
    wire N__75724;
    wire N__75721;
    wire N__75718;
    wire N__75715;
    wire N__75714;
    wire N__75709;
    wire N__75706;
    wire N__75697;
    wire N__75690;
    wire N__75687;
    wire N__75684;
    wire N__75683;
    wire N__75678;
    wire N__75675;
    wire N__75672;
    wire N__75669;
    wire N__75666;
    wire N__75663;
    wire N__75660;
    wire N__75657;
    wire N__75654;
    wire N__75651;
    wire N__75648;
    wire N__75645;
    wire N__75642;
    wire N__75639;
    wire N__75636;
    wire N__75633;
    wire N__75630;
    wire N__75627;
    wire N__75624;
    wire N__75621;
    wire N__75618;
    wire N__75615;
    wire N__75614;
    wire N__75613;
    wire N__75610;
    wire N__75607;
    wire N__75604;
    wire N__75597;
    wire N__75594;
    wire N__75591;
    wire N__75588;
    wire N__75585;
    wire N__75582;
    wire N__75579;
    wire N__75576;
    wire N__75573;
    wire N__75570;
    wire N__75569;
    wire N__75568;
    wire N__75567;
    wire N__75566;
    wire N__75565;
    wire N__75562;
    wire N__75559;
    wire N__75556;
    wire N__75553;
    wire N__75550;
    wire N__75547;
    wire N__75542;
    wire N__75533;
    wire N__75528;
    wire N__75527;
    wire N__75526;
    wire N__75523;
    wire N__75520;
    wire N__75517;
    wire N__75514;
    wire N__75507;
    wire N__75504;
    wire N__75503;
    wire N__75500;
    wire N__75499;
    wire N__75496;
    wire N__75493;
    wire N__75490;
    wire N__75483;
    wire N__75480;
    wire N__75479;
    wire N__75478;
    wire N__75475;
    wire N__75472;
    wire N__75469;
    wire N__75462;
    wire N__75459;
    wire N__75458;
    wire N__75457;
    wire N__75454;
    wire N__75451;
    wire N__75448;
    wire N__75441;
    wire N__75438;
    wire N__75437;
    wire N__75436;
    wire N__75433;
    wire N__75430;
    wire N__75427;
    wire N__75420;
    wire N__75417;
    wire N__75416;
    wire N__75415;
    wire N__75412;
    wire N__75409;
    wire N__75406;
    wire N__75399;
    wire N__75396;
    wire N__75393;
    wire N__75392;
    wire N__75391;
    wire N__75388;
    wire N__75385;
    wire N__75380;
    wire N__75377;
    wire N__75372;
    wire N__75371;
    wire N__75370;
    wire N__75369;
    wire N__75366;
    wire N__75365;
    wire N__75364;
    wire N__75363;
    wire N__75362;
    wire N__75361;
    wire N__75360;
    wire N__75359;
    wire N__75358;
    wire N__75355;
    wire N__75352;
    wire N__75351;
    wire N__75348;
    wire N__75345;
    wire N__75344;
    wire N__75343;
    wire N__75340;
    wire N__75339;
    wire N__75336;
    wire N__75335;
    wire N__75330;
    wire N__75327;
    wire N__75326;
    wire N__75325;
    wire N__75324;
    wire N__75321;
    wire N__75320;
    wire N__75319;
    wire N__75318;
    wire N__75317;
    wire N__75316;
    wire N__75311;
    wire N__75306;
    wire N__75303;
    wire N__75300;
    wire N__75297;
    wire N__75296;
    wire N__75293;
    wire N__75290;
    wire N__75289;
    wire N__75286;
    wire N__75283;
    wire N__75280;
    wire N__75277;
    wire N__75274;
    wire N__75271;
    wire N__75270;
    wire N__75269;
    wire N__75266;
    wire N__75263;
    wire N__75260;
    wire N__75257;
    wire N__75254;
    wire N__75249;
    wire N__75244;
    wire N__75241;
    wire N__75238;
    wire N__75231;
    wire N__75230;
    wire N__75229;
    wire N__75224;
    wire N__75221;
    wire N__75218;
    wire N__75213;
    wire N__75210;
    wire N__75203;
    wire N__75202;
    wire N__75197;
    wire N__75194;
    wire N__75191;
    wire N__75186;
    wire N__75173;
    wire N__75170;
    wire N__75167;
    wire N__75164;
    wire N__75161;
    wire N__75156;
    wire N__75151;
    wire N__75148;
    wire N__75145;
    wire N__75136;
    wire N__75125;
    wire N__75122;
    wire N__75111;
    wire N__75110;
    wire N__75107;
    wire N__75106;
    wire N__75103;
    wire N__75098;
    wire N__75093;
    wire N__75090;
    wire N__75089;
    wire N__75088;
    wire N__75087;
    wire N__75086;
    wire N__75085;
    wire N__75084;
    wire N__75083;
    wire N__75080;
    wire N__75079;
    wire N__75076;
    wire N__75073;
    wire N__75072;
    wire N__75067;
    wire N__75066;
    wire N__75063;
    wire N__75062;
    wire N__75061;
    wire N__75058;
    wire N__75055;
    wire N__75054;
    wire N__75053;
    wire N__75052;
    wire N__75051;
    wire N__75050;
    wire N__75049;
    wire N__75048;
    wire N__75045;
    wire N__75042;
    wire N__75039;
    wire N__75036;
    wire N__75033;
    wire N__75030;
    wire N__75027;
    wire N__75024;
    wire N__75021;
    wire N__75018;
    wire N__75015;
    wire N__75012;
    wire N__75011;
    wire N__75010;
    wire N__75009;
    wire N__75008;
    wire N__75005;
    wire N__75002;
    wire N__74999;
    wire N__74996;
    wire N__74993;
    wire N__74992;
    wire N__74987;
    wire N__74982;
    wire N__74975;
    wire N__74972;
    wire N__74965;
    wire N__74962;
    wire N__74959;
    wire N__74956;
    wire N__74953;
    wire N__74950;
    wire N__74949;
    wire N__74948;
    wire N__74947;
    wire N__74946;
    wire N__74943;
    wire N__74940;
    wire N__74937;
    wire N__74934;
    wire N__74931;
    wire N__74928;
    wire N__74925;
    wire N__74922;
    wire N__74917;
    wire N__74912;
    wire N__74909;
    wire N__74904;
    wire N__74901;
    wire N__74896;
    wire N__74895;
    wire N__74894;
    wire N__74893;
    wire N__74890;
    wire N__74887;
    wire N__74882;
    wire N__74877;
    wire N__74874;
    wire N__74871;
    wire N__74864;
    wire N__74855;
    wire N__74848;
    wire N__74843;
    wire N__74840;
    wire N__74825;
    wire N__74822;
    wire N__74819;
    wire N__74808;
    wire N__74807;
    wire N__74806;
    wire N__74803;
    wire N__74800;
    wire N__74797;
    wire N__74794;
    wire N__74791;
    wire N__74790;
    wire N__74787;
    wire N__74782;
    wire N__74779;
    wire N__74776;
    wire N__74771;
    wire N__74768;
    wire N__74765;
    wire N__74760;
    wire N__74759;
    wire N__74756;
    wire N__74753;
    wire N__74752;
    wire N__74749;
    wire N__74744;
    wire N__74741;
    wire N__74736;
    wire N__74733;
    wire N__74730;
    wire N__74727;
    wire N__74726;
    wire N__74725;
    wire N__74722;
    wire N__74719;
    wire N__74716;
    wire N__74715;
    wire N__74714;
    wire N__74709;
    wire N__74706;
    wire N__74703;
    wire N__74700;
    wire N__74693;
    wire N__74690;
    wire N__74687;
    wire N__74684;
    wire N__74681;
    wire N__74678;
    wire N__74673;
    wire N__74670;
    wire N__74667;
    wire N__74666;
    wire N__74663;
    wire N__74660;
    wire N__74659;
    wire N__74654;
    wire N__74651;
    wire N__74646;
    wire N__74645;
    wire N__74642;
    wire N__74639;
    wire N__74638;
    wire N__74633;
    wire N__74630;
    wire N__74625;
    wire N__74624;
    wire N__74623;
    wire N__74620;
    wire N__74617;
    wire N__74614;
    wire N__74609;
    wire N__74606;
    wire N__74601;
    wire N__74598;
    wire N__74597;
    wire N__74594;
    wire N__74591;
    wire N__74590;
    wire N__74587;
    wire N__74584;
    wire N__74581;
    wire N__74574;
    wire N__74571;
    wire N__74568;
    wire N__74565;
    wire N__74564;
    wire N__74561;
    wire N__74558;
    wire N__74555;
    wire N__74550;
    wire N__74549;
    wire N__74544;
    wire N__74543;
    wire N__74540;
    wire N__74537;
    wire N__74534;
    wire N__74531;
    wire N__74528;
    wire N__74523;
    wire N__74522;
    wire N__74519;
    wire N__74516;
    wire N__74515;
    wire N__74512;
    wire N__74509;
    wire N__74506;
    wire N__74499;
    wire N__74496;
    wire N__74493;
    wire N__74492;
    wire N__74489;
    wire N__74486;
    wire N__74483;
    wire N__74480;
    wire N__74475;
    wire N__74474;
    wire N__74471;
    wire N__74468;
    wire N__74465;
    wire N__74462;
    wire N__74457;
    wire N__74456;
    wire N__74455;
    wire N__74454;
    wire N__74453;
    wire N__74450;
    wire N__74449;
    wire N__74446;
    wire N__74445;
    wire N__74442;
    wire N__74441;
    wire N__74436;
    wire N__74433;
    wire N__74428;
    wire N__74425;
    wire N__74420;
    wire N__74417;
    wire N__74414;
    wire N__74411;
    wire N__74408;
    wire N__74403;
    wire N__74400;
    wire N__74397;
    wire N__74394;
    wire N__74391;
    wire N__74390;
    wire N__74387;
    wire N__74380;
    wire N__74377;
    wire N__74370;
    wire N__74367;
    wire N__74366;
    wire N__74363;
    wire N__74360;
    wire N__74355;
    wire N__74354;
    wire N__74351;
    wire N__74348;
    wire N__74347;
    wire N__74346;
    wire N__74345;
    wire N__74342;
    wire N__74341;
    wire N__74340;
    wire N__74337;
    wire N__74330;
    wire N__74327;
    wire N__74322;
    wire N__74319;
    wire N__74316;
    wire N__74315;
    wire N__74310;
    wire N__74307;
    wire N__74304;
    wire N__74301;
    wire N__74292;
    wire N__74291;
    wire N__74290;
    wire N__74287;
    wire N__74286;
    wire N__74283;
    wire N__74280;
    wire N__74279;
    wire N__74274;
    wire N__74273;
    wire N__74270;
    wire N__74267;
    wire N__74264;
    wire N__74263;
    wire N__74260;
    wire N__74257;
    wire N__74252;
    wire N__74247;
    wire N__74246;
    wire N__74237;
    wire N__74234;
    wire N__74231;
    wire N__74226;
    wire N__74225;
    wire N__74222;
    wire N__74219;
    wire N__74218;
    wire N__74215;
    wire N__74212;
    wire N__74209;
    wire N__74204;
    wire N__74201;
    wire N__74198;
    wire N__74195;
    wire N__74192;
    wire N__74187;
    wire N__74184;
    wire N__74181;
    wire N__74178;
    wire N__74175;
    wire N__74174;
    wire N__74173;
    wire N__74168;
    wire N__74165;
    wire N__74162;
    wire N__74157;
    wire N__74156;
    wire N__74153;
    wire N__74152;
    wire N__74151;
    wire N__74148;
    wire N__74145;
    wire N__74142;
    wire N__74139;
    wire N__74136;
    wire N__74127;
    wire N__74124;
    wire N__74123;
    wire N__74120;
    wire N__74119;
    wire N__74116;
    wire N__74113;
    wire N__74110;
    wire N__74107;
    wire N__74104;
    wire N__74101;
    wire N__74094;
    wire N__74093;
    wire N__74092;
    wire N__74089;
    wire N__74086;
    wire N__74083;
    wire N__74080;
    wire N__74077;
    wire N__74074;
    wire N__74069;
    wire N__74066;
    wire N__74061;
    wire N__74060;
    wire N__74057;
    wire N__74054;
    wire N__74051;
    wire N__74046;
    wire N__74043;
    wire N__74042;
    wire N__74039;
    wire N__74038;
    wire N__74035;
    wire N__74030;
    wire N__74025;
    wire N__74022;
    wire N__74019;
    wire N__74018;
    wire N__74013;
    wire N__74010;
    wire N__74007;
    wire N__74004;
    wire N__74001;
    wire N__74000;
    wire N__73997;
    wire N__73994;
    wire N__73991;
    wire N__73988;
    wire N__73985;
    wire N__73980;
    wire N__73979;
    wire N__73978;
    wire N__73977;
    wire N__73974;
    wire N__73967;
    wire N__73964;
    wire N__73961;
    wire N__73958;
    wire N__73955;
    wire N__73950;
    wire N__73949;
    wire N__73948;
    wire N__73947;
    wire N__73946;
    wire N__73943;
    wire N__73942;
    wire N__73941;
    wire N__73938;
    wire N__73937;
    wire N__73936;
    wire N__73935;
    wire N__73934;
    wire N__73931;
    wire N__73930;
    wire N__73929;
    wire N__73928;
    wire N__73927;
    wire N__73926;
    wire N__73923;
    wire N__73922;
    wire N__73921;
    wire N__73920;
    wire N__73915;
    wire N__73914;
    wire N__73911;
    wire N__73910;
    wire N__73909;
    wire N__73908;
    wire N__73907;
    wire N__73906;
    wire N__73903;
    wire N__73898;
    wire N__73893;
    wire N__73890;
    wire N__73887;
    wire N__73884;
    wire N__73881;
    wire N__73880;
    wire N__73879;
    wire N__73878;
    wire N__73875;
    wire N__73872;
    wire N__73869;
    wire N__73864;
    wire N__73861;
    wire N__73858;
    wire N__73855;
    wire N__73852;
    wire N__73849;
    wire N__73848;
    wire N__73847;
    wire N__73844;
    wire N__73841;
    wire N__73834;
    wire N__73829;
    wire N__73826;
    wire N__73823;
    wire N__73818;
    wire N__73817;
    wire N__73808;
    wire N__73805;
    wire N__73802;
    wire N__73799;
    wire N__73796;
    wire N__73793;
    wire N__73788;
    wire N__73785;
    wire N__73782;
    wire N__73781;
    wire N__73778;
    wire N__73773;
    wire N__73768;
    wire N__73765;
    wire N__73760;
    wire N__73757;
    wire N__73754;
    wire N__73747;
    wire N__73742;
    wire N__73737;
    wire N__73732;
    wire N__73729;
    wire N__73726;
    wire N__73723;
    wire N__73714;
    wire N__73707;
    wire N__73702;
    wire N__73689;
    wire N__73688;
    wire N__73685;
    wire N__73682;
    wire N__73679;
    wire N__73674;
    wire N__73673;
    wire N__73672;
    wire N__73671;
    wire N__73668;
    wire N__73665;
    wire N__73662;
    wire N__73659;
    wire N__73656;
    wire N__73655;
    wire N__73652;
    wire N__73647;
    wire N__73644;
    wire N__73641;
    wire N__73640;
    wire N__73639;
    wire N__73638;
    wire N__73637;
    wire N__73636;
    wire N__73635;
    wire N__73634;
    wire N__73633;
    wire N__73626;
    wire N__73625;
    wire N__73624;
    wire N__73623;
    wire N__73622;
    wire N__73621;
    wire N__73618;
    wire N__73617;
    wire N__73616;
    wire N__73613;
    wire N__73606;
    wire N__73601;
    wire N__73598;
    wire N__73597;
    wire N__73596;
    wire N__73595;
    wire N__73594;
    wire N__73593;
    wire N__73590;
    wire N__73587;
    wire N__73584;
    wire N__73581;
    wire N__73578;
    wire N__73577;
    wire N__73574;
    wire N__73571;
    wire N__73568;
    wire N__73565;
    wire N__73562;
    wire N__73559;
    wire N__73556;
    wire N__73551;
    wire N__73546;
    wire N__73545;
    wire N__73540;
    wire N__73535;
    wire N__73528;
    wire N__73525;
    wire N__73524;
    wire N__73523;
    wire N__73522;
    wire N__73519;
    wire N__73518;
    wire N__73515;
    wire N__73508;
    wire N__73501;
    wire N__73498;
    wire N__73495;
    wire N__73492;
    wire N__73487;
    wire N__73484;
    wire N__73481;
    wire N__73480;
    wire N__73477;
    wire N__73474;
    wire N__73471;
    wire N__73468;
    wire N__73465;
    wire N__73460;
    wire N__73455;
    wire N__73452;
    wire N__73449;
    wire N__73442;
    wire N__73439;
    wire N__73434;
    wire N__73429;
    wire N__73420;
    wire N__73415;
    wire N__73404;
    wire N__73403;
    wire N__73400;
    wire N__73399;
    wire N__73396;
    wire N__73393;
    wire N__73390;
    wire N__73387;
    wire N__73382;
    wire N__73379;
    wire N__73376;
    wire N__73371;
    wire N__73368;
    wire N__73367;
    wire N__73364;
    wire N__73361;
    wire N__73358;
    wire N__73353;
    wire N__73352;
    wire N__73351;
    wire N__73348;
    wire N__73347;
    wire N__73344;
    wire N__73341;
    wire N__73338;
    wire N__73335;
    wire N__73326;
    wire N__73323;
    wire N__73322;
    wire N__73321;
    wire N__73318;
    wire N__73313;
    wire N__73312;
    wire N__73307;
    wire N__73304;
    wire N__73299;
    wire N__73298;
    wire N__73293;
    wire N__73292;
    wire N__73291;
    wire N__73288;
    wire N__73285;
    wire N__73282;
    wire N__73279;
    wire N__73274;
    wire N__73269;
    wire N__73268;
    wire N__73265;
    wire N__73262;
    wire N__73257;
    wire N__73256;
    wire N__73253;
    wire N__73250;
    wire N__73247;
    wire N__73244;
    wire N__73241;
    wire N__73236;
    wire N__73233;
    wire N__73232;
    wire N__73231;
    wire N__73228;
    wire N__73225;
    wire N__73222;
    wire N__73221;
    wire N__73218;
    wire N__73215;
    wire N__73212;
    wire N__73211;
    wire N__73208;
    wire N__73205;
    wire N__73202;
    wire N__73199;
    wire N__73196;
    wire N__73185;
    wire N__73182;
    wire N__73179;
    wire N__73176;
    wire N__73173;
    wire N__73170;
    wire N__73169;
    wire N__73166;
    wire N__73163;
    wire N__73162;
    wire N__73159;
    wire N__73156;
    wire N__73153;
    wire N__73148;
    wire N__73143;
    wire N__73140;
    wire N__73137;
    wire N__73134;
    wire N__73133;
    wire N__73132;
    wire N__73131;
    wire N__73128;
    wire N__73123;
    wire N__73120;
    wire N__73115;
    wire N__73110;
    wire N__73107;
    wire N__73104;
    wire N__73101;
    wire N__73098;
    wire N__73097;
    wire N__73094;
    wire N__73091;
    wire N__73090;
    wire N__73087;
    wire N__73084;
    wire N__73081;
    wire N__73080;
    wire N__73079;
    wire N__73076;
    wire N__73073;
    wire N__73070;
    wire N__73067;
    wire N__73064;
    wire N__73055;
    wire N__73050;
    wire N__73047;
    wire N__73046;
    wire N__73045;
    wire N__73042;
    wire N__73041;
    wire N__73040;
    wire N__73039;
    wire N__73038;
    wire N__73037;
    wire N__73036;
    wire N__73033;
    wire N__73032;
    wire N__73031;
    wire N__73030;
    wire N__73029;
    wire N__73028;
    wire N__73027;
    wire N__73026;
    wire N__73025;
    wire N__73024;
    wire N__73023;
    wire N__73022;
    wire N__73021;
    wire N__73020;
    wire N__73019;
    wire N__73018;
    wire N__73017;
    wire N__73016;
    wire N__73015;
    wire N__73014;
    wire N__73013;
    wire N__73012;
    wire N__73011;
    wire N__73010;
    wire N__73009;
    wire N__73008;
    wire N__73007;
    wire N__73006;
    wire N__73003;
    wire N__73000;
    wire N__72995;
    wire N__72992;
    wire N__72987;
    wire N__72986;
    wire N__72985;
    wire N__72984;
    wire N__72983;
    wire N__72982;
    wire N__72979;
    wire N__72976;
    wire N__72975;
    wire N__72972;
    wire N__72969;
    wire N__72964;
    wire N__72961;
    wire N__72958;
    wire N__72955;
    wire N__72944;
    wire N__72937;
    wire N__72926;
    wire N__72925;
    wire N__72924;
    wire N__72913;
    wire N__72910;
    wire N__72907;
    wire N__72904;
    wire N__72903;
    wire N__72902;
    wire N__72897;
    wire N__72892;
    wire N__72889;
    wire N__72886;
    wire N__72881;
    wire N__72880;
    wire N__72879;
    wire N__72876;
    wire N__72871;
    wire N__72870;
    wire N__72869;
    wire N__72868;
    wire N__72867;
    wire N__72866;
    wire N__72863;
    wire N__72860;
    wire N__72851;
    wire N__72842;
    wire N__72837;
    wire N__72834;
    wire N__72831;
    wire N__72828;
    wire N__72825;
    wire N__72820;
    wire N__72817;
    wire N__72812;
    wire N__72807;
    wire N__72804;
    wire N__72803;
    wire N__72800;
    wire N__72799;
    wire N__72796;
    wire N__72793;
    wire N__72790;
    wire N__72785;
    wire N__72780;
    wire N__72771;
    wire N__72766;
    wire N__72763;
    wire N__72750;
    wire N__72745;
    wire N__72740;
    wire N__72735;
    wire N__72726;
    wire N__72719;
    wire N__72708;
    wire N__72705;
    wire N__72704;
    wire N__72701;
    wire N__72700;
    wire N__72697;
    wire N__72694;
    wire N__72691;
    wire N__72684;
    wire N__72681;
    wire N__72678;
    wire N__72675;
    wire N__72672;
    wire N__72669;
    wire N__72666;
    wire N__72663;
    wire N__72662;
    wire N__72661;
    wire N__72660;
    wire N__72655;
    wire N__72652;
    wire N__72651;
    wire N__72650;
    wire N__72647;
    wire N__72644;
    wire N__72641;
    wire N__72636;
    wire N__72631;
    wire N__72624;
    wire N__72623;
    wire N__72618;
    wire N__72615;
    wire N__72612;
    wire N__72609;
    wire N__72606;
    wire N__72603;
    wire N__72600;
    wire N__72597;
    wire N__72596;
    wire N__72593;
    wire N__72590;
    wire N__72589;
    wire N__72588;
    wire N__72585;
    wire N__72582;
    wire N__72579;
    wire N__72576;
    wire N__72575;
    wire N__72572;
    wire N__72569;
    wire N__72566;
    wire N__72563;
    wire N__72560;
    wire N__72557;
    wire N__72550;
    wire N__72543;
    wire N__72540;
    wire N__72537;
    wire N__72534;
    wire N__72531;
    wire N__72528;
    wire N__72525;
    wire N__72522;
    wire N__72521;
    wire N__72516;
    wire N__72515;
    wire N__72512;
    wire N__72509;
    wire N__72506;
    wire N__72503;
    wire N__72500;
    wire N__72495;
    wire N__72492;
    wire N__72489;
    wire N__72486;
    wire N__72483;
    wire N__72480;
    wire N__72477;
    wire N__72474;
    wire N__72471;
    wire N__72468;
    wire N__72465;
    wire N__72464;
    wire N__72461;
    wire N__72460;
    wire N__72457;
    wire N__72456;
    wire N__72455;
    wire N__72454;
    wire N__72451;
    wire N__72448;
    wire N__72445;
    wire N__72438;
    wire N__72429;
    wire N__72426;
    wire N__72425;
    wire N__72422;
    wire N__72419;
    wire N__72418;
    wire N__72417;
    wire N__72416;
    wire N__72415;
    wire N__72412;
    wire N__72409;
    wire N__72406;
    wire N__72401;
    wire N__72398;
    wire N__72393;
    wire N__72388;
    wire N__72381;
    wire N__72380;
    wire N__72379;
    wire N__72376;
    wire N__72373;
    wire N__72370;
    wire N__72367;
    wire N__72366;
    wire N__72363;
    wire N__72362;
    wire N__72359;
    wire N__72356;
    wire N__72353;
    wire N__72350;
    wire N__72347;
    wire N__72344;
    wire N__72333;
    wire N__72330;
    wire N__72329;
    wire N__72326;
    wire N__72323;
    wire N__72318;
    wire N__72315;
    wire N__72312;
    wire N__72309;
    wire N__72308;
    wire N__72305;
    wire N__72304;
    wire N__72303;
    wire N__72302;
    wire N__72299;
    wire N__72296;
    wire N__72293;
    wire N__72288;
    wire N__72279;
    wire N__72278;
    wire N__72275;
    wire N__72274;
    wire N__72273;
    wire N__72270;
    wire N__72267;
    wire N__72264;
    wire N__72261;
    wire N__72260;
    wire N__72253;
    wire N__72250;
    wire N__72247;
    wire N__72244;
    wire N__72237;
    wire N__72234;
    wire N__72231;
    wire N__72228;
    wire N__72225;
    wire N__72222;
    wire N__72221;
    wire N__72218;
    wire N__72215;
    wire N__72212;
    wire N__72207;
    wire N__72204;
    wire N__72203;
    wire N__72202;
    wire N__72201;
    wire N__72198;
    wire N__72197;
    wire N__72194;
    wire N__72189;
    wire N__72188;
    wire N__72185;
    wire N__72182;
    wire N__72177;
    wire N__72174;
    wire N__72171;
    wire N__72166;
    wire N__72159;
    wire N__72158;
    wire N__72155;
    wire N__72154;
    wire N__72153;
    wire N__72152;
    wire N__72149;
    wire N__72148;
    wire N__72145;
    wire N__72138;
    wire N__72135;
    wire N__72132;
    wire N__72129;
    wire N__72126;
    wire N__72117;
    wire N__72114;
    wire N__72111;
    wire N__72108;
    wire N__72105;
    wire N__72102;
    wire N__72099;
    wire N__72098;
    wire N__72095;
    wire N__72092;
    wire N__72087;
    wire N__72084;
    wire N__72081;
    wire N__72078;
    wire N__72077;
    wire N__72074;
    wire N__72073;
    wire N__72070;
    wire N__72069;
    wire N__72066;
    wire N__72063;
    wire N__72062;
    wire N__72059;
    wire N__72056;
    wire N__72053;
    wire N__72050;
    wire N__72047;
    wire N__72046;
    wire N__72043;
    wire N__72040;
    wire N__72033;
    wire N__72030;
    wire N__72027;
    wire N__72022;
    wire N__72015;
    wire N__72012;
    wire N__72009;
    wire N__72008;
    wire N__72005;
    wire N__72004;
    wire N__72003;
    wire N__72002;
    wire N__72001;
    wire N__71998;
    wire N__71995;
    wire N__71992;
    wire N__71989;
    wire N__71984;
    wire N__71983;
    wire N__71980;
    wire N__71977;
    wire N__71974;
    wire N__71971;
    wire N__71968;
    wire N__71965;
    wire N__71960;
    wire N__71955;
    wire N__71952;
    wire N__71943;
    wire N__71940;
    wire N__71937;
    wire N__71934;
    wire N__71931;
    wire N__71928;
    wire N__71925;
    wire N__71922;
    wire N__71919;
    wire N__71918;
    wire N__71915;
    wire N__71912;
    wire N__71909;
    wire N__71904;
    wire N__71901;
    wire N__71898;
    wire N__71895;
    wire N__71892;
    wire N__71891;
    wire N__71890;
    wire N__71889;
    wire N__71886;
    wire N__71883;
    wire N__71880;
    wire N__71877;
    wire N__71872;
    wire N__71871;
    wire N__71868;
    wire N__71863;
    wire N__71860;
    wire N__71853;
    wire N__71852;
    wire N__71849;
    wire N__71846;
    wire N__71841;
    wire N__71840;
    wire N__71837;
    wire N__71834;
    wire N__71829;
    wire N__71826;
    wire N__71823;
    wire N__71820;
    wire N__71817;
    wire N__71816;
    wire N__71811;
    wire N__71808;
    wire N__71805;
    wire N__71804;
    wire N__71801;
    wire N__71800;
    wire N__71797;
    wire N__71794;
    wire N__71791;
    wire N__71790;
    wire N__71787;
    wire N__71782;
    wire N__71779;
    wire N__71774;
    wire N__71769;
    wire N__71766;
    wire N__71763;
    wire N__71760;
    wire N__71757;
    wire N__71756;
    wire N__71753;
    wire N__71750;
    wire N__71745;
    wire N__71742;
    wire N__71739;
    wire N__71736;
    wire N__71733;
    wire N__71730;
    wire N__71727;
    wire N__71724;
    wire N__71721;
    wire N__71718;
    wire N__71717;
    wire N__71714;
    wire N__71711;
    wire N__71708;
    wire N__71703;
    wire N__71700;
    wire N__71697;
    wire N__71694;
    wire N__71691;
    wire N__71690;
    wire N__71689;
    wire N__71688;
    wire N__71685;
    wire N__71682;
    wire N__71677;
    wire N__71676;
    wire N__71673;
    wire N__71670;
    wire N__71667;
    wire N__71666;
    wire N__71663;
    wire N__71662;
    wire N__71655;
    wire N__71652;
    wire N__71651;
    wire N__71648;
    wire N__71645;
    wire N__71640;
    wire N__71637;
    wire N__71634;
    wire N__71631;
    wire N__71628;
    wire N__71625;
    wire N__71616;
    wire N__71613;
    wire N__71610;
    wire N__71609;
    wire N__71606;
    wire N__71603;
    wire N__71600;
    wire N__71595;
    wire N__71592;
    wire N__71589;
    wire N__71586;
    wire N__71583;
    wire N__71580;
    wire N__71577;
    wire N__71574;
    wire N__71571;
    wire N__71568;
    wire N__71565;
    wire N__71562;
    wire N__71559;
    wire N__71556;
    wire N__71553;
    wire N__71550;
    wire N__71547;
    wire N__71544;
    wire N__71541;
    wire N__71538;
    wire N__71537;
    wire N__71532;
    wire N__71529;
    wire N__71526;
    wire N__71523;
    wire N__71520;
    wire N__71517;
    wire N__71514;
    wire N__71511;
    wire N__71508;
    wire N__71505;
    wire N__71504;
    wire N__71503;
    wire N__71502;
    wire N__71501;
    wire N__71500;
    wire N__71499;
    wire N__71498;
    wire N__71497;
    wire N__71496;
    wire N__71495;
    wire N__71494;
    wire N__71493;
    wire N__71492;
    wire N__71491;
    wire N__71490;
    wire N__71489;
    wire N__71488;
    wire N__71485;
    wire N__71482;
    wire N__71479;
    wire N__71476;
    wire N__71475;
    wire N__71474;
    wire N__71473;
    wire N__71472;
    wire N__71469;
    wire N__71466;
    wire N__71463;
    wire N__71460;
    wire N__71457;
    wire N__71454;
    wire N__71451;
    wire N__71448;
    wire N__71447;
    wire N__71446;
    wire N__71445;
    wire N__71444;
    wire N__71441;
    wire N__71438;
    wire N__71435;
    wire N__71432;
    wire N__71429;
    wire N__71426;
    wire N__71417;
    wire N__71414;
    wire N__71411;
    wire N__71410;
    wire N__71407;
    wire N__71404;
    wire N__71401;
    wire N__71394;
    wire N__71385;
    wire N__71382;
    wire N__71379;
    wire N__71376;
    wire N__71373;
    wire N__71368;
    wire N__71363;
    wire N__71356;
    wire N__71351;
    wire N__71348;
    wire N__71337;
    wire N__71332;
    wire N__71323;
    wire N__71322;
    wire N__71317;
    wire N__71316;
    wire N__71313;
    wire N__71310;
    wire N__71305;
    wire N__71302;
    wire N__71299;
    wire N__71296;
    wire N__71293;
    wire N__71290;
    wire N__71287;
    wire N__71282;
    wire N__71271;
    wire N__71270;
    wire N__71267;
    wire N__71264;
    wire N__71263;
    wire N__71262;
    wire N__71259;
    wire N__71256;
    wire N__71251;
    wire N__71248;
    wire N__71245;
    wire N__71242;
    wire N__71239;
    wire N__71234;
    wire N__71233;
    wire N__71230;
    wire N__71227;
    wire N__71224;
    wire N__71221;
    wire N__71218;
    wire N__71211;
    wire N__71208;
    wire N__71205;
    wire N__71202;
    wire N__71199;
    wire N__71196;
    wire N__71193;
    wire N__71190;
    wire N__71187;
    wire N__71184;
    wire N__71181;
    wire N__71178;
    wire N__71175;
    wire N__71172;
    wire N__71169;
    wire N__71166;
    wire N__71163;
    wire N__71160;
    wire N__71159;
    wire N__71156;
    wire N__71155;
    wire N__71154;
    wire N__71151;
    wire N__71148;
    wire N__71147;
    wire N__71146;
    wire N__71143;
    wire N__71140;
    wire N__71137;
    wire N__71134;
    wire N__71131;
    wire N__71128;
    wire N__71125;
    wire N__71124;
    wire N__71121;
    wire N__71118;
    wire N__71115;
    wire N__71114;
    wire N__71113;
    wire N__71112;
    wire N__71109;
    wire N__71106;
    wire N__71103;
    wire N__71100;
    wire N__71097;
    wire N__71092;
    wire N__71085;
    wire N__71070;
    wire N__71069;
    wire N__71066;
    wire N__71063;
    wire N__71062;
    wire N__71057;
    wire N__71054;
    wire N__71049;
    wire N__71048;
    wire N__71045;
    wire N__71042;
    wire N__71041;
    wire N__71036;
    wire N__71033;
    wire N__71030;
    wire N__71027;
    wire N__71022;
    wire N__71019;
    wire N__71016;
    wire N__71015;
    wire N__71012;
    wire N__71009;
    wire N__71004;
    wire N__71003;
    wire N__71000;
    wire N__70997;
    wire N__70992;
    wire N__70991;
    wire N__70988;
    wire N__70985;
    wire N__70980;
    wire N__70979;
    wire N__70976;
    wire N__70973;
    wire N__70968;
    wire N__70965;
    wire N__70962;
    wire N__70961;
    wire N__70958;
    wire N__70955;
    wire N__70952;
    wire N__70949;
    wire N__70948;
    wire N__70943;
    wire N__70940;
    wire N__70935;
    wire N__70934;
    wire N__70933;
    wire N__70930;
    wire N__70925;
    wire N__70920;
    wire N__70917;
    wire N__70914;
    wire N__70911;
    wire N__70910;
    wire N__70907;
    wire N__70904;
    wire N__70903;
    wire N__70898;
    wire N__70895;
    wire N__70892;
    wire N__70889;
    wire N__70884;
    wire N__70883;
    wire N__70880;
    wire N__70877;
    wire N__70872;
    wire N__70871;
    wire N__70868;
    wire N__70865;
    wire N__70860;
    wire N__70857;
    wire N__70856;
    wire N__70853;
    wire N__70850;
    wire N__70849;
    wire N__70844;
    wire N__70841;
    wire N__70836;
    wire N__70835;
    wire N__70834;
    wire N__70833;
    wire N__70830;
    wire N__70827;
    wire N__70824;
    wire N__70821;
    wire N__70820;
    wire N__70819;
    wire N__70818;
    wire N__70817;
    wire N__70816;
    wire N__70815;
    wire N__70814;
    wire N__70813;
    wire N__70808;
    wire N__70803;
    wire N__70800;
    wire N__70797;
    wire N__70794;
    wire N__70791;
    wire N__70788;
    wire N__70785;
    wire N__70782;
    wire N__70779;
    wire N__70778;
    wire N__70777;
    wire N__70772;
    wire N__70763;
    wire N__70754;
    wire N__70751;
    wire N__70748;
    wire N__70741;
    wire N__70736;
    wire N__70731;
    wire N__70728;
    wire N__70727;
    wire N__70724;
    wire N__70721;
    wire N__70716;
    wire N__70715;
    wire N__70712;
    wire N__70709;
    wire N__70704;
    wire N__70701;
    wire N__70698;
    wire N__70697;
    wire N__70696;
    wire N__70693;
    wire N__70690;
    wire N__70687;
    wire N__70684;
    wire N__70677;
    wire N__70674;
    wire N__70671;
    wire N__70668;
    wire N__70667;
    wire N__70666;
    wire N__70663;
    wire N__70660;
    wire N__70657;
    wire N__70654;
    wire N__70647;
    wire N__70644;
    wire N__70641;
    wire N__70638;
    wire N__70635;
    wire N__70632;
    wire N__70629;
    wire N__70628;
    wire N__70627;
    wire N__70624;
    wire N__70621;
    wire N__70618;
    wire N__70615;
    wire N__70610;
    wire N__70607;
    wire N__70602;
    wire N__70601;
    wire N__70598;
    wire N__70595;
    wire N__70594;
    wire N__70589;
    wire N__70586;
    wire N__70581;
    wire N__70578;
    wire N__70575;
    wire N__70572;
    wire N__70569;
    wire N__70566;
    wire N__70563;
    wire N__70560;
    wire N__70559;
    wire N__70556;
    wire N__70553;
    wire N__70552;
    wire N__70547;
    wire N__70544;
    wire N__70539;
    wire N__70536;
    wire N__70535;
    wire N__70532;
    wire N__70529;
    wire N__70524;
    wire N__70523;
    wire N__70520;
    wire N__70517;
    wire N__70512;
    wire N__70509;
    wire N__70508;
    wire N__70505;
    wire N__70502;
    wire N__70497;
    wire N__70496;
    wire N__70493;
    wire N__70490;
    wire N__70485;
    wire N__70484;
    wire N__70481;
    wire N__70478;
    wire N__70477;
    wire N__70472;
    wire N__70469;
    wire N__70466;
    wire N__70463;
    wire N__70458;
    wire N__70455;
    wire N__70454;
    wire N__70451;
    wire N__70448;
    wire N__70447;
    wire N__70442;
    wire N__70439;
    wire N__70436;
    wire N__70433;
    wire N__70428;
    wire N__70425;
    wire N__70424;
    wire N__70421;
    wire N__70418;
    wire N__70417;
    wire N__70412;
    wire N__70409;
    wire N__70404;
    wire N__70401;
    wire N__70400;
    wire N__70397;
    wire N__70394;
    wire N__70393;
    wire N__70388;
    wire N__70385;
    wire N__70382;
    wire N__70379;
    wire N__70374;
    wire N__70373;
    wire N__70370;
    wire N__70367;
    wire N__70364;
    wire N__70363;
    wire N__70358;
    wire N__70355;
    wire N__70350;
    wire N__70347;
    wire N__70346;
    wire N__70343;
    wire N__70340;
    wire N__70339;
    wire N__70334;
    wire N__70331;
    wire N__70326;
    wire N__70323;
    wire N__70322;
    wire N__70319;
    wire N__70316;
    wire N__70315;
    wire N__70310;
    wire N__70307;
    wire N__70302;
    wire N__70299;
    wire N__70298;
    wire N__70295;
    wire N__70292;
    wire N__70291;
    wire N__70286;
    wire N__70283;
    wire N__70278;
    wire N__70277;
    wire N__70274;
    wire N__70273;
    wire N__70270;
    wire N__70267;
    wire N__70264;
    wire N__70259;
    wire N__70256;
    wire N__70251;
    wire N__70248;
    wire N__70247;
    wire N__70246;
    wire N__70243;
    wire N__70240;
    wire N__70237;
    wire N__70232;
    wire N__70229;
    wire N__70224;
    wire N__70223;
    wire N__70220;
    wire N__70217;
    wire N__70214;
    wire N__70213;
    wire N__70208;
    wire N__70205;
    wire N__70200;
    wire N__70197;
    wire N__70194;
    wire N__70191;
    wire N__70188;
    wire N__70185;
    wire N__70182;
    wire N__70181;
    wire N__70178;
    wire N__70175;
    wire N__70172;
    wire N__70169;
    wire N__70168;
    wire N__70163;
    wire N__70160;
    wire N__70155;
    wire N__70152;
    wire N__70151;
    wire N__70148;
    wire N__70145;
    wire N__70144;
    wire N__70139;
    wire N__70136;
    wire N__70133;
    wire N__70130;
    wire N__70125;
    wire N__70122;
    wire N__70121;
    wire N__70118;
    wire N__70115;
    wire N__70114;
    wire N__70109;
    wire N__70106;
    wire N__70101;
    wire N__70098;
    wire N__70097;
    wire N__70094;
    wire N__70091;
    wire N__70088;
    wire N__70087;
    wire N__70082;
    wire N__70079;
    wire N__70074;
    wire N__70071;
    wire N__70070;
    wire N__70069;
    wire N__70066;
    wire N__70063;
    wire N__70060;
    wire N__70053;
    wire N__70050;
    wire N__70049;
    wire N__70046;
    wire N__70043;
    wire N__70040;
    wire N__70039;
    wire N__70034;
    wire N__70031;
    wire N__70026;
    wire N__70023;
    wire N__70022;
    wire N__70021;
    wire N__70018;
    wire N__70015;
    wire N__70012;
    wire N__70007;
    wire N__70004;
    wire N__69999;
    wire N__69996;
    wire N__69993;
    wire N__69992;
    wire N__69991;
    wire N__69988;
    wire N__69985;
    wire N__69982;
    wire N__69975;
    wire N__69972;
    wire N__69971;
    wire N__69970;
    wire N__69969;
    wire N__69968;
    wire N__69967;
    wire N__69964;
    wire N__69961;
    wire N__69958;
    wire N__69955;
    wire N__69952;
    wire N__69949;
    wire N__69944;
    wire N__69935;
    wire N__69930;
    wire N__69929;
    wire N__69926;
    wire N__69923;
    wire N__69920;
    wire N__69919;
    wire N__69914;
    wire N__69911;
    wire N__69906;
    wire N__69903;
    wire N__69902;
    wire N__69899;
    wire N__69896;
    wire N__69895;
    wire N__69890;
    wire N__69887;
    wire N__69882;
    wire N__69879;
    wire N__69876;
    wire N__69875;
    wire N__69872;
    wire N__69869;
    wire N__69866;
    wire N__69863;
    wire N__69862;
    wire N__69859;
    wire N__69856;
    wire N__69853;
    wire N__69846;
    wire N__69843;
    wire N__69840;
    wire N__69837;
    wire N__69836;
    wire N__69835;
    wire N__69832;
    wire N__69829;
    wire N__69826;
    wire N__69823;
    wire N__69818;
    wire N__69813;
    wire N__69810;
    wire N__69809;
    wire N__69806;
    wire N__69805;
    wire N__69802;
    wire N__69799;
    wire N__69796;
    wire N__69793;
    wire N__69790;
    wire N__69785;
    wire N__69780;
    wire N__69777;
    wire N__69774;
    wire N__69773;
    wire N__69772;
    wire N__69769;
    wire N__69766;
    wire N__69763;
    wire N__69760;
    wire N__69753;
    wire N__69750;
    wire N__69747;
    wire N__69744;
    wire N__69741;
    wire N__69738;
    wire N__69735;
    wire N__69732;
    wire N__69731;
    wire N__69728;
    wire N__69725;
    wire N__69724;
    wire N__69721;
    wire N__69718;
    wire N__69715;
    wire N__69708;
    wire N__69705;
    wire N__69704;
    wire N__69701;
    wire N__69698;
    wire N__69697;
    wire N__69692;
    wire N__69689;
    wire N__69684;
    wire N__69681;
    wire N__69678;
    wire N__69677;
    wire N__69674;
    wire N__69671;
    wire N__69670;
    wire N__69667;
    wire N__69664;
    wire N__69661;
    wire N__69654;
    wire N__69651;
    wire N__69648;
    wire N__69647;
    wire N__69646;
    wire N__69643;
    wire N__69640;
    wire N__69637;
    wire N__69630;
    wire N__69627;
    wire N__69624;
    wire N__69621;
    wire N__69620;
    wire N__69619;
    wire N__69616;
    wire N__69613;
    wire N__69610;
    wire N__69607;
    wire N__69602;
    wire N__69597;
    wire N__69594;
    wire N__69593;
    wire N__69592;
    wire N__69589;
    wire N__69586;
    wire N__69583;
    wire N__69580;
    wire N__69575;
    wire N__69570;
    wire N__69569;
    wire N__69568;
    wire N__69567;
    wire N__69566;
    wire N__69565;
    wire N__69562;
    wire N__69559;
    wire N__69556;
    wire N__69553;
    wire N__69550;
    wire N__69547;
    wire N__69542;
    wire N__69533;
    wire N__69528;
    wire N__69525;
    wire N__69524;
    wire N__69523;
    wire N__69522;
    wire N__69521;
    wire N__69520;
    wire N__69519;
    wire N__69518;
    wire N__69517;
    wire N__69516;
    wire N__69515;
    wire N__69512;
    wire N__69509;
    wire N__69506;
    wire N__69503;
    wire N__69500;
    wire N__69497;
    wire N__69494;
    wire N__69491;
    wire N__69488;
    wire N__69485;
    wire N__69482;
    wire N__69477;
    wire N__69476;
    wire N__69473;
    wire N__69464;
    wire N__69455;
    wire N__69452;
    wire N__69449;
    wire N__69438;
    wire N__69435;
    wire N__69432;
    wire N__69429;
    wire N__69426;
    wire N__69425;
    wire N__69424;
    wire N__69421;
    wire N__69418;
    wire N__69415;
    wire N__69410;
    wire N__69407;
    wire N__69402;
    wire N__69399;
    wire N__69398;
    wire N__69395;
    wire N__69392;
    wire N__69391;
    wire N__69386;
    wire N__69383;
    wire N__69378;
    wire N__69375;
    wire N__69374;
    wire N__69371;
    wire N__69368;
    wire N__69367;
    wire N__69362;
    wire N__69359;
    wire N__69354;
    wire N__69351;
    wire N__69350;
    wire N__69349;
    wire N__69346;
    wire N__69343;
    wire N__69340;
    wire N__69333;
    wire N__69330;
    wire N__69327;
    wire N__69324;
    wire N__69321;
    wire N__69318;
    wire N__69315;
    wire N__69312;
    wire N__69311;
    wire N__69306;
    wire N__69303;
    wire N__69300;
    wire N__69299;
    wire N__69296;
    wire N__69293;
    wire N__69292;
    wire N__69289;
    wire N__69284;
    wire N__69279;
    wire N__69276;
    wire N__69275;
    wire N__69272;
    wire N__69269;
    wire N__69264;
    wire N__69261;
    wire N__69258;
    wire N__69255;
    wire N__69252;
    wire N__69249;
    wire N__69248;
    wire N__69245;
    wire N__69244;
    wire N__69241;
    wire N__69238;
    wire N__69235;
    wire N__69232;
    wire N__69229;
    wire N__69226;
    wire N__69221;
    wire N__69218;
    wire N__69213;
    wire N__69212;
    wire N__69209;
    wire N__69206;
    wire N__69203;
    wire N__69200;
    wire N__69195;
    wire N__69192;
    wire N__69189;
    wire N__69186;
    wire N__69183;
    wire N__69180;
    wire N__69179;
    wire N__69176;
    wire N__69173;
    wire N__69170;
    wire N__69167;
    wire N__69162;
    wire N__69159;
    wire N__69158;
    wire N__69155;
    wire N__69152;
    wire N__69147;
    wire N__69144;
    wire N__69141;
    wire N__69138;
    wire N__69135;
    wire N__69134;
    wire N__69131;
    wire N__69130;
    wire N__69129;
    wire N__69126;
    wire N__69123;
    wire N__69118;
    wire N__69111;
    wire N__69110;
    wire N__69109;
    wire N__69106;
    wire N__69101;
    wire N__69096;
    wire N__69095;
    wire N__69092;
    wire N__69087;
    wire N__69084;
    wire N__69083;
    wire N__69080;
    wire N__69079;
    wire N__69076;
    wire N__69075;
    wire N__69072;
    wire N__69069;
    wire N__69066;
    wire N__69063;
    wire N__69058;
    wire N__69055;
    wire N__69050;
    wire N__69045;
    wire N__69044;
    wire N__69041;
    wire N__69038;
    wire N__69035;
    wire N__69034;
    wire N__69029;
    wire N__69026;
    wire N__69021;
    wire N__69018;
    wire N__69017;
    wire N__69014;
    wire N__69013;
    wire N__69012;
    wire N__69009;
    wire N__69006;
    wire N__69001;
    wire N__68998;
    wire N__68991;
    wire N__68988;
    wire N__68985;
    wire N__68984;
    wire N__68981;
    wire N__68978;
    wire N__68973;
    wire N__68972;
    wire N__68969;
    wire N__68966;
    wire N__68963;
    wire N__68960;
    wire N__68955;
    wire N__68954;
    wire N__68953;
    wire N__68948;
    wire N__68945;
    wire N__68940;
    wire N__68939;
    wire N__68936;
    wire N__68933;
    wire N__68930;
    wire N__68927;
    wire N__68924;
    wire N__68921;
    wire N__68918;
    wire N__68913;
    wire N__68912;
    wire N__68911;
    wire N__68910;
    wire N__68905;
    wire N__68902;
    wire N__68899;
    wire N__68896;
    wire N__68895;
    wire N__68892;
    wire N__68887;
    wire N__68884;
    wire N__68881;
    wire N__68878;
    wire N__68871;
    wire N__68868;
    wire N__68865;
    wire N__68862;
    wire N__68859;
    wire N__68856;
    wire N__68853;
    wire N__68850;
    wire N__68847;
    wire N__68844;
    wire N__68841;
    wire N__68838;
    wire N__68835;
    wire N__68832;
    wire N__68829;
    wire N__68826;
    wire N__68825;
    wire N__68822;
    wire N__68821;
    wire N__68818;
    wire N__68813;
    wire N__68808;
    wire N__68807;
    wire N__68804;
    wire N__68801;
    wire N__68798;
    wire N__68793;
    wire N__68790;
    wire N__68789;
    wire N__68786;
    wire N__68785;
    wire N__68782;
    wire N__68779;
    wire N__68776;
    wire N__68773;
    wire N__68766;
    wire N__68763;
    wire N__68760;
    wire N__68757;
    wire N__68754;
    wire N__68751;
    wire N__68748;
    wire N__68745;
    wire N__68742;
    wire N__68739;
    wire N__68738;
    wire N__68735;
    wire N__68732;
    wire N__68731;
    wire N__68728;
    wire N__68723;
    wire N__68718;
    wire N__68715;
    wire N__68714;
    wire N__68711;
    wire N__68710;
    wire N__68707;
    wire N__68706;
    wire N__68703;
    wire N__68700;
    wire N__68695;
    wire N__68688;
    wire N__68687;
    wire N__68684;
    wire N__68681;
    wire N__68678;
    wire N__68675;
    wire N__68672;
    wire N__68667;
    wire N__68664;
    wire N__68663;
    wire N__68662;
    wire N__68659;
    wire N__68656;
    wire N__68655;
    wire N__68652;
    wire N__68647;
    wire N__68644;
    wire N__68641;
    wire N__68638;
    wire N__68631;
    wire N__68630;
    wire N__68625;
    wire N__68622;
    wire N__68619;
    wire N__68618;
    wire N__68615;
    wire N__68612;
    wire N__68609;
    wire N__68604;
    wire N__68601;
    wire N__68600;
    wire N__68595;
    wire N__68594;
    wire N__68591;
    wire N__68590;
    wire N__68589;
    wire N__68588;
    wire N__68585;
    wire N__68582;
    wire N__68581;
    wire N__68580;
    wire N__68575;
    wire N__68572;
    wire N__68567;
    wire N__68564;
    wire N__68563;
    wire N__68560;
    wire N__68557;
    wire N__68554;
    wire N__68551;
    wire N__68548;
    wire N__68545;
    wire N__68540;
    wire N__68535;
    wire N__68532;
    wire N__68523;
    wire N__68520;
    wire N__68519;
    wire N__68516;
    wire N__68515;
    wire N__68514;
    wire N__68511;
    wire N__68508;
    wire N__68505;
    wire N__68502;
    wire N__68499;
    wire N__68496;
    wire N__68491;
    wire N__68484;
    wire N__68481;
    wire N__68478;
    wire N__68475;
    wire N__68474;
    wire N__68473;
    wire N__68470;
    wire N__68467;
    wire N__68464;
    wire N__68461;
    wire N__68458;
    wire N__68455;
    wire N__68448;
    wire N__68445;
    wire N__68442;
    wire N__68439;
    wire N__68436;
    wire N__68433;
    wire N__68430;
    wire N__68427;
    wire N__68424;
    wire N__68421;
    wire N__68420;
    wire N__68415;
    wire N__68412;
    wire N__68409;
    wire N__68406;
    wire N__68403;
    wire N__68400;
    wire N__68399;
    wire N__68396;
    wire N__68393;
    wire N__68388;
    wire N__68387;
    wire N__68384;
    wire N__68381;
    wire N__68376;
    wire N__68373;
    wire N__68370;
    wire N__68367;
    wire N__68366;
    wire N__68363;
    wire N__68360;
    wire N__68355;
    wire N__68352;
    wire N__68349;
    wire N__68346;
    wire N__68343;
    wire N__68340;
    wire N__68337;
    wire N__68334;
    wire N__68331;
    wire N__68328;
    wire N__68325;
    wire N__68322;
    wire N__68319;
    wire N__68316;
    wire N__68313;
    wire N__68310;
    wire N__68307;
    wire N__68306;
    wire N__68305;
    wire N__68304;
    wire N__68303;
    wire N__68298;
    wire N__68297;
    wire N__68296;
    wire N__68293;
    wire N__68290;
    wire N__68287;
    wire N__68284;
    wire N__68281;
    wire N__68278;
    wire N__68273;
    wire N__68272;
    wire N__68269;
    wire N__68266;
    wire N__68265;
    wire N__68262;
    wire N__68259;
    wire N__68256;
    wire N__68253;
    wire N__68248;
    wire N__68245;
    wire N__68242;
    wire N__68235;
    wire N__68232;
    wire N__68227;
    wire N__68224;
    wire N__68217;
    wire N__68214;
    wire N__68213;
    wire N__68210;
    wire N__68207;
    wire N__68204;
    wire N__68201;
    wire N__68198;
    wire N__68193;
    wire N__68190;
    wire N__68187;
    wire N__68184;
    wire N__68183;
    wire N__68180;
    wire N__68177;
    wire N__68174;
    wire N__68171;
    wire N__68170;
    wire N__68169;
    wire N__68168;
    wire N__68165;
    wire N__68162;
    wire N__68159;
    wire N__68156;
    wire N__68153;
    wire N__68150;
    wire N__68145;
    wire N__68142;
    wire N__68133;
    wire N__68130;
    wire N__68127;
    wire N__68126;
    wire N__68121;
    wire N__68118;
    wire N__68115;
    wire N__68112;
    wire N__68111;
    wire N__68108;
    wire N__68105;
    wire N__68102;
    wire N__68097;
    wire N__68094;
    wire N__68093;
    wire N__68092;
    wire N__68089;
    wire N__68086;
    wire N__68083;
    wire N__68080;
    wire N__68079;
    wire N__68074;
    wire N__68073;
    wire N__68072;
    wire N__68069;
    wire N__68066;
    wire N__68063;
    wire N__68058;
    wire N__68049;
    wire N__68048;
    wire N__68045;
    wire N__68042;
    wire N__68037;
    wire N__68034;
    wire N__68031;
    wire N__68030;
    wire N__68029;
    wire N__68028;
    wire N__68025;
    wire N__68022;
    wire N__68019;
    wire N__68018;
    wire N__68015;
    wire N__68010;
    wire N__68007;
    wire N__68004;
    wire N__67995;
    wire N__67994;
    wire N__67991;
    wire N__67988;
    wire N__67985;
    wire N__67980;
    wire N__67977;
    wire N__67974;
    wire N__67971;
    wire N__67970;
    wire N__67965;
    wire N__67962;
    wire N__67959;
    wire N__67956;
    wire N__67953;
    wire N__67950;
    wire N__67947;
    wire N__67944;
    wire N__67941;
    wire N__67940;
    wire N__67939;
    wire N__67938;
    wire N__67937;
    wire N__67936;
    wire N__67933;
    wire N__67930;
    wire N__67925;
    wire N__67922;
    wire N__67919;
    wire N__67914;
    wire N__67909;
    wire N__67906;
    wire N__67903;
    wire N__67900;
    wire N__67893;
    wire N__67890;
    wire N__67889;
    wire N__67886;
    wire N__67883;
    wire N__67880;
    wire N__67875;
    wire N__67872;
    wire N__67871;
    wire N__67870;
    wire N__67867;
    wire N__67866;
    wire N__67863;
    wire N__67860;
    wire N__67857;
    wire N__67852;
    wire N__67849;
    wire N__67846;
    wire N__67839;
    wire N__67838;
    wire N__67835;
    wire N__67830;
    wire N__67827;
    wire N__67824;
    wire N__67821;
    wire N__67818;
    wire N__67815;
    wire N__67814;
    wire N__67811;
    wire N__67808;
    wire N__67805;
    wire N__67802;
    wire N__67799;
    wire N__67798;
    wire N__67793;
    wire N__67790;
    wire N__67789;
    wire N__67788;
    wire N__67785;
    wire N__67782;
    wire N__67777;
    wire N__67770;
    wire N__67767;
    wire N__67764;
    wire N__67763;
    wire N__67760;
    wire N__67757;
    wire N__67754;
    wire N__67749;
    wire N__67746;
    wire N__67743;
    wire N__67740;
    wire N__67737;
    wire N__67734;
    wire N__67731;
    wire N__67728;
    wire N__67725;
    wire N__67722;
    wire N__67719;
    wire N__67716;
    wire N__67715;
    wire N__67712;
    wire N__67709;
    wire N__67706;
    wire N__67701;
    wire N__67698;
    wire N__67695;
    wire N__67692;
    wire N__67689;
    wire N__67686;
    wire N__67683;
    wire N__67680;
    wire N__67677;
    wire N__67674;
    wire N__67673;
    wire N__67670;
    wire N__67667;
    wire N__67662;
    wire N__67659;
    wire N__67656;
    wire N__67653;
    wire N__67652;
    wire N__67651;
    wire N__67650;
    wire N__67649;
    wire N__67648;
    wire N__67647;
    wire N__67646;
    wire N__67645;
    wire N__67644;
    wire N__67643;
    wire N__67642;
    wire N__67639;
    wire N__67636;
    wire N__67635;
    wire N__67634;
    wire N__67633;
    wire N__67630;
    wire N__67627;
    wire N__67624;
    wire N__67621;
    wire N__67618;
    wire N__67615;
    wire N__67612;
    wire N__67609;
    wire N__67606;
    wire N__67603;
    wire N__67598;
    wire N__67595;
    wire N__67592;
    wire N__67589;
    wire N__67588;
    wire N__67583;
    wire N__67574;
    wire N__67565;
    wire N__67562;
    wire N__67553;
    wire N__67542;
    wire N__67539;
    wire N__67536;
    wire N__67535;
    wire N__67532;
    wire N__67529;
    wire N__67524;
    wire N__67521;
    wire N__67518;
    wire N__67515;
    wire N__67512;
    wire N__67509;
    wire N__67506;
    wire N__67503;
    wire N__67500;
    wire N__67497;
    wire N__67494;
    wire N__67491;
    wire N__67488;
    wire N__67485;
    wire N__67482;
    wire N__67479;
    wire N__67478;
    wire N__67473;
    wire N__67470;
    wire N__67467;
    wire N__67464;
    wire N__67463;
    wire N__67460;
    wire N__67457;
    wire N__67454;
    wire N__67449;
    wire N__67446;
    wire N__67443;
    wire N__67440;
    wire N__67437;
    wire N__67434;
    wire N__67431;
    wire N__67428;
    wire N__67427;
    wire N__67426;
    wire N__67425;
    wire N__67424;
    wire N__67423;
    wire N__67420;
    wire N__67417;
    wire N__67414;
    wire N__67411;
    wire N__67408;
    wire N__67405;
    wire N__67400;
    wire N__67391;
    wire N__67386;
    wire N__67383;
    wire N__67380;
    wire N__67377;
    wire N__67374;
    wire N__67371;
    wire N__67368;
    wire N__67365;
    wire N__67362;
    wire N__67359;
    wire N__67356;
    wire N__67353;
    wire N__67350;
    wire N__67347;
    wire N__67344;
    wire N__67341;
    wire N__67338;
    wire N__67335;
    wire N__67332;
    wire N__67329;
    wire N__67326;
    wire N__67323;
    wire N__67320;
    wire N__67317;
    wire N__67314;
    wire N__67311;
    wire N__67310;
    wire N__67309;
    wire N__67306;
    wire N__67303;
    wire N__67300;
    wire N__67295;
    wire N__67292;
    wire N__67287;
    wire N__67284;
    wire N__67283;
    wire N__67282;
    wire N__67279;
    wire N__67276;
    wire N__67273;
    wire N__67268;
    wire N__67265;
    wire N__67260;
    wire N__67257;
    wire N__67256;
    wire N__67253;
    wire N__67250;
    wire N__67245;
    wire N__67244;
    wire N__67241;
    wire N__67238;
    wire N__67233;
    wire N__67230;
    wire N__67229;
    wire N__67226;
    wire N__67223;
    wire N__67222;
    wire N__67217;
    wire N__67214;
    wire N__67209;
    wire N__67206;
    wire N__67205;
    wire N__67202;
    wire N__67199;
    wire N__67196;
    wire N__67195;
    wire N__67192;
    wire N__67189;
    wire N__67186;
    wire N__67179;
    wire N__67178;
    wire N__67177;
    wire N__67176;
    wire N__67175;
    wire N__67174;
    wire N__67173;
    wire N__67172;
    wire N__67171;
    wire N__67170;
    wire N__67169;
    wire N__67168;
    wire N__67167;
    wire N__67164;
    wire N__67161;
    wire N__67158;
    wire N__67155;
    wire N__67152;
    wire N__67149;
    wire N__67146;
    wire N__67143;
    wire N__67140;
    wire N__67137;
    wire N__67134;
    wire N__67131;
    wire N__67128;
    wire N__67123;
    wire N__67120;
    wire N__67115;
    wire N__67106;
    wire N__67097;
    wire N__67094;
    wire N__67083;
    wire N__67080;
    wire N__67077;
    wire N__67074;
    wire N__67071;
    wire N__67070;
    wire N__67067;
    wire N__67064;
    wire N__67063;
    wire N__67058;
    wire N__67055;
    wire N__67050;
    wire N__67049;
    wire N__67048;
    wire N__67047;
    wire N__67046;
    wire N__67045;
    wire N__67042;
    wire N__67039;
    wire N__67036;
    wire N__67033;
    wire N__67030;
    wire N__67027;
    wire N__67022;
    wire N__67013;
    wire N__67008;
    wire N__67005;
    wire N__67004;
    wire N__67001;
    wire N__66998;
    wire N__66997;
    wire N__66992;
    wire N__66989;
    wire N__66986;
    wire N__66983;
    wire N__66978;
    wire N__66975;
    wire N__66974;
    wire N__66971;
    wire N__66968;
    wire N__66967;
    wire N__66962;
    wire N__66959;
    wire N__66954;
    wire N__66951;
    wire N__66950;
    wire N__66947;
    wire N__66944;
    wire N__66943;
    wire N__66938;
    wire N__66935;
    wire N__66930;
    wire N__66927;
    wire N__66924;
    wire N__66923;
    wire N__66920;
    wire N__66917;
    wire N__66916;
    wire N__66911;
    wire N__66908;
    wire N__66905;
    wire N__66902;
    wire N__66897;
    wire N__66894;
    wire N__66893;
    wire N__66892;
    wire N__66889;
    wire N__66886;
    wire N__66883;
    wire N__66878;
    wire N__66875;
    wire N__66872;
    wire N__66869;
    wire N__66864;
    wire N__66861;
    wire N__66860;
    wire N__66857;
    wire N__66854;
    wire N__66849;
    wire N__66848;
    wire N__66845;
    wire N__66842;
    wire N__66837;
    wire N__66834;
    wire N__66833;
    wire N__66830;
    wire N__66827;
    wire N__66822;
    wire N__66821;
    wire N__66818;
    wire N__66815;
    wire N__66810;
    wire N__66807;
    wire N__66804;
    wire N__66801;
    wire N__66800;
    wire N__66799;
    wire N__66796;
    wire N__66791;
    wire N__66788;
    wire N__66785;
    wire N__66780;
    wire N__66777;
    wire N__66774;
    wire N__66773;
    wire N__66772;
    wire N__66769;
    wire N__66766;
    wire N__66763;
    wire N__66760;
    wire N__66753;
    wire N__66750;
    wire N__66749;
    wire N__66746;
    wire N__66743;
    wire N__66738;
    wire N__66737;
    wire N__66734;
    wire N__66731;
    wire N__66726;
    wire N__66723;
    wire N__66722;
    wire N__66719;
    wire N__66716;
    wire N__66711;
    wire N__66710;
    wire N__66707;
    wire N__66704;
    wire N__66699;
    wire N__66696;
    wire N__66695;
    wire N__66692;
    wire N__66689;
    wire N__66688;
    wire N__66683;
    wire N__66680;
    wire N__66675;
    wire N__66672;
    wire N__66671;
    wire N__66668;
    wire N__66665;
    wire N__66664;
    wire N__66659;
    wire N__66656;
    wire N__66651;
    wire N__66648;
    wire N__66647;
    wire N__66644;
    wire N__66641;
    wire N__66640;
    wire N__66635;
    wire N__66632;
    wire N__66627;
    wire N__66624;
    wire N__66623;
    wire N__66622;
    wire N__66619;
    wire N__66616;
    wire N__66613;
    wire N__66610;
    wire N__66603;
    wire N__66600;
    wire N__66597;
    wire N__66594;
    wire N__66593;
    wire N__66590;
    wire N__66587;
    wire N__66586;
    wire N__66581;
    wire N__66578;
    wire N__66573;
    wire N__66570;
    wire N__66569;
    wire N__66568;
    wire N__66565;
    wire N__66562;
    wire N__66559;
    wire N__66552;
    wire N__66549;
    wire N__66548;
    wire N__66547;
    wire N__66544;
    wire N__66541;
    wire N__66538;
    wire N__66535;
    wire N__66528;
    wire N__66525;
    wire N__66524;
    wire N__66521;
    wire N__66520;
    wire N__66517;
    wire N__66514;
    wire N__66511;
    wire N__66506;
    wire N__66503;
    wire N__66498;
    wire N__66495;
    wire N__66492;
    wire N__66491;
    wire N__66490;
    wire N__66487;
    wire N__66484;
    wire N__66481;
    wire N__66478;
    wire N__66471;
    wire N__66468;
    wire N__66467;
    wire N__66466;
    wire N__66463;
    wire N__66460;
    wire N__66457;
    wire N__66450;
    wire N__66447;
    wire N__66446;
    wire N__66445;
    wire N__66442;
    wire N__66439;
    wire N__66436;
    wire N__66429;
    wire N__66426;
    wire N__66425;
    wire N__66424;
    wire N__66421;
    wire N__66418;
    wire N__66415;
    wire N__66408;
    wire N__66405;
    wire N__66402;
    wire N__66401;
    wire N__66398;
    wire N__66395;
    wire N__66390;
    wire N__66387;
    wire N__66386;
    wire N__66383;
    wire N__66380;
    wire N__66375;
    wire N__66372;
    wire N__66371;
    wire N__66368;
    wire N__66367;
    wire N__66364;
    wire N__66361;
    wire N__66358;
    wire N__66355;
    wire N__66350;
    wire N__66345;
    wire N__66342;
    wire N__66341;
    wire N__66340;
    wire N__66337;
    wire N__66334;
    wire N__66331;
    wire N__66328;
    wire N__66321;
    wire N__66318;
    wire N__66317;
    wire N__66314;
    wire N__66313;
    wire N__66310;
    wire N__66307;
    wire N__66304;
    wire N__66299;
    wire N__66296;
    wire N__66291;
    wire N__66288;
    wire N__66287;
    wire N__66284;
    wire N__66283;
    wire N__66280;
    wire N__66277;
    wire N__66274;
    wire N__66267;
    wire N__66264;
    wire N__66263;
    wire N__66262;
    wire N__66259;
    wire N__66256;
    wire N__66253;
    wire N__66246;
    wire N__66243;
    wire N__66242;
    wire N__66241;
    wire N__66238;
    wire N__66235;
    wire N__66232;
    wire N__66225;
    wire N__66222;
    wire N__66221;
    wire N__66220;
    wire N__66217;
    wire N__66214;
    wire N__66211;
    wire N__66204;
    wire N__66201;
    wire N__66198;
    wire N__66195;
    wire N__66192;
    wire N__66189;
    wire N__66186;
    wire N__66183;
    wire N__66180;
    wire N__66177;
    wire N__66174;
    wire N__66173;
    wire N__66170;
    wire N__66167;
    wire N__66162;
    wire N__66159;
    wire N__66156;
    wire N__66153;
    wire N__66150;
    wire N__66147;
    wire N__66144;
    wire N__66141;
    wire N__66138;
    wire N__66135;
    wire N__66134;
    wire N__66133;
    wire N__66130;
    wire N__66127;
    wire N__66124;
    wire N__66121;
    wire N__66116;
    wire N__66113;
    wire N__66110;
    wire N__66105;
    wire N__66104;
    wire N__66101;
    wire N__66098;
    wire N__66095;
    wire N__66092;
    wire N__66089;
    wire N__66084;
    wire N__66083;
    wire N__66080;
    wire N__66079;
    wire N__66076;
    wire N__66075;
    wire N__66070;
    wire N__66067;
    wire N__66064;
    wire N__66057;
    wire N__66056;
    wire N__66053;
    wire N__66050;
    wire N__66047;
    wire N__66042;
    wire N__66041;
    wire N__66036;
    wire N__66033;
    wire N__66030;
    wire N__66027;
    wire N__66026;
    wire N__66025;
    wire N__66022;
    wire N__66019;
    wire N__66018;
    wire N__66017;
    wire N__66014;
    wire N__66011;
    wire N__66008;
    wire N__66005;
    wire N__66002;
    wire N__65999;
    wire N__65996;
    wire N__65991;
    wire N__65988;
    wire N__65979;
    wire N__65976;
    wire N__65973;
    wire N__65970;
    wire N__65967;
    wire N__65964;
    wire N__65961;
    wire N__65960;
    wire N__65957;
    wire N__65954;
    wire N__65949;
    wire N__65946;
    wire N__65943;
    wire N__65942;
    wire N__65939;
    wire N__65938;
    wire N__65937;
    wire N__65934;
    wire N__65931;
    wire N__65928;
    wire N__65925;
    wire N__65920;
    wire N__65917;
    wire N__65910;
    wire N__65907;
    wire N__65904;
    wire N__65901;
    wire N__65898;
    wire N__65895;
    wire N__65892;
    wire N__65891;
    wire N__65888;
    wire N__65885;
    wire N__65880;
    wire N__65879;
    wire N__65876;
    wire N__65875;
    wire N__65872;
    wire N__65869;
    wire N__65866;
    wire N__65863;
    wire N__65860;
    wire N__65857;
    wire N__65852;
    wire N__65847;
    wire N__65846;
    wire N__65843;
    wire N__65840;
    wire N__65837;
    wire N__65836;
    wire N__65833;
    wire N__65830;
    wire N__65827;
    wire N__65820;
    wire N__65817;
    wire N__65814;
    wire N__65811;
    wire N__65808;
    wire N__65805;
    wire N__65802;
    wire N__65799;
    wire N__65796;
    wire N__65793;
    wire N__65790;
    wire N__65787;
    wire N__65784;
    wire N__65781;
    wire N__65778;
    wire N__65775;
    wire N__65772;
    wire N__65771;
    wire N__65768;
    wire N__65765;
    wire N__65762;
    wire N__65761;
    wire N__65758;
    wire N__65755;
    wire N__65752;
    wire N__65745;
    wire N__65744;
    wire N__65739;
    wire N__65736;
    wire N__65735;
    wire N__65732;
    wire N__65731;
    wire N__65728;
    wire N__65723;
    wire N__65722;
    wire N__65719;
    wire N__65716;
    wire N__65713;
    wire N__65706;
    wire N__65703;
    wire N__65700;
    wire N__65697;
    wire N__65694;
    wire N__65691;
    wire N__65688;
    wire N__65685;
    wire N__65682;
    wire N__65679;
    wire N__65678;
    wire N__65677;
    wire N__65674;
    wire N__65673;
    wire N__65668;
    wire N__65665;
    wire N__65662;
    wire N__65659;
    wire N__65656;
    wire N__65653;
    wire N__65650;
    wire N__65647;
    wire N__65640;
    wire N__65639;
    wire N__65636;
    wire N__65633;
    wire N__65630;
    wire N__65627;
    wire N__65624;
    wire N__65621;
    wire N__65616;
    wire N__65613;
    wire N__65610;
    wire N__65607;
    wire N__65604;
    wire N__65601;
    wire N__65598;
    wire N__65595;
    wire N__65592;
    wire N__65589;
    wire N__65588;
    wire N__65585;
    wire N__65584;
    wire N__65581;
    wire N__65578;
    wire N__65575;
    wire N__65572;
    wire N__65569;
    wire N__65564;
    wire N__65559;
    wire N__65556;
    wire N__65553;
    wire N__65550;
    wire N__65549;
    wire N__65546;
    wire N__65543;
    wire N__65540;
    wire N__65535;
    wire N__65532;
    wire N__65529;
    wire N__65526;
    wire N__65525;
    wire N__65524;
    wire N__65523;
    wire N__65522;
    wire N__65521;
    wire N__65518;
    wire N__65511;
    wire N__65508;
    wire N__65505;
    wire N__65502;
    wire N__65499;
    wire N__65496;
    wire N__65493;
    wire N__65488;
    wire N__65485;
    wire N__65478;
    wire N__65475;
    wire N__65474;
    wire N__65473;
    wire N__65472;
    wire N__65471;
    wire N__65468;
    wire N__65465;
    wire N__65458;
    wire N__65455;
    wire N__65450;
    wire N__65445;
    wire N__65442;
    wire N__65439;
    wire N__65436;
    wire N__65435;
    wire N__65432;
    wire N__65429;
    wire N__65424;
    wire N__65421;
    wire N__65418;
    wire N__65415;
    wire N__65412;
    wire N__65411;
    wire N__65408;
    wire N__65405;
    wire N__65402;
    wire N__65399;
    wire N__65396;
    wire N__65393;
    wire N__65390;
    wire N__65387;
    wire N__65384;
    wire N__65379;
    wire N__65376;
    wire N__65373;
    wire N__65370;
    wire N__65367;
    wire N__65364;
    wire N__65363;
    wire N__65360;
    wire N__65357;
    wire N__65356;
    wire N__65351;
    wire N__65348;
    wire N__65345;
    wire N__65342;
    wire N__65339;
    wire N__65336;
    wire N__65331;
    wire N__65328;
    wire N__65325;
    wire N__65324;
    wire N__65321;
    wire N__65318;
    wire N__65317;
    wire N__65314;
    wire N__65309;
    wire N__65304;
    wire N__65301;
    wire N__65298;
    wire N__65295;
    wire N__65292;
    wire N__65289;
    wire N__65286;
    wire N__65283;
    wire N__65280;
    wire N__65277;
    wire N__65274;
    wire N__65273;
    wire N__65272;
    wire N__65269;
    wire N__65266;
    wire N__65263;
    wire N__65262;
    wire N__65259;
    wire N__65254;
    wire N__65251;
    wire N__65246;
    wire N__65243;
    wire N__65240;
    wire N__65235;
    wire N__65232;
    wire N__65229;
    wire N__65226;
    wire N__65223;
    wire N__65220;
    wire N__65217;
    wire N__65216;
    wire N__65213;
    wire N__65210;
    wire N__65205;
    wire N__65204;
    wire N__65201;
    wire N__65198;
    wire N__65193;
    wire N__65190;
    wire N__65187;
    wire N__65184;
    wire N__65181;
    wire N__65178;
    wire N__65175;
    wire N__65172;
    wire N__65169;
    wire N__65168;
    wire N__65165;
    wire N__65162;
    wire N__65159;
    wire N__65154;
    wire N__65151;
    wire N__65148;
    wire N__65147;
    wire N__65146;
    wire N__65145;
    wire N__65142;
    wire N__65139;
    wire N__65138;
    wire N__65137;
    wire N__65136;
    wire N__65135;
    wire N__65130;
    wire N__65127;
    wire N__65124;
    wire N__65123;
    wire N__65122;
    wire N__65121;
    wire N__65116;
    wire N__65111;
    wire N__65104;
    wire N__65097;
    wire N__65088;
    wire N__65085;
    wire N__65082;
    wire N__65081;
    wire N__65080;
    wire N__65079;
    wire N__65078;
    wire N__65077;
    wire N__65076;
    wire N__65075;
    wire N__65074;
    wire N__65073;
    wire N__65070;
    wire N__65063;
    wire N__65058;
    wire N__65053;
    wire N__65048;
    wire N__65037;
    wire N__65036;
    wire N__65033;
    wire N__65030;
    wire N__65025;
    wire N__65022;
    wire N__65019;
    wire N__65016;
    wire N__65013;
    wire N__65010;
    wire N__65007;
    wire N__65004;
    wire N__65001;
    wire N__65000;
    wire N__64999;
    wire N__64998;
    wire N__64997;
    wire N__64996;
    wire N__64995;
    wire N__64994;
    wire N__64993;
    wire N__64990;
    wire N__64989;
    wire N__64986;
    wire N__64985;
    wire N__64982;
    wire N__64981;
    wire N__64978;
    wire N__64977;
    wire N__64974;
    wire N__64973;
    wire N__64970;
    wire N__64969;
    wire N__64966;
    wire N__64965;
    wire N__64962;
    wire N__64961;
    wire N__64960;
    wire N__64959;
    wire N__64958;
    wire N__64957;
    wire N__64954;
    wire N__64937;
    wire N__64920;
    wire N__64917;
    wire N__64916;
    wire N__64913;
    wire N__64912;
    wire N__64909;
    wire N__64908;
    wire N__64905;
    wire N__64904;
    wire N__64903;
    wire N__64896;
    wire N__64879;
    wire N__64878;
    wire N__64877;
    wire N__64876;
    wire N__64873;
    wire N__64872;
    wire N__64871;
    wire N__64870;
    wire N__64869;
    wire N__64864;
    wire N__64855;
    wire N__64846;
    wire N__64839;
    wire N__64836;
    wire N__64833;
    wire N__64830;
    wire N__64829;
    wire N__64828;
    wire N__64827;
    wire N__64826;
    wire N__64825;
    wire N__64822;
    wire N__64819;
    wire N__64816;
    wire N__64813;
    wire N__64810;
    wire N__64807;
    wire N__64804;
    wire N__64801;
    wire N__64794;
    wire N__64791;
    wire N__64788;
    wire N__64783;
    wire N__64776;
    wire N__64773;
    wire N__64770;
    wire N__64767;
    wire N__64764;
    wire N__64761;
    wire N__64758;
    wire N__64755;
    wire N__64754;
    wire N__64751;
    wire N__64748;
    wire N__64745;
    wire N__64740;
    wire N__64739;
    wire N__64738;
    wire N__64735;
    wire N__64732;
    wire N__64731;
    wire N__64728;
    wire N__64725;
    wire N__64722;
    wire N__64719;
    wire N__64716;
    wire N__64713;
    wire N__64712;
    wire N__64711;
    wire N__64706;
    wire N__64701;
    wire N__64698;
    wire N__64695;
    wire N__64692;
    wire N__64683;
    wire N__64680;
    wire N__64677;
    wire N__64674;
    wire N__64671;
    wire N__64668;
    wire N__64665;
    wire N__64662;
    wire N__64659;
    wire N__64656;
    wire N__64653;
    wire N__64650;
    wire N__64647;
    wire N__64644;
    wire N__64641;
    wire N__64638;
    wire N__64635;
    wire N__64632;
    wire N__64629;
    wire N__64626;
    wire N__64623;
    wire N__64620;
    wire N__64617;
    wire N__64614;
    wire N__64611;
    wire N__64608;
    wire N__64605;
    wire N__64602;
    wire N__64599;
    wire N__64596;
    wire N__64593;
    wire N__64590;
    wire N__64587;
    wire N__64584;
    wire N__64581;
    wire N__64578;
    wire N__64575;
    wire N__64572;
    wire N__64569;
    wire N__64566;
    wire N__64563;
    wire N__64560;
    wire N__64559;
    wire N__64558;
    wire N__64555;
    wire N__64552;
    wire N__64549;
    wire N__64542;
    wire N__64541;
    wire N__64538;
    wire N__64537;
    wire N__64534;
    wire N__64531;
    wire N__64528;
    wire N__64521;
    wire N__64518;
    wire N__64515;
    wire N__64514;
    wire N__64513;
    wire N__64512;
    wire N__64511;
    wire N__64510;
    wire N__64509;
    wire N__64508;
    wire N__64505;
    wire N__64502;
    wire N__64499;
    wire N__64496;
    wire N__64493;
    wire N__64490;
    wire N__64487;
    wire N__64484;
    wire N__64477;
    wire N__64472;
    wire N__64465;
    wire N__64460;
    wire N__64455;
    wire N__64452;
    wire N__64451;
    wire N__64450;
    wire N__64449;
    wire N__64448;
    wire N__64447;
    wire N__64444;
    wire N__64441;
    wire N__64438;
    wire N__64435;
    wire N__64432;
    wire N__64429;
    wire N__64424;
    wire N__64415;
    wire N__64410;
    wire N__64407;
    wire N__64406;
    wire N__64405;
    wire N__64402;
    wire N__64399;
    wire N__64396;
    wire N__64393;
    wire N__64390;
    wire N__64383;
    wire N__64382;
    wire N__64381;
    wire N__64378;
    wire N__64375;
    wire N__64372;
    wire N__64369;
    wire N__64362;
    wire N__64359;
    wire N__64356;
    wire N__64353;
    wire N__64352;
    wire N__64351;
    wire N__64348;
    wire N__64345;
    wire N__64342;
    wire N__64339;
    wire N__64332;
    wire N__64331;
    wire N__64330;
    wire N__64327;
    wire N__64324;
    wire N__64321;
    wire N__64318;
    wire N__64311;
    wire N__64310;
    wire N__64309;
    wire N__64306;
    wire N__64303;
    wire N__64300;
    wire N__64297;
    wire N__64290;
    wire N__64287;
    wire N__64286;
    wire N__64285;
    wire N__64282;
    wire N__64279;
    wire N__64276;
    wire N__64269;
    wire N__64266;
    wire N__64263;
    wire N__64260;
    wire N__64257;
    wire N__64254;
    wire N__64251;
    wire N__64248;
    wire N__64245;
    wire N__64242;
    wire N__64239;
    wire N__64236;
    wire N__64233;
    wire N__64230;
    wire N__64227;
    wire N__64226;
    wire N__64225;
    wire N__64224;
    wire N__64223;
    wire N__64222;
    wire N__64219;
    wire N__64216;
    wire N__64213;
    wire N__64210;
    wire N__64207;
    wire N__64204;
    wire N__64199;
    wire N__64190;
    wire N__64185;
    wire N__64182;
    wire N__64179;
    wire N__64176;
    wire N__64175;
    wire N__64174;
    wire N__64171;
    wire N__64168;
    wire N__64165;
    wire N__64160;
    wire N__64157;
    wire N__64154;
    wire N__64149;
    wire N__64146;
    wire N__64145;
    wire N__64144;
    wire N__64141;
    wire N__64138;
    wire N__64135;
    wire N__64132;
    wire N__64127;
    wire N__64124;
    wire N__64119;
    wire N__64116;
    wire N__64113;
    wire N__64110;
    wire N__64109;
    wire N__64108;
    wire N__64105;
    wire N__64102;
    wire N__64099;
    wire N__64096;
    wire N__64093;
    wire N__64088;
    wire N__64083;
    wire N__64080;
    wire N__64079;
    wire N__64078;
    wire N__64075;
    wire N__64072;
    wire N__64069;
    wire N__64066;
    wire N__64061;
    wire N__64058;
    wire N__64053;
    wire N__64050;
    wire N__64049;
    wire N__64048;
    wire N__64045;
    wire N__64042;
    wire N__64039;
    wire N__64036;
    wire N__64031;
    wire N__64028;
    wire N__64023;
    wire N__64020;
    wire N__64019;
    wire N__64018;
    wire N__64015;
    wire N__64012;
    wire N__64009;
    wire N__64006;
    wire N__64003;
    wire N__64000;
    wire N__63997;
    wire N__63990;
    wire N__63989;
    wire N__63988;
    wire N__63987;
    wire N__63986;
    wire N__63983;
    wire N__63980;
    wire N__63977;
    wire N__63974;
    wire N__63971;
    wire N__63970;
    wire N__63969;
    wire N__63964;
    wire N__63957;
    wire N__63954;
    wire N__63951;
    wire N__63946;
    wire N__63941;
    wire N__63938;
    wire N__63935;
    wire N__63930;
    wire N__63927;
    wire N__63926;
    wire N__63925;
    wire N__63922;
    wire N__63921;
    wire N__63918;
    wire N__63915;
    wire N__63912;
    wire N__63909;
    wire N__63904;
    wire N__63901;
    wire N__63894;
    wire N__63893;
    wire N__63892;
    wire N__63889;
    wire N__63886;
    wire N__63883;
    wire N__63876;
    wire N__63875;
    wire N__63874;
    wire N__63871;
    wire N__63868;
    wire N__63865;
    wire N__63858;
    wire N__63857;
    wire N__63856;
    wire N__63853;
    wire N__63850;
    wire N__63847;
    wire N__63840;
    wire N__63839;
    wire N__63838;
    wire N__63835;
    wire N__63832;
    wire N__63829;
    wire N__63826;
    wire N__63819;
    wire N__63818;
    wire N__63817;
    wire N__63814;
    wire N__63811;
    wire N__63808;
    wire N__63801;
    wire N__63800;
    wire N__63797;
    wire N__63794;
    wire N__63793;
    wire N__63788;
    wire N__63785;
    wire N__63780;
    wire N__63777;
    wire N__63776;
    wire N__63773;
    wire N__63770;
    wire N__63769;
    wire N__63764;
    wire N__63761;
    wire N__63756;
    wire N__63755;
    wire N__63754;
    wire N__63753;
    wire N__63750;
    wire N__63747;
    wire N__63744;
    wire N__63741;
    wire N__63740;
    wire N__63739;
    wire N__63734;
    wire N__63729;
    wire N__63726;
    wire N__63723;
    wire N__63718;
    wire N__63713;
    wire N__63708;
    wire N__63705;
    wire N__63704;
    wire N__63701;
    wire N__63698;
    wire N__63697;
    wire N__63692;
    wire N__63689;
    wire N__63688;
    wire N__63685;
    wire N__63682;
    wire N__63679;
    wire N__63676;
    wire N__63673;
    wire N__63666;
    wire N__63663;
    wire N__63662;
    wire N__63659;
    wire N__63658;
    wire N__63655;
    wire N__63652;
    wire N__63649;
    wire N__63646;
    wire N__63643;
    wire N__63640;
    wire N__63637;
    wire N__63634;
    wire N__63627;
    wire N__63624;
    wire N__63623;
    wire N__63622;
    wire N__63619;
    wire N__63616;
    wire N__63613;
    wire N__63610;
    wire N__63607;
    wire N__63604;
    wire N__63597;
    wire N__63594;
    wire N__63591;
    wire N__63588;
    wire N__63587;
    wire N__63586;
    wire N__63583;
    wire N__63580;
    wire N__63577;
    wire N__63574;
    wire N__63569;
    wire N__63566;
    wire N__63561;
    wire N__63558;
    wire N__63555;
    wire N__63552;
    wire N__63551;
    wire N__63550;
    wire N__63547;
    wire N__63544;
    wire N__63541;
    wire N__63538;
    wire N__63531;
    wire N__63528;
    wire N__63525;
    wire N__63524;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63514;
    wire N__63511;
    wire N__63508;
    wire N__63505;
    wire N__63502;
    wire N__63495;
    wire N__63492;
    wire N__63489;
    wire N__63488;
    wire N__63487;
    wire N__63484;
    wire N__63481;
    wire N__63478;
    wire N__63475;
    wire N__63472;
    wire N__63469;
    wire N__63466;
    wire N__63459;
    wire N__63456;
    wire N__63455;
    wire N__63454;
    wire N__63451;
    wire N__63448;
    wire N__63445;
    wire N__63442;
    wire N__63437;
    wire N__63434;
    wire N__63429;
    wire N__63426;
    wire N__63425;
    wire N__63424;
    wire N__63421;
    wire N__63418;
    wire N__63415;
    wire N__63412;
    wire N__63409;
    wire N__63406;
    wire N__63403;
    wire N__63396;
    wire N__63393;
    wire N__63392;
    wire N__63391;
    wire N__63388;
    wire N__63385;
    wire N__63382;
    wire N__63379;
    wire N__63374;
    wire N__63371;
    wire N__63366;
    wire N__63365;
    wire N__63364;
    wire N__63363;
    wire N__63362;
    wire N__63361;
    wire N__63358;
    wire N__63355;
    wire N__63352;
    wire N__63349;
    wire N__63346;
    wire N__63343;
    wire N__63338;
    wire N__63329;
    wire N__63324;
    wire N__63321;
    wire N__63320;
    wire N__63319;
    wire N__63316;
    wire N__63313;
    wire N__63310;
    wire N__63307;
    wire N__63304;
    wire N__63301;
    wire N__63298;
    wire N__63291;
    wire N__63288;
    wire N__63287;
    wire N__63286;
    wire N__63283;
    wire N__63280;
    wire N__63277;
    wire N__63272;
    wire N__63269;
    wire N__63264;
    wire N__63261;
    wire N__63260;
    wire N__63259;
    wire N__63256;
    wire N__63253;
    wire N__63250;
    wire N__63245;
    wire N__63242;
    wire N__63237;
    wire N__63234;
    wire N__63233;
    wire N__63232;
    wire N__63229;
    wire N__63226;
    wire N__63223;
    wire N__63218;
    wire N__63215;
    wire N__63212;
    wire N__63209;
    wire N__63204;
    wire N__63201;
    wire N__63200;
    wire N__63199;
    wire N__63196;
    wire N__63193;
    wire N__63190;
    wire N__63187;
    wire N__63184;
    wire N__63181;
    wire N__63176;
    wire N__63173;
    wire N__63168;
    wire N__63165;
    wire N__63164;
    wire N__63161;
    wire N__63160;
    wire N__63157;
    wire N__63154;
    wire N__63151;
    wire N__63148;
    wire N__63145;
    wire N__63142;
    wire N__63137;
    wire N__63134;
    wire N__63129;
    wire N__63128;
    wire N__63127;
    wire N__63124;
    wire N__63121;
    wire N__63118;
    wire N__63117;
    wire N__63116;
    wire N__63113;
    wire N__63108;
    wire N__63105;
    wire N__63102;
    wire N__63097;
    wire N__63092;
    wire N__63087;
    wire N__63084;
    wire N__63081;
    wire N__63078;
    wire N__63075;
    wire N__63072;
    wire N__63069;
    wire N__63066;
    wire N__63063;
    wire N__63060;
    wire N__63057;
    wire N__63054;
    wire N__63053;
    wire N__63052;
    wire N__63049;
    wire N__63048;
    wire N__63045;
    wire N__63042;
    wire N__63039;
    wire N__63036;
    wire N__63027;
    wire N__63024;
    wire N__63023;
    wire N__63020;
    wire N__63017;
    wire N__63016;
    wire N__63011;
    wire N__63008;
    wire N__63003;
    wire N__63000;
    wire N__62999;
    wire N__62998;
    wire N__62997;
    wire N__62994;
    wire N__62991;
    wire N__62988;
    wire N__62985;
    wire N__62982;
    wire N__62973;
    wire N__62970;
    wire N__62969;
    wire N__62966;
    wire N__62963;
    wire N__62958;
    wire N__62957;
    wire N__62954;
    wire N__62951;
    wire N__62946;
    wire N__62943;
    wire N__62940;
    wire N__62939;
    wire N__62938;
    wire N__62935;
    wire N__62932;
    wire N__62929;
    wire N__62926;
    wire N__62923;
    wire N__62920;
    wire N__62915;
    wire N__62912;
    wire N__62907;
    wire N__62904;
    wire N__62903;
    wire N__62902;
    wire N__62899;
    wire N__62896;
    wire N__62893;
    wire N__62890;
    wire N__62887;
    wire N__62882;
    wire N__62879;
    wire N__62876;
    wire N__62871;
    wire N__62868;
    wire N__62867;
    wire N__62866;
    wire N__62863;
    wire N__62860;
    wire N__62857;
    wire N__62854;
    wire N__62849;
    wire N__62844;
    wire N__62841;
    wire N__62838;
    wire N__62837;
    wire N__62836;
    wire N__62833;
    wire N__62830;
    wire N__62827;
    wire N__62822;
    wire N__62819;
    wire N__62816;
    wire N__62813;
    wire N__62808;
    wire N__62805;
    wire N__62804;
    wire N__62803;
    wire N__62800;
    wire N__62797;
    wire N__62794;
    wire N__62791;
    wire N__62788;
    wire N__62785;
    wire N__62780;
    wire N__62777;
    wire N__62772;
    wire N__62771;
    wire N__62770;
    wire N__62769;
    wire N__62768;
    wire N__62767;
    wire N__62764;
    wire N__62761;
    wire N__62758;
    wire N__62755;
    wire N__62752;
    wire N__62749;
    wire N__62744;
    wire N__62735;
    wire N__62730;
    wire N__62727;
    wire N__62726;
    wire N__62725;
    wire N__62722;
    wire N__62719;
    wire N__62716;
    wire N__62711;
    wire N__62708;
    wire N__62705;
    wire N__62702;
    wire N__62697;
    wire N__62694;
    wire N__62691;
    wire N__62688;
    wire N__62685;
    wire N__62682;
    wire N__62679;
    wire N__62676;
    wire N__62673;
    wire N__62670;
    wire N__62667;
    wire N__62664;
    wire N__62661;
    wire N__62658;
    wire N__62655;
    wire N__62652;
    wire N__62649;
    wire N__62646;
    wire N__62643;
    wire N__62640;
    wire N__62637;
    wire N__62634;
    wire N__62631;
    wire N__62628;
    wire N__62625;
    wire N__62622;
    wire N__62619;
    wire N__62618;
    wire N__62615;
    wire N__62612;
    wire N__62611;
    wire N__62610;
    wire N__62609;
    wire N__62608;
    wire N__62607;
    wire N__62606;
    wire N__62605;
    wire N__62604;
    wire N__62601;
    wire N__62598;
    wire N__62595;
    wire N__62592;
    wire N__62589;
    wire N__62586;
    wire N__62583;
    wire N__62580;
    wire N__62577;
    wire N__62574;
    wire N__62573;
    wire N__62572;
    wire N__62567;
    wire N__62558;
    wire N__62549;
    wire N__62546;
    wire N__62543;
    wire N__62536;
    wire N__62531;
    wire N__62526;
    wire N__62523;
    wire N__62520;
    wire N__62517;
    wire N__62514;
    wire N__62511;
    wire N__62508;
    wire N__62505;
    wire N__62504;
    wire N__62501;
    wire N__62498;
    wire N__62497;
    wire N__62496;
    wire N__62495;
    wire N__62494;
    wire N__62489;
    wire N__62486;
    wire N__62483;
    wire N__62480;
    wire N__62477;
    wire N__62474;
    wire N__62465;
    wire N__62460;
    wire N__62457;
    wire N__62454;
    wire N__62451;
    wire N__62448;
    wire N__62447;
    wire N__62444;
    wire N__62441;
    wire N__62438;
    wire N__62435;
    wire N__62432;
    wire N__62431;
    wire N__62426;
    wire N__62423;
    wire N__62420;
    wire N__62415;
    wire N__62412;
    wire N__62411;
    wire N__62408;
    wire N__62407;
    wire N__62404;
    wire N__62401;
    wire N__62398;
    wire N__62395;
    wire N__62388;
    wire N__62385;
    wire N__62382;
    wire N__62379;
    wire N__62376;
    wire N__62373;
    wire N__62370;
    wire N__62367;
    wire N__62364;
    wire N__62361;
    wire N__62358;
    wire N__62355;
    wire N__62352;
    wire N__62349;
    wire N__62346;
    wire N__62345;
    wire N__62342;
    wire N__62339;
    wire N__62336;
    wire N__62333;
    wire N__62330;
    wire N__62325;
    wire N__62324;
    wire N__62321;
    wire N__62320;
    wire N__62317;
    wire N__62316;
    wire N__62313;
    wire N__62310;
    wire N__62309;
    wire N__62306;
    wire N__62303;
    wire N__62300;
    wire N__62297;
    wire N__62294;
    wire N__62291;
    wire N__62284;
    wire N__62281;
    wire N__62278;
    wire N__62275;
    wire N__62268;
    wire N__62267;
    wire N__62266;
    wire N__62265;
    wire N__62262;
    wire N__62261;
    wire N__62260;
    wire N__62259;
    wire N__62258;
    wire N__62255;
    wire N__62254;
    wire N__62253;
    wire N__62250;
    wire N__62247;
    wire N__62246;
    wire N__62245;
    wire N__62242;
    wire N__62241;
    wire N__62240;
    wire N__62239;
    wire N__62236;
    wire N__62233;
    wire N__62230;
    wire N__62229;
    wire N__62226;
    wire N__62225;
    wire N__62224;
    wire N__62221;
    wire N__62218;
    wire N__62215;
    wire N__62212;
    wire N__62205;
    wire N__62202;
    wire N__62199;
    wire N__62196;
    wire N__62193;
    wire N__62188;
    wire N__62185;
    wire N__62182;
    wire N__62179;
    wire N__62178;
    wire N__62177;
    wire N__62174;
    wire N__62173;
    wire N__62172;
    wire N__62169;
    wire N__62166;
    wire N__62163;
    wire N__62160;
    wire N__62155;
    wire N__62150;
    wire N__62149;
    wire N__62144;
    wire N__62141;
    wire N__62134;
    wire N__62131;
    wire N__62130;
    wire N__62127;
    wire N__62124;
    wire N__62119;
    wire N__62114;
    wire N__62109;
    wire N__62106;
    wire N__62103;
    wire N__62100;
    wire N__62095;
    wire N__62092;
    wire N__62087;
    wire N__62072;
    wire N__62071;
    wire N__62066;
    wire N__62063;
    wire N__62058;
    wire N__62055;
    wire N__62050;
    wire N__62045;
    wire N__62040;
    wire N__62039;
    wire N__62036;
    wire N__62033;
    wire N__62030;
    wire N__62027;
    wire N__62026;
    wire N__62025;
    wire N__62022;
    wire N__62019;
    wire N__62014;
    wire N__62007;
    wire N__62004;
    wire N__62003;
    wire N__62000;
    wire N__61999;
    wire N__61996;
    wire N__61993;
    wire N__61992;
    wire N__61989;
    wire N__61986;
    wire N__61983;
    wire N__61980;
    wire N__61977;
    wire N__61972;
    wire N__61965;
    wire N__61962;
    wire N__61961;
    wire N__61960;
    wire N__61959;
    wire N__61958;
    wire N__61957;
    wire N__61956;
    wire N__61955;
    wire N__61954;
    wire N__61951;
    wire N__61950;
    wire N__61947;
    wire N__61946;
    wire N__61943;
    wire N__61942;
    wire N__61939;
    wire N__61938;
    wire N__61937;
    wire N__61934;
    wire N__61933;
    wire N__61930;
    wire N__61929;
    wire N__61926;
    wire N__61925;
    wire N__61922;
    wire N__61921;
    wire N__61920;
    wire N__61919;
    wire N__61918;
    wire N__61917;
    wire N__61916;
    wire N__61915;
    wire N__61914;
    wire N__61911;
    wire N__61894;
    wire N__61877;
    wire N__61874;
    wire N__61873;
    wire N__61870;
    wire N__61869;
    wire N__61866;
    wire N__61865;
    wire N__61862;
    wire N__61861;
    wire N__61858;
    wire N__61855;
    wire N__61854;
    wire N__61851;
    wire N__61850;
    wire N__61847;
    wire N__61846;
    wire N__61845;
    wire N__61838;
    wire N__61821;
    wire N__61818;
    wire N__61803;
    wire N__61798;
    wire N__61793;
    wire N__61790;
    wire N__61787;
    wire N__61784;
    wire N__61781;
    wire N__61776;
    wire N__61773;
    wire N__61770;
    wire N__61767;
    wire N__61764;
    wire N__61761;
    wire N__61758;
    wire N__61755;
    wire N__61752;
    wire N__61749;
    wire N__61746;
    wire N__61743;
    wire N__61740;
    wire N__61739;
    wire N__61736;
    wire N__61733;
    wire N__61730;
    wire N__61727;
    wire N__61722;
    wire N__61721;
    wire N__61720;
    wire N__61719;
    wire N__61716;
    wire N__61711;
    wire N__61708;
    wire N__61701;
    wire N__61700;
    wire N__61699;
    wire N__61698;
    wire N__61695;
    wire N__61690;
    wire N__61687;
    wire N__61684;
    wire N__61679;
    wire N__61674;
    wire N__61671;
    wire N__61670;
    wire N__61667;
    wire N__61664;
    wire N__61663;
    wire N__61660;
    wire N__61659;
    wire N__61656;
    wire N__61653;
    wire N__61650;
    wire N__61647;
    wire N__61638;
    wire N__61635;
    wire N__61632;
    wire N__61631;
    wire N__61628;
    wire N__61625;
    wire N__61620;
    wire N__61617;
    wire N__61616;
    wire N__61615;
    wire N__61612;
    wire N__61609;
    wire N__61608;
    wire N__61605;
    wire N__61600;
    wire N__61597;
    wire N__61592;
    wire N__61587;
    wire N__61584;
    wire N__61581;
    wire N__61578;
    wire N__61575;
    wire N__61572;
    wire N__61569;
    wire N__61566;
    wire N__61563;
    wire N__61560;
    wire N__61557;
    wire N__61554;
    wire N__61551;
    wire N__61548;
    wire N__61545;
    wire N__61542;
    wire N__61539;
    wire N__61536;
    wire N__61533;
    wire N__61530;
    wire N__61527;
    wire N__61524;
    wire N__61521;
    wire N__61518;
    wire N__61515;
    wire N__61512;
    wire N__61509;
    wire N__61506;
    wire N__61503;
    wire N__61500;
    wire N__61497;
    wire N__61494;
    wire N__61491;
    wire N__61488;
    wire N__61485;
    wire N__61482;
    wire N__61479;
    wire N__61476;
    wire N__61473;
    wire N__61470;
    wire N__61467;
    wire N__61464;
    wire N__61461;
    wire N__61458;
    wire N__61457;
    wire N__61454;
    wire N__61453;
    wire N__61452;
    wire N__61449;
    wire N__61444;
    wire N__61441;
    wire N__61440;
    wire N__61439;
    wire N__61438;
    wire N__61437;
    wire N__61430;
    wire N__61425;
    wire N__61422;
    wire N__61419;
    wire N__61416;
    wire N__61411;
    wire N__61408;
    wire N__61405;
    wire N__61402;
    wire N__61395;
    wire N__61392;
    wire N__61391;
    wire N__61388;
    wire N__61385;
    wire N__61382;
    wire N__61377;
    wire N__61376;
    wire N__61373;
    wire N__61370;
    wire N__61367;
    wire N__61362;
    wire N__61359;
    wire N__61356;
    wire N__61353;
    wire N__61350;
    wire N__61347;
    wire N__61344;
    wire N__61341;
    wire N__61340;
    wire N__61337;
    wire N__61334;
    wire N__61331;
    wire N__61328;
    wire N__61325;
    wire N__61320;
    wire N__61319;
    wire N__61314;
    wire N__61311;
    wire N__61308;
    wire N__61305;
    wire N__61304;
    wire N__61299;
    wire N__61296;
    wire N__61293;
    wire N__61290;
    wire N__61287;
    wire N__61286;
    wire N__61283;
    wire N__61280;
    wire N__61277;
    wire N__61272;
    wire N__61269;
    wire N__61266;
    wire N__61263;
    wire N__61260;
    wire N__61257;
    wire N__61254;
    wire N__61251;
    wire N__61248;
    wire N__61247;
    wire N__61244;
    wire N__61241;
    wire N__61238;
    wire N__61233;
    wire N__61230;
    wire N__61227;
    wire N__61226;
    wire N__61223;
    wire N__61220;
    wire N__61215;
    wire N__61214;
    wire N__61211;
    wire N__61210;
    wire N__61209;
    wire N__61206;
    wire N__61203;
    wire N__61200;
    wire N__61197;
    wire N__61190;
    wire N__61185;
    wire N__61184;
    wire N__61181;
    wire N__61178;
    wire N__61177;
    wire N__61176;
    wire N__61173;
    wire N__61170;
    wire N__61167;
    wire N__61164;
    wire N__61161;
    wire N__61158;
    wire N__61155;
    wire N__61152;
    wire N__61149;
    wire N__61146;
    wire N__61143;
    wire N__61140;
    wire N__61137;
    wire N__61134;
    wire N__61129;
    wire N__61122;
    wire N__61119;
    wire N__61118;
    wire N__61115;
    wire N__61112;
    wire N__61107;
    wire N__61106;
    wire N__61103;
    wire N__61100;
    wire N__61095;
    wire N__61092;
    wire N__61091;
    wire N__61088;
    wire N__61085;
    wire N__61082;
    wire N__61077;
    wire N__61074;
    wire N__61071;
    wire N__61070;
    wire N__61067;
    wire N__61064;
    wire N__61059;
    wire N__61058;
    wire N__61055;
    wire N__61052;
    wire N__61047;
    wire N__61044;
    wire N__61041;
    wire N__61038;
    wire N__61035;
    wire N__61034;
    wire N__61031;
    wire N__61028;
    wire N__61023;
    wire N__61020;
    wire N__61017;
    wire N__61016;
    wire N__61013;
    wire N__61010;
    wire N__61005;
    wire N__61004;
    wire N__60999;
    wire N__60996;
    wire N__60993;
    wire N__60992;
    wire N__60987;
    wire N__60984;
    wire N__60981;
    wire N__60978;
    wire N__60975;
    wire N__60972;
    wire N__60969;
    wire N__60966;
    wire N__60963;
    wire N__60960;
    wire N__60957;
    wire N__60954;
    wire N__60951;
    wire N__60948;
    wire N__60947;
    wire N__60944;
    wire N__60941;
    wire N__60936;
    wire N__60935;
    wire N__60932;
    wire N__60929;
    wire N__60924;
    wire N__60923;
    wire N__60920;
    wire N__60917;
    wire N__60912;
    wire N__60911;
    wire N__60908;
    wire N__60905;
    wire N__60904;
    wire N__60899;
    wire N__60896;
    wire N__60893;
    wire N__60890;
    wire N__60885;
    wire N__60882;
    wire N__60881;
    wire N__60878;
    wire N__60875;
    wire N__60870;
    wire N__60869;
    wire N__60866;
    wire N__60863;
    wire N__60858;
    wire N__60855;
    wire N__60854;
    wire N__60851;
    wire N__60848;
    wire N__60843;
    wire N__60842;
    wire N__60839;
    wire N__60836;
    wire N__60831;
    wire N__60828;
    wire N__60827;
    wire N__60826;
    wire N__60823;
    wire N__60820;
    wire N__60817;
    wire N__60810;
    wire N__60807;
    wire N__60804;
    wire N__60801;
    wire N__60798;
    wire N__60797;
    wire N__60794;
    wire N__60791;
    wire N__60786;
    wire N__60785;
    wire N__60782;
    wire N__60779;
    wire N__60774;
    wire N__60773;
    wire N__60768;
    wire N__60765;
    wire N__60762;
    wire N__60759;
    wire N__60756;
    wire N__60753;
    wire N__60752;
    wire N__60749;
    wire N__60746;
    wire N__60741;
    wire N__60740;
    wire N__60737;
    wire N__60734;
    wire N__60729;
    wire N__60726;
    wire N__60725;
    wire N__60722;
    wire N__60719;
    wire N__60716;
    wire N__60713;
    wire N__60712;
    wire N__60707;
    wire N__60704;
    wire N__60699;
    wire N__60696;
    wire N__60695;
    wire N__60692;
    wire N__60689;
    wire N__60684;
    wire N__60683;
    wire N__60680;
    wire N__60677;
    wire N__60672;
    wire N__60669;
    wire N__60668;
    wire N__60665;
    wire N__60662;
    wire N__60661;
    wire N__60656;
    wire N__60653;
    wire N__60650;
    wire N__60647;
    wire N__60642;
    wire N__60639;
    wire N__60638;
    wire N__60635;
    wire N__60632;
    wire N__60627;
    wire N__60626;
    wire N__60623;
    wire N__60620;
    wire N__60615;
    wire N__60612;
    wire N__60611;
    wire N__60610;
    wire N__60607;
    wire N__60604;
    wire N__60601;
    wire N__60596;
    wire N__60593;
    wire N__60590;
    wire N__60587;
    wire N__60582;
    wire N__60579;
    wire N__60578;
    wire N__60575;
    wire N__60572;
    wire N__60571;
    wire N__60566;
    wire N__60563;
    wire N__60560;
    wire N__60557;
    wire N__60552;
    wire N__60549;
    wire N__60548;
    wire N__60545;
    wire N__60542;
    wire N__60537;
    wire N__60536;
    wire N__60533;
    wire N__60530;
    wire N__60525;
    wire N__60522;
    wire N__60519;
    wire N__60518;
    wire N__60515;
    wire N__60512;
    wire N__60511;
    wire N__60506;
    wire N__60503;
    wire N__60502;
    wire N__60499;
    wire N__60496;
    wire N__60493;
    wire N__60490;
    wire N__60487;
    wire N__60480;
    wire N__60477;
    wire N__60476;
    wire N__60475;
    wire N__60472;
    wire N__60469;
    wire N__60466;
    wire N__60461;
    wire N__60458;
    wire N__60457;
    wire N__60454;
    wire N__60451;
    wire N__60448;
    wire N__60443;
    wire N__60438;
    wire N__60435;
    wire N__60434;
    wire N__60433;
    wire N__60430;
    wire N__60427;
    wire N__60424;
    wire N__60421;
    wire N__60416;
    wire N__60413;
    wire N__60412;
    wire N__60407;
    wire N__60404;
    wire N__60401;
    wire N__60396;
    wire N__60393;
    wire N__60392;
    wire N__60391;
    wire N__60388;
    wire N__60385;
    wire N__60382;
    wire N__60379;
    wire N__60376;
    wire N__60373;
    wire N__60372;
    wire N__60365;
    wire N__60362;
    wire N__60359;
    wire N__60354;
    wire N__60351;
    wire N__60350;
    wire N__60349;
    wire N__60346;
    wire N__60343;
    wire N__60340;
    wire N__60335;
    wire N__60332;
    wire N__60331;
    wire N__60326;
    wire N__60323;
    wire N__60320;
    wire N__60315;
    wire N__60312;
    wire N__60309;
    wire N__60308;
    wire N__60307;
    wire N__60304;
    wire N__60301;
    wire N__60298;
    wire N__60293;
    wire N__60290;
    wire N__60289;
    wire N__60284;
    wire N__60281;
    wire N__60278;
    wire N__60273;
    wire N__60272;
    wire N__60269;
    wire N__60266;
    wire N__60263;
    wire N__60260;
    wire N__60257;
    wire N__60252;
    wire N__60249;
    wire N__60248;
    wire N__60245;
    wire N__60242;
    wire N__60239;
    wire N__60234;
    wire N__60233;
    wire N__60230;
    wire N__60227;
    wire N__60226;
    wire N__60221;
    wire N__60218;
    wire N__60215;
    wire N__60212;
    wire N__60207;
    wire N__60204;
    wire N__60203;
    wire N__60202;
    wire N__60199;
    wire N__60196;
    wire N__60195;
    wire N__60192;
    wire N__60189;
    wire N__60186;
    wire N__60183;
    wire N__60180;
    wire N__60177;
    wire N__60174;
    wire N__60169;
    wire N__60162;
    wire N__60159;
    wire N__60156;
    wire N__60153;
    wire N__60150;
    wire N__60147;
    wire N__60146;
    wire N__60145;
    wire N__60142;
    wire N__60139;
    wire N__60136;
    wire N__60135;
    wire N__60130;
    wire N__60127;
    wire N__60124;
    wire N__60119;
    wire N__60114;
    wire N__60111;
    wire N__60108;
    wire N__60107;
    wire N__60106;
    wire N__60103;
    wire N__60100;
    wire N__60097;
    wire N__60094;
    wire N__60093;
    wire N__60088;
    wire N__60085;
    wire N__60082;
    wire N__60079;
    wire N__60076;
    wire N__60071;
    wire N__60066;
    wire N__60063;
    wire N__60062;
    wire N__60061;
    wire N__60058;
    wire N__60055;
    wire N__60052;
    wire N__60045;
    wire N__60044;
    wire N__60041;
    wire N__60038;
    wire N__60035;
    wire N__60030;
    wire N__60027;
    wire N__60026;
    wire N__60025;
    wire N__60022;
    wire N__60019;
    wire N__60016;
    wire N__60011;
    wire N__60008;
    wire N__60007;
    wire N__60004;
    wire N__60001;
    wire N__59998;
    wire N__59995;
    wire N__59992;
    wire N__59985;
    wire N__59984;
    wire N__59983;
    wire N__59980;
    wire N__59979;
    wire N__59976;
    wire N__59973;
    wire N__59970;
    wire N__59967;
    wire N__59962;
    wire N__59959;
    wire N__59952;
    wire N__59949;
    wire N__59948;
    wire N__59947;
    wire N__59946;
    wire N__59943;
    wire N__59940;
    wire N__59937;
    wire N__59934;
    wire N__59929;
    wire N__59926;
    wire N__59919;
    wire N__59916;
    wire N__59915;
    wire N__59914;
    wire N__59913;
    wire N__59910;
    wire N__59907;
    wire N__59904;
    wire N__59901;
    wire N__59894;
    wire N__59889;
    wire N__59886;
    wire N__59883;
    wire N__59882;
    wire N__59881;
    wire N__59880;
    wire N__59877;
    wire N__59874;
    wire N__59871;
    wire N__59868;
    wire N__59861;
    wire N__59856;
    wire N__59853;
    wire N__59852;
    wire N__59849;
    wire N__59846;
    wire N__59845;
    wire N__59840;
    wire N__59837;
    wire N__59836;
    wire N__59833;
    wire N__59830;
    wire N__59827;
    wire N__59824;
    wire N__59821;
    wire N__59814;
    wire N__59811;
    wire N__59810;
    wire N__59807;
    wire N__59804;
    wire N__59799;
    wire N__59796;
    wire N__59795;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59785;
    wire N__59782;
    wire N__59779;
    wire N__59772;
    wire N__59769;
    wire N__59768;
    wire N__59767;
    wire N__59764;
    wire N__59761;
    wire N__59758;
    wire N__59755;
    wire N__59750;
    wire N__59747;
    wire N__59746;
    wire N__59743;
    wire N__59740;
    wire N__59737;
    wire N__59734;
    wire N__59731;
    wire N__59724;
    wire N__59721;
    wire N__59720;
    wire N__59719;
    wire N__59716;
    wire N__59713;
    wire N__59710;
    wire N__59705;
    wire N__59702;
    wire N__59699;
    wire N__59696;
    wire N__59695;
    wire N__59692;
    wire N__59689;
    wire N__59686;
    wire N__59683;
    wire N__59680;
    wire N__59673;
    wire N__59670;
    wire N__59669;
    wire N__59666;
    wire N__59663;
    wire N__59662;
    wire N__59661;
    wire N__59656;
    wire N__59653;
    wire N__59650;
    wire N__59647;
    wire N__59644;
    wire N__59639;
    wire N__59636;
    wire N__59631;
    wire N__59628;
    wire N__59627;
    wire N__59624;
    wire N__59621;
    wire N__59616;
    wire N__59613;
    wire N__59610;
    wire N__59607;
    wire N__59604;
    wire N__59603;
    wire N__59600;
    wire N__59597;
    wire N__59592;
    wire N__59589;
    wire N__59588;
    wire N__59585;
    wire N__59582;
    wire N__59577;
    wire N__59574;
    wire N__59573;
    wire N__59570;
    wire N__59567;
    wire N__59564;
    wire N__59559;
    wire N__59556;
    wire N__59555;
    wire N__59552;
    wire N__59549;
    wire N__59544;
    wire N__59541;
    wire N__59538;
    wire N__59535;
    wire N__59534;
    wire N__59531;
    wire N__59528;
    wire N__59523;
    wire N__59520;
    wire N__59517;
    wire N__59514;
    wire N__59513;
    wire N__59510;
    wire N__59507;
    wire N__59502;
    wire N__59499;
    wire N__59496;
    wire N__59493;
    wire N__59492;
    wire N__59489;
    wire N__59486;
    wire N__59481;
    wire N__59478;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59468;
    wire N__59467;
    wire N__59464;
    wire N__59459;
    wire N__59454;
    wire N__59451;
    wire N__59448;
    wire N__59447;
    wire N__59446;
    wire N__59443;
    wire N__59440;
    wire N__59439;
    wire N__59436;
    wire N__59433;
    wire N__59428;
    wire N__59423;
    wire N__59420;
    wire N__59419;
    wire N__59416;
    wire N__59413;
    wire N__59410;
    wire N__59407;
    wire N__59404;
    wire N__59397;
    wire N__59394;
    wire N__59393;
    wire N__59390;
    wire N__59387;
    wire N__59386;
    wire N__59383;
    wire N__59380;
    wire N__59377;
    wire N__59374;
    wire N__59367;
    wire N__59366;
    wire N__59363;
    wire N__59362;
    wire N__59359;
    wire N__59356;
    wire N__59353;
    wire N__59352;
    wire N__59349;
    wire N__59348;
    wire N__59347;
    wire N__59346;
    wire N__59343;
    wire N__59340;
    wire N__59337;
    wire N__59334;
    wire N__59327;
    wire N__59316;
    wire N__59315;
    wire N__59312;
    wire N__59309;
    wire N__59308;
    wire N__59307;
    wire N__59302;
    wire N__59299;
    wire N__59296;
    wire N__59293;
    wire N__59288;
    wire N__59283;
    wire N__59280;
    wire N__59277;
    wire N__59276;
    wire N__59273;
    wire N__59270;
    wire N__59267;
    wire N__59264;
    wire N__59259;
    wire N__59256;
    wire N__59253;
    wire N__59250;
    wire N__59247;
    wire N__59244;
    wire N__59241;
    wire N__59238;
    wire N__59235;
    wire N__59232;
    wire N__59229;
    wire N__59228;
    wire N__59225;
    wire N__59224;
    wire N__59221;
    wire N__59220;
    wire N__59217;
    wire N__59214;
    wire N__59211;
    wire N__59208;
    wire N__59203;
    wire N__59198;
    wire N__59195;
    wire N__59192;
    wire N__59189;
    wire N__59184;
    wire N__59181;
    wire N__59178;
    wire N__59177;
    wire N__59174;
    wire N__59171;
    wire N__59168;
    wire N__59165;
    wire N__59160;
    wire N__59157;
    wire N__59154;
    wire N__59151;
    wire N__59150;
    wire N__59147;
    wire N__59144;
    wire N__59141;
    wire N__59138;
    wire N__59137;
    wire N__59134;
    wire N__59131;
    wire N__59128;
    wire N__59121;
    wire N__59118;
    wire N__59115;
    wire N__59112;
    wire N__59109;
    wire N__59108;
    wire N__59105;
    wire N__59102;
    wire N__59099;
    wire N__59096;
    wire N__59091;
    wire N__59090;
    wire N__59087;
    wire N__59084;
    wire N__59081;
    wire N__59076;
    wire N__59075;
    wire N__59070;
    wire N__59067;
    wire N__59064;
    wire N__59061;
    wire N__59058;
    wire N__59057;
    wire N__59056;
    wire N__59053;
    wire N__59048;
    wire N__59043;
    wire N__59042;
    wire N__59039;
    wire N__59036;
    wire N__59033;
    wire N__59030;
    wire N__59025;
    wire N__59022;
    wire N__59021;
    wire N__59018;
    wire N__59015;
    wire N__59012;
    wire N__59009;
    wire N__59006;
    wire N__59001;
    wire N__58998;
    wire N__58995;
    wire N__58992;
    wire N__58989;
    wire N__58986;
    wire N__58983;
    wire N__58980;
    wire N__58977;
    wire N__58974;
    wire N__58971;
    wire N__58968;
    wire N__58965;
    wire N__58962;
    wire N__58959;
    wire N__58958;
    wire N__58957;
    wire N__58956;
    wire N__58955;
    wire N__58950;
    wire N__58945;
    wire N__58942;
    wire N__58939;
    wire N__58936;
    wire N__58929;
    wire N__58928;
    wire N__58923;
    wire N__58922;
    wire N__58921;
    wire N__58920;
    wire N__58917;
    wire N__58914;
    wire N__58911;
    wire N__58908;
    wire N__58905;
    wire N__58902;
    wire N__58893;
    wire N__58890;
    wire N__58887;
    wire N__58884;
    wire N__58883;
    wire N__58882;
    wire N__58875;
    wire N__58872;
    wire N__58871;
    wire N__58868;
    wire N__58865;
    wire N__58862;
    wire N__58857;
    wire N__58854;
    wire N__58851;
    wire N__58848;
    wire N__58847;
    wire N__58842;
    wire N__58839;
    wire N__58836;
    wire N__58833;
    wire N__58830;
    wire N__58827;
    wire N__58824;
    wire N__58821;
    wire N__58820;
    wire N__58817;
    wire N__58814;
    wire N__58811;
    wire N__58806;
    wire N__58803;
    wire N__58800;
    wire N__58797;
    wire N__58794;
    wire N__58793;
    wire N__58790;
    wire N__58789;
    wire N__58786;
    wire N__58783;
    wire N__58782;
    wire N__58779;
    wire N__58776;
    wire N__58773;
    wire N__58770;
    wire N__58767;
    wire N__58758;
    wire N__58755;
    wire N__58752;
    wire N__58749;
    wire N__58746;
    wire N__58743;
    wire N__58740;
    wire N__58737;
    wire N__58734;
    wire N__58733;
    wire N__58730;
    wire N__58727;
    wire N__58726;
    wire N__58721;
    wire N__58718;
    wire N__58713;
    wire N__58710;
    wire N__58709;
    wire N__58706;
    wire N__58703;
    wire N__58700;
    wire N__58697;
    wire N__58694;
    wire N__58689;
    wire N__58688;
    wire N__58685;
    wire N__58682;
    wire N__58681;
    wire N__58680;
    wire N__58679;
    wire N__58678;
    wire N__58675;
    wire N__58672;
    wire N__58669;
    wire N__58666;
    wire N__58663;
    wire N__58660;
    wire N__58653;
    wire N__58650;
    wire N__58647;
    wire N__58644;
    wire N__58641;
    wire N__58638;
    wire N__58629;
    wire N__58626;
    wire N__58623;
    wire N__58620;
    wire N__58617;
    wire N__58614;
    wire N__58611;
    wire N__58608;
    wire N__58605;
    wire N__58602;
    wire N__58601;
    wire N__58598;
    wire N__58595;
    wire N__58592;
    wire N__58587;
    wire N__58584;
    wire N__58583;
    wire N__58580;
    wire N__58577;
    wire N__58572;
    wire N__58569;
    wire N__58566;
    wire N__58563;
    wire N__58560;
    wire N__58559;
    wire N__58556;
    wire N__58555;
    wire N__58554;
    wire N__58551;
    wire N__58548;
    wire N__58543;
    wire N__58536;
    wire N__58533;
    wire N__58530;
    wire N__58529;
    wire N__58526;
    wire N__58525;
    wire N__58524;
    wire N__58521;
    wire N__58518;
    wire N__58513;
    wire N__58506;
    wire N__58503;
    wire N__58500;
    wire N__58499;
    wire N__58498;
    wire N__58497;
    wire N__58494;
    wire N__58487;
    wire N__58482;
    wire N__58479;
    wire N__58478;
    wire N__58475;
    wire N__58472;
    wire N__58469;
    wire N__58466;
    wire N__58461;
    wire N__58458;
    wire N__58457;
    wire N__58454;
    wire N__58451;
    wire N__58448;
    wire N__58445;
    wire N__58440;
    wire N__58439;
    wire N__58438;
    wire N__58437;
    wire N__58436;
    wire N__58433;
    wire N__58432;
    wire N__58431;
    wire N__58430;
    wire N__58429;
    wire N__58428;
    wire N__58427;
    wire N__58426;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58416;
    wire N__58415;
    wire N__58414;
    wire N__58413;
    wire N__58412;
    wire N__58411;
    wire N__58410;
    wire N__58407;
    wire N__58406;
    wire N__58405;
    wire N__58404;
    wire N__58403;
    wire N__58402;
    wire N__58401;
    wire N__58396;
    wire N__58391;
    wire N__58384;
    wire N__58383;
    wire N__58382;
    wire N__58381;
    wire N__58380;
    wire N__58379;
    wire N__58378;
    wire N__58377;
    wire N__58374;
    wire N__58369;
    wire N__58368;
    wire N__58367;
    wire N__58366;
    wire N__58365;
    wire N__58364;
    wire N__58363;
    wire N__58362;
    wire N__58361;
    wire N__58358;
    wire N__58349;
    wire N__58344;
    wire N__58341;
    wire N__58338;
    wire N__58335;
    wire N__58332;
    wire N__58323;
    wire N__58322;
    wire N__58321;
    wire N__58320;
    wire N__58319;
    wire N__58318;
    wire N__58317;
    wire N__58316;
    wire N__58313;
    wire N__58308;
    wire N__58303;
    wire N__58302;
    wire N__58301;
    wire N__58300;
    wire N__58299;
    wire N__58298;
    wire N__58295;
    wire N__58288;
    wire N__58287;
    wire N__58284;
    wire N__58279;
    wire N__58276;
    wire N__58273;
    wire N__58270;
    wire N__58267;
    wire N__58258;
    wire N__58249;
    wire N__58240;
    wire N__58237;
    wire N__58234;
    wire N__58227;
    wire N__58222;
    wire N__58215;
    wire N__58210;
    wire N__58207;
    wire N__58206;
    wire N__58205;
    wire N__58204;
    wire N__58199;
    wire N__58196;
    wire N__58193;
    wire N__58190;
    wire N__58179;
    wire N__58176;
    wire N__58169;
    wire N__58166;
    wire N__58157;
    wire N__58154;
    wire N__58151;
    wire N__58148;
    wire N__58143;
    wire N__58140;
    wire N__58135;
    wire N__58130;
    wire N__58125;
    wire N__58120;
    wire N__58115;
    wire N__58098;
    wire N__58097;
    wire N__58094;
    wire N__58091;
    wire N__58088;
    wire N__58087;
    wire N__58082;
    wire N__58079;
    wire N__58076;
    wire N__58073;
    wire N__58070;
    wire N__58065;
    wire N__58062;
    wire N__58061;
    wire N__58058;
    wire N__58055;
    wire N__58054;
    wire N__58049;
    wire N__58046;
    wire N__58043;
    wire N__58038;
    wire N__58037;
    wire N__58034;
    wire N__58031;
    wire N__58028;
    wire N__58023;
    wire N__58020;
    wire N__58017;
    wire N__58016;
    wire N__58013;
    wire N__58010;
    wire N__58009;
    wire N__58006;
    wire N__58005;
    wire N__58002;
    wire N__57999;
    wire N__57996;
    wire N__57993;
    wire N__57988;
    wire N__57981;
    wire N__57980;
    wire N__57979;
    wire N__57978;
    wire N__57977;
    wire N__57976;
    wire N__57973;
    wire N__57972;
    wire N__57971;
    wire N__57968;
    wire N__57967;
    wire N__57966;
    wire N__57965;
    wire N__57964;
    wire N__57963;
    wire N__57962;
    wire N__57959;
    wire N__57958;
    wire N__57957;
    wire N__57956;
    wire N__57955;
    wire N__57954;
    wire N__57953;
    wire N__57952;
    wire N__57949;
    wire N__57946;
    wire N__57945;
    wire N__57942;
    wire N__57937;
    wire N__57930;
    wire N__57923;
    wire N__57914;
    wire N__57913;
    wire N__57912;
    wire N__57911;
    wire N__57910;
    wire N__57909;
    wire N__57908;
    wire N__57907;
    wire N__57904;
    wire N__57901;
    wire N__57900;
    wire N__57891;
    wire N__57886;
    wire N__57883;
    wire N__57880;
    wire N__57871;
    wire N__57870;
    wire N__57863;
    wire N__57858;
    wire N__57853;
    wire N__57848;
    wire N__57845;
    wire N__57842;
    wire N__57839;
    wire N__57838;
    wire N__57835;
    wire N__57830;
    wire N__57829;
    wire N__57826;
    wire N__57823;
    wire N__57816;
    wire N__57809;
    wire N__57806;
    wire N__57801;
    wire N__57798;
    wire N__57797;
    wire N__57794;
    wire N__57789;
    wire N__57788;
    wire N__57787;
    wire N__57784;
    wire N__57779;
    wire N__57776;
    wire N__57773;
    wire N__57772;
    wire N__57771;
    wire N__57768;
    wire N__57765;
    wire N__57762;
    wire N__57759;
    wire N__57756;
    wire N__57751;
    wire N__57748;
    wire N__57743;
    wire N__57736;
    wire N__57723;
    wire N__57722;
    wire N__57719;
    wire N__57718;
    wire N__57715;
    wire N__57710;
    wire N__57705;
    wire N__57702;
    wire N__57699;
    wire N__57696;
    wire N__57695;
    wire N__57692;
    wire N__57689;
    wire N__57684;
    wire N__57681;
    wire N__57678;
    wire N__57675;
    wire N__57672;
    wire N__57669;
    wire N__57668;
    wire N__57667;
    wire N__57664;
    wire N__57661;
    wire N__57658;
    wire N__57653;
    wire N__57648;
    wire N__57645;
    wire N__57642;
    wire N__57641;
    wire N__57640;
    wire N__57639;
    wire N__57636;
    wire N__57633;
    wire N__57630;
    wire N__57627;
    wire N__57624;
    wire N__57621;
    wire N__57618;
    wire N__57615;
    wire N__57612;
    wire N__57607;
    wire N__57600;
    wire N__57599;
    wire N__57596;
    wire N__57593;
    wire N__57588;
    wire N__57587;
    wire N__57584;
    wire N__57581;
    wire N__57576;
    wire N__57573;
    wire N__57570;
    wire N__57567;
    wire N__57566;
    wire N__57563;
    wire N__57560;
    wire N__57557;
    wire N__57552;
    wire N__57549;
    wire N__57546;
    wire N__57543;
    wire N__57540;
    wire N__57537;
    wire N__57534;
    wire N__57531;
    wire N__57528;
    wire N__57527;
    wire N__57524;
    wire N__57521;
    wire N__57516;
    wire N__57515;
    wire N__57510;
    wire N__57507;
    wire N__57506;
    wire N__57503;
    wire N__57500;
    wire N__57495;
    wire N__57492;
    wire N__57491;
    wire N__57490;
    wire N__57483;
    wire N__57480;
    wire N__57477;
    wire N__57476;
    wire N__57473;
    wire N__57470;
    wire N__57465;
    wire N__57462;
    wire N__57459;
    wire N__57458;
    wire N__57453;
    wire N__57450;
    wire N__57447;
    wire N__57444;
    wire N__57441;
    wire N__57438;
    wire N__57435;
    wire N__57432;
    wire N__57429;
    wire N__57426;
    wire N__57423;
    wire N__57420;
    wire N__57419;
    wire N__57416;
    wire N__57413;
    wire N__57408;
    wire N__57407;
    wire N__57402;
    wire N__57399;
    wire N__57396;
    wire N__57393;
    wire N__57392;
    wire N__57389;
    wire N__57388;
    wire N__57385;
    wire N__57382;
    wire N__57379;
    wire N__57376;
    wire N__57373;
    wire N__57366;
    wire N__57363;
    wire N__57360;
    wire N__57357;
    wire N__57356;
    wire N__57355;
    wire N__57352;
    wire N__57347;
    wire N__57344;
    wire N__57339;
    wire N__57336;
    wire N__57333;
    wire N__57330;
    wire N__57327;
    wire N__57324;
    wire N__57321;
    wire N__57318;
    wire N__57317;
    wire N__57316;
    wire N__57313;
    wire N__57310;
    wire N__57307;
    wire N__57300;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57285;
    wire N__57282;
    wire N__57279;
    wire N__57276;
    wire N__57273;
    wire N__57270;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57258;
    wire N__57255;
    wire N__57252;
    wire N__57249;
    wire N__57246;
    wire N__57243;
    wire N__57240;
    wire N__57237;
    wire N__57234;
    wire N__57231;
    wire N__57228;
    wire N__57225;
    wire N__57222;
    wire N__57219;
    wire N__57216;
    wire N__57213;
    wire N__57210;
    wire N__57207;
    wire N__57204;
    wire N__57201;
    wire N__57198;
    wire N__57195;
    wire N__57192;
    wire N__57189;
    wire N__57186;
    wire N__57183;
    wire N__57180;
    wire N__57177;
    wire N__57174;
    wire N__57171;
    wire N__57168;
    wire N__57165;
    wire N__57162;
    wire N__57161;
    wire N__57158;
    wire N__57155;
    wire N__57154;
    wire N__57151;
    wire N__57146;
    wire N__57143;
    wire N__57138;
    wire N__57135;
    wire N__57132;
    wire N__57129;
    wire N__57128;
    wire N__57127;
    wire N__57124;
    wire N__57121;
    wire N__57118;
    wire N__57115;
    wire N__57108;
    wire N__57105;
    wire N__57102;
    wire N__57099;
    wire N__57096;
    wire N__57095;
    wire N__57094;
    wire N__57091;
    wire N__57088;
    wire N__57085;
    wire N__57082;
    wire N__57075;
    wire N__57072;
    wire N__57069;
    wire N__57066;
    wire N__57065;
    wire N__57062;
    wire N__57059;
    wire N__57054;
    wire N__57053;
    wire N__57050;
    wire N__57047;
    wire N__57042;
    wire N__57039;
    wire N__57038;
    wire N__57037;
    wire N__57036;
    wire N__57033;
    wire N__57030;
    wire N__57027;
    wire N__57024;
    wire N__57023;
    wire N__57020;
    wire N__57015;
    wire N__57010;
    wire N__57003;
    wire N__57002;
    wire N__57001;
    wire N__57000;
    wire N__56999;
    wire N__56998;
    wire N__56995;
    wire N__56992;
    wire N__56989;
    wire N__56986;
    wire N__56983;
    wire N__56980;
    wire N__56975;
    wire N__56966;
    wire N__56961;
    wire N__56958;
    wire N__56955;
    wire N__56952;
    wire N__56949;
    wire N__56946;
    wire N__56943;
    wire N__56940;
    wire N__56937;
    wire N__56934;
    wire N__56931;
    wire N__56928;
    wire N__56925;
    wire N__56922;
    wire N__56919;
    wire N__56916;
    wire N__56913;
    wire N__56912;
    wire N__56909;
    wire N__56906;
    wire N__56903;
    wire N__56900;
    wire N__56895;
    wire N__56892;
    wire N__56891;
    wire N__56888;
    wire N__56885;
    wire N__56880;
    wire N__56879;
    wire N__56876;
    wire N__56873;
    wire N__56868;
    wire N__56865;
    wire N__56864;
    wire N__56863;
    wire N__56860;
    wire N__56857;
    wire N__56854;
    wire N__56851;
    wire N__56844;
    wire N__56841;
    wire N__56840;
    wire N__56839;
    wire N__56836;
    wire N__56833;
    wire N__56830;
    wire N__56823;
    wire N__56820;
    wire N__56819;
    wire N__56818;
    wire N__56815;
    wire N__56812;
    wire N__56809;
    wire N__56802;
    wire N__56799;
    wire N__56798;
    wire N__56797;
    wire N__56794;
    wire N__56791;
    wire N__56788;
    wire N__56781;
    wire N__56778;
    wire N__56777;
    wire N__56774;
    wire N__56771;
    wire N__56770;
    wire N__56765;
    wire N__56762;
    wire N__56757;
    wire N__56754;
    wire N__56753;
    wire N__56750;
    wire N__56747;
    wire N__56746;
    wire N__56741;
    wire N__56738;
    wire N__56733;
    wire N__56730;
    wire N__56729;
    wire N__56728;
    wire N__56725;
    wire N__56722;
    wire N__56721;
    wire N__56718;
    wire N__56717;
    wire N__56714;
    wire N__56711;
    wire N__56708;
    wire N__56705;
    wire N__56702;
    wire N__56695;
    wire N__56688;
    wire N__56687;
    wire N__56684;
    wire N__56681;
    wire N__56678;
    wire N__56673;
    wire N__56670;
    wire N__56667;
    wire N__56664;
    wire N__56661;
    wire N__56658;
    wire N__56655;
    wire N__56652;
    wire N__56649;
    wire N__56646;
    wire N__56643;
    wire N__56640;
    wire N__56637;
    wire N__56634;
    wire N__56631;
    wire N__56628;
    wire N__56625;
    wire N__56624;
    wire N__56619;
    wire N__56616;
    wire N__56613;
    wire N__56610;
    wire N__56609;
    wire N__56608;
    wire N__56605;
    wire N__56600;
    wire N__56597;
    wire N__56594;
    wire N__56591;
    wire N__56586;
    wire N__56585;
    wire N__56580;
    wire N__56577;
    wire N__56574;
    wire N__56571;
    wire N__56568;
    wire N__56567;
    wire N__56564;
    wire N__56561;
    wire N__56560;
    wire N__56555;
    wire N__56552;
    wire N__56549;
    wire N__56546;
    wire N__56541;
    wire N__56538;
    wire N__56535;
    wire N__56532;
    wire N__56529;
    wire N__56526;
    wire N__56523;
    wire N__56520;
    wire N__56517;
    wire N__56516;
    wire N__56513;
    wire N__56510;
    wire N__56505;
    wire N__56502;
    wire N__56499;
    wire N__56496;
    wire N__56493;
    wire N__56492;
    wire N__56489;
    wire N__56488;
    wire N__56485;
    wire N__56482;
    wire N__56481;
    wire N__56478;
    wire N__56475;
    wire N__56472;
    wire N__56467;
    wire N__56460;
    wire N__56457;
    wire N__56456;
    wire N__56455;
    wire N__56454;
    wire N__56451;
    wire N__56448;
    wire N__56443;
    wire N__56438;
    wire N__56435;
    wire N__56432;
    wire N__56427;
    wire N__56424;
    wire N__56421;
    wire N__56418;
    wire N__56415;
    wire N__56414;
    wire N__56411;
    wire N__56408;
    wire N__56405;
    wire N__56402;
    wire N__56397;
    wire N__56394;
    wire N__56391;
    wire N__56390;
    wire N__56385;
    wire N__56382;
    wire N__56381;
    wire N__56376;
    wire N__56373;
    wire N__56372;
    wire N__56369;
    wire N__56368;
    wire N__56365;
    wire N__56362;
    wire N__56359;
    wire N__56352;
    wire N__56351;
    wire N__56350;
    wire N__56345;
    wire N__56342;
    wire N__56339;
    wire N__56334;
    wire N__56331;
    wire N__56330;
    wire N__56329;
    wire N__56324;
    wire N__56321;
    wire N__56318;
    wire N__56315;
    wire N__56310;
    wire N__56307;
    wire N__56304;
    wire N__56301;
    wire N__56300;
    wire N__56297;
    wire N__56292;
    wire N__56291;
    wire N__56290;
    wire N__56287;
    wire N__56282;
    wire N__56277;
    wire N__56274;
    wire N__56273;
    wire N__56272;
    wire N__56269;
    wire N__56264;
    wire N__56259;
    wire N__56256;
    wire N__56253;
    wire N__56250;
    wire N__56249;
    wire N__56248;
    wire N__56245;
    wire N__56242;
    wire N__56239;
    wire N__56236;
    wire N__56229;
    wire N__56228;
    wire N__56227;
    wire N__56224;
    wire N__56221;
    wire N__56220;
    wire N__56217;
    wire N__56214;
    wire N__56209;
    wire N__56206;
    wire N__56199;
    wire N__56196;
    wire N__56193;
    wire N__56192;
    wire N__56189;
    wire N__56186;
    wire N__56181;
    wire N__56178;
    wire N__56177;
    wire N__56174;
    wire N__56171;
    wire N__56166;
    wire N__56165;
    wire N__56162;
    wire N__56159;
    wire N__56156;
    wire N__56151;
    wire N__56148;
    wire N__56145;
    wire N__56142;
    wire N__56139;
    wire N__56136;
    wire N__56135;
    wire N__56130;
    wire N__56127;
    wire N__56124;
    wire N__56121;
    wire N__56118;
    wire N__56115;
    wire N__56114;
    wire N__56113;
    wire N__56110;
    wire N__56105;
    wire N__56100;
    wire N__56097;
    wire N__56094;
    wire N__56091;
    wire N__56088;
    wire N__56087;
    wire N__56084;
    wire N__56081;
    wire N__56076;
    wire N__56075;
    wire N__56072;
    wire N__56069;
    wire N__56068;
    wire N__56063;
    wire N__56060;
    wire N__56059;
    wire N__56056;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56040;
    wire N__56037;
    wire N__56034;
    wire N__56031;
    wire N__56028;
    wire N__56027;
    wire N__56022;
    wire N__56021;
    wire N__56018;
    wire N__56015;
    wire N__56012;
    wire N__56007;
    wire N__56004;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55992;
    wire N__55991;
    wire N__55988;
    wire N__55987;
    wire N__55986;
    wire N__55983;
    wire N__55980;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55968;
    wire N__55963;
    wire N__55956;
    wire N__55953;
    wire N__55950;
    wire N__55947;
    wire N__55944;
    wire N__55941;
    wire N__55938;
    wire N__55935;
    wire N__55934;
    wire N__55933;
    wire N__55932;
    wire N__55931;
    wire N__55930;
    wire N__55929;
    wire N__55928;
    wire N__55927;
    wire N__55926;
    wire N__55923;
    wire N__55920;
    wire N__55917;
    wire N__55916;
    wire N__55913;
    wire N__55908;
    wire N__55905;
    wire N__55902;
    wire N__55899;
    wire N__55898;
    wire N__55895;
    wire N__55892;
    wire N__55887;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55869;
    wire N__55866;
    wire N__55863;
    wire N__55860;
    wire N__55855;
    wire N__55852;
    wire N__55849;
    wire N__55846;
    wire N__55841;
    wire N__55838;
    wire N__55835;
    wire N__55830;
    wire N__55827;
    wire N__55824;
    wire N__55819;
    wire N__55814;
    wire N__55811;
    wire N__55806;
    wire N__55803;
    wire N__55802;
    wire N__55801;
    wire N__55800;
    wire N__55795;
    wire N__55792;
    wire N__55789;
    wire N__55782;
    wire N__55779;
    wire N__55776;
    wire N__55775;
    wire N__55774;
    wire N__55771;
    wire N__55768;
    wire N__55765;
    wire N__55762;
    wire N__55759;
    wire N__55756;
    wire N__55753;
    wire N__55750;
    wire N__55743;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55733;
    wire N__55730;
    wire N__55729;
    wire N__55728;
    wire N__55725;
    wire N__55722;
    wire N__55719;
    wire N__55716;
    wire N__55709;
    wire N__55706;
    wire N__55703;
    wire N__55698;
    wire N__55695;
    wire N__55692;
    wire N__55691;
    wire N__55688;
    wire N__55687;
    wire N__55684;
    wire N__55681;
    wire N__55676;
    wire N__55673;
    wire N__55670;
    wire N__55665;
    wire N__55662;
    wire N__55659;
    wire N__55656;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55646;
    wire N__55643;
    wire N__55640;
    wire N__55635;
    wire N__55632;
    wire N__55629;
    wire N__55626;
    wire N__55625;
    wire N__55624;
    wire N__55623;
    wire N__55620;
    wire N__55617;
    wire N__55614;
    wire N__55613;
    wire N__55610;
    wire N__55607;
    wire N__55606;
    wire N__55603;
    wire N__55600;
    wire N__55597;
    wire N__55592;
    wire N__55589;
    wire N__55584;
    wire N__55581;
    wire N__55578;
    wire N__55571;
    wire N__55566;
    wire N__55563;
    wire N__55562;
    wire N__55559;
    wire N__55558;
    wire N__55557;
    wire N__55554;
    wire N__55551;
    wire N__55550;
    wire N__55549;
    wire N__55548;
    wire N__55545;
    wire N__55542;
    wire N__55539;
    wire N__55536;
    wire N__55533;
    wire N__55530;
    wire N__55527;
    wire N__55520;
    wire N__55517;
    wire N__55506;
    wire N__55503;
    wire N__55500;
    wire N__55497;
    wire N__55494;
    wire N__55491;
    wire N__55490;
    wire N__55489;
    wire N__55486;
    wire N__55481;
    wire N__55476;
    wire N__55473;
    wire N__55470;
    wire N__55467;
    wire N__55464;
    wire N__55461;
    wire N__55458;
    wire N__55455;
    wire N__55452;
    wire N__55449;
    wire N__55448;
    wire N__55447;
    wire N__55446;
    wire N__55443;
    wire N__55440;
    wire N__55437;
    wire N__55436;
    wire N__55435;
    wire N__55432;
    wire N__55429;
    wire N__55424;
    wire N__55421;
    wire N__55418;
    wire N__55407;
    wire N__55404;
    wire N__55401;
    wire N__55400;
    wire N__55399;
    wire N__55398;
    wire N__55395;
    wire N__55390;
    wire N__55387;
    wire N__55382;
    wire N__55379;
    wire N__55376;
    wire N__55371;
    wire N__55370;
    wire N__55367;
    wire N__55364;
    wire N__55361;
    wire N__55358;
    wire N__55353;
    wire N__55350;
    wire N__55347;
    wire N__55344;
    wire N__55341;
    wire N__55338;
    wire N__55335;
    wire N__55332;
    wire N__55329;
    wire N__55326;
    wire N__55325;
    wire N__55322;
    wire N__55319;
    wire N__55314;
    wire N__55313;
    wire N__55308;
    wire N__55305;
    wire N__55302;
    wire N__55299;
    wire N__55296;
    wire N__55293;
    wire N__55290;
    wire N__55289;
    wire N__55284;
    wire N__55281;
    wire N__55278;
    wire N__55275;
    wire N__55272;
    wire N__55269;
    wire N__55266;
    wire N__55263;
    wire N__55260;
    wire N__55257;
    wire N__55254;
    wire N__55251;
    wire N__55248;
    wire N__55245;
    wire N__55242;
    wire N__55239;
    wire N__55236;
    wire N__55235;
    wire N__55232;
    wire N__55231;
    wire N__55228;
    wire N__55225;
    wire N__55222;
    wire N__55219;
    wire N__55216;
    wire N__55213;
    wire N__55210;
    wire N__55207;
    wire N__55204;
    wire N__55197;
    wire N__55196;
    wire N__55191;
    wire N__55188;
    wire N__55187;
    wire N__55182;
    wire N__55179;
    wire N__55176;
    wire N__55173;
    wire N__55170;
    wire N__55167;
    wire N__55164;
    wire N__55163;
    wire N__55158;
    wire N__55155;
    wire N__55152;
    wire N__55149;
    wire N__55146;
    wire N__55143;
    wire N__55140;
    wire N__55139;
    wire N__55136;
    wire N__55133;
    wire N__55130;
    wire N__55127;
    wire N__55124;
    wire N__55119;
    wire N__55118;
    wire N__55115;
    wire N__55112;
    wire N__55109;
    wire N__55104;
    wire N__55103;
    wire N__55100;
    wire N__55097;
    wire N__55092;
    wire N__55091;
    wire N__55088;
    wire N__55085;
    wire N__55080;
    wire N__55079;
    wire N__55076;
    wire N__55073;
    wire N__55068;
    wire N__55065;
    wire N__55064;
    wire N__55063;
    wire N__55056;
    wire N__55053;
    wire N__55050;
    wire N__55049;
    wire N__55046;
    wire N__55043;
    wire N__55040;
    wire N__55037;
    wire N__55034;
    wire N__55029;
    wire N__55026;
    wire N__55023;
    wire N__55020;
    wire N__55017;
    wire N__55014;
    wire N__55011;
    wire N__55008;
    wire N__55007;
    wire N__55004;
    wire N__55001;
    wire N__54998;
    wire N__54993;
    wire N__54990;
    wire N__54987;
    wire N__54984;
    wire N__54981;
    wire N__54980;
    wire N__54977;
    wire N__54974;
    wire N__54973;
    wire N__54968;
    wire N__54965;
    wire N__54960;
    wire N__54957;
    wire N__54956;
    wire N__54953;
    wire N__54950;
    wire N__54949;
    wire N__54944;
    wire N__54941;
    wire N__54936;
    wire N__54933;
    wire N__54932;
    wire N__54931;
    wire N__54928;
    wire N__54925;
    wire N__54922;
    wire N__54917;
    wire N__54914;
    wire N__54909;
    wire N__54906;
    wire N__54905;
    wire N__54902;
    wire N__54899;
    wire N__54898;
    wire N__54893;
    wire N__54890;
    wire N__54885;
    wire N__54882;
    wire N__54881;
    wire N__54878;
    wire N__54875;
    wire N__54874;
    wire N__54869;
    wire N__54866;
    wire N__54861;
    wire N__54858;
    wire N__54857;
    wire N__54854;
    wire N__54851;
    wire N__54850;
    wire N__54845;
    wire N__54842;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54834;
    wire N__54833;
    wire N__54832;
    wire N__54831;
    wire N__54830;
    wire N__54829;
    wire N__54828;
    wire N__54827;
    wire N__54826;
    wire N__54825;
    wire N__54824;
    wire N__54823;
    wire N__54822;
    wire N__54821;
    wire N__54818;
    wire N__54815;
    wire N__54812;
    wire N__54809;
    wire N__54806;
    wire N__54803;
    wire N__54800;
    wire N__54797;
    wire N__54794;
    wire N__54791;
    wire N__54788;
    wire N__54785;
    wire N__54782;
    wire N__54779;
    wire N__54776;
    wire N__54773;
    wire N__54770;
    wire N__54769;
    wire N__54762;
    wire N__54753;
    wire N__54744;
    wire N__54735;
    wire N__54730;
    wire N__54727;
    wire N__54714;
    wire N__54711;
    wire N__54708;
    wire N__54705;
    wire N__54702;
    wire N__54699;
    wire N__54698;
    wire N__54697;
    wire N__54696;
    wire N__54695;
    wire N__54694;
    wire N__54691;
    wire N__54688;
    wire N__54685;
    wire N__54682;
    wire N__54679;
    wire N__54676;
    wire N__54671;
    wire N__54662;
    wire N__54657;
    wire N__54656;
    wire N__54655;
    wire N__54654;
    wire N__54653;
    wire N__54652;
    wire N__54651;
    wire N__54650;
    wire N__54649;
    wire N__54648;
    wire N__54645;
    wire N__54642;
    wire N__54639;
    wire N__54636;
    wire N__54633;
    wire N__54630;
    wire N__54627;
    wire N__54624;
    wire N__54621;
    wire N__54618;
    wire N__54611;
    wire N__54602;
    wire N__54597;
    wire N__54594;
    wire N__54585;
    wire N__54582;
    wire N__54579;
    wire N__54576;
    wire N__54575;
    wire N__54574;
    wire N__54571;
    wire N__54568;
    wire N__54565;
    wire N__54560;
    wire N__54557;
    wire N__54552;
    wire N__54549;
    wire N__54546;
    wire N__54543;
    wire N__54542;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54532;
    wire N__54527;
    wire N__54524;
    wire N__54519;
    wire N__54516;
    wire N__54513;
    wire N__54510;
    wire N__54509;
    wire N__54508;
    wire N__54505;
    wire N__54502;
    wire N__54499;
    wire N__54494;
    wire N__54491;
    wire N__54486;
    wire N__54483;
    wire N__54482;
    wire N__54479;
    wire N__54476;
    wire N__54475;
    wire N__54470;
    wire N__54467;
    wire N__54462;
    wire N__54459;
    wire N__54458;
    wire N__54455;
    wire N__54452;
    wire N__54451;
    wire N__54446;
    wire N__54443;
    wire N__54438;
    wire N__54435;
    wire N__54432;
    wire N__54429;
    wire N__54428;
    wire N__54425;
    wire N__54422;
    wire N__54421;
    wire N__54416;
    wire N__54413;
    wire N__54408;
    wire N__54405;
    wire N__54402;
    wire N__54399;
    wire N__54398;
    wire N__54395;
    wire N__54392;
    wire N__54391;
    wire N__54386;
    wire N__54383;
    wire N__54378;
    wire N__54375;
    wire N__54374;
    wire N__54371;
    wire N__54368;
    wire N__54363;
    wire N__54362;
    wire N__54359;
    wire N__54356;
    wire N__54351;
    wire N__54348;
    wire N__54347;
    wire N__54346;
    wire N__54343;
    wire N__54340;
    wire N__54337;
    wire N__54332;
    wire N__54329;
    wire N__54324;
    wire N__54321;
    wire N__54320;
    wire N__54317;
    wire N__54314;
    wire N__54313;
    wire N__54308;
    wire N__54305;
    wire N__54300;
    wire N__54297;
    wire N__54296;
    wire N__54295;
    wire N__54292;
    wire N__54289;
    wire N__54286;
    wire N__54281;
    wire N__54278;
    wire N__54273;
    wire N__54270;
    wire N__54269;
    wire N__54266;
    wire N__54263;
    wire N__54262;
    wire N__54257;
    wire N__54254;
    wire N__54249;
    wire N__54246;
    wire N__54245;
    wire N__54242;
    wire N__54239;
    wire N__54238;
    wire N__54233;
    wire N__54230;
    wire N__54225;
    wire N__54222;
    wire N__54221;
    wire N__54218;
    wire N__54215;
    wire N__54214;
    wire N__54209;
    wire N__54206;
    wire N__54201;
    wire N__54200;
    wire N__54199;
    wire N__54198;
    wire N__54197;
    wire N__54196;
    wire N__54193;
    wire N__54190;
    wire N__54187;
    wire N__54184;
    wire N__54181;
    wire N__54178;
    wire N__54173;
    wire N__54164;
    wire N__54159;
    wire N__54156;
    wire N__54155;
    wire N__54152;
    wire N__54149;
    wire N__54148;
    wire N__54143;
    wire N__54140;
    wire N__54135;
    wire N__54132;
    wire N__54131;
    wire N__54128;
    wire N__54125;
    wire N__54120;
    wire N__54119;
    wire N__54116;
    wire N__54113;
    wire N__54108;
    wire N__54105;
    wire N__54102;
    wire N__54099;
    wire N__54098;
    wire N__54095;
    wire N__54092;
    wire N__54089;
    wire N__54084;
    wire N__54081;
    wire N__54080;
    wire N__54077;
    wire N__54074;
    wire N__54073;
    wire N__54070;
    wire N__54067;
    wire N__54064;
    wire N__54057;
    wire N__54054;
    wire N__54051;
    wire N__54048;
    wire N__54045;
    wire N__54044;
    wire N__54043;
    wire N__54040;
    wire N__54037;
    wire N__54034;
    wire N__54027;
    wire N__54024;
    wire N__54021;
    wire N__54018;
    wire N__54015;
    wire N__54012;
    wire N__54011;
    wire N__54010;
    wire N__54009;
    wire N__54006;
    wire N__54005;
    wire N__54002;
    wire N__53999;
    wire N__53998;
    wire N__53995;
    wire N__53994;
    wire N__53991;
    wire N__53988;
    wire N__53983;
    wire N__53976;
    wire N__53967;
    wire N__53966;
    wire N__53963;
    wire N__53960;
    wire N__53957;
    wire N__53952;
    wire N__53949;
    wire N__53946;
    wire N__53943;
    wire N__53942;
    wire N__53941;
    wire N__53938;
    wire N__53935;
    wire N__53932;
    wire N__53929;
    wire N__53926;
    wire N__53923;
    wire N__53916;
    wire N__53913;
    wire N__53910;
    wire N__53907;
    wire N__53906;
    wire N__53905;
    wire N__53904;
    wire N__53901;
    wire N__53900;
    wire N__53897;
    wire N__53896;
    wire N__53893;
    wire N__53892;
    wire N__53891;
    wire N__53888;
    wire N__53883;
    wire N__53872;
    wire N__53865;
    wire N__53862;
    wire N__53859;
    wire N__53856;
    wire N__53853;
    wire N__53850;
    wire N__53847;
    wire N__53846;
    wire N__53843;
    wire N__53840;
    wire N__53835;
    wire N__53832;
    wire N__53829;
    wire N__53826;
    wire N__53825;
    wire N__53820;
    wire N__53817;
    wire N__53814;
    wire N__53813;
    wire N__53812;
    wire N__53809;
    wire N__53804;
    wire N__53803;
    wire N__53798;
    wire N__53795;
    wire N__53792;
    wire N__53787;
    wire N__53784;
    wire N__53783;
    wire N__53782;
    wire N__53779;
    wire N__53774;
    wire N__53769;
    wire N__53766;
    wire N__53765;
    wire N__53764;
    wire N__53763;
    wire N__53758;
    wire N__53755;
    wire N__53752;
    wire N__53749;
    wire N__53744;
    wire N__53739;
    wire N__53738;
    wire N__53733;
    wire N__53730;
    wire N__53727;
    wire N__53726;
    wire N__53723;
    wire N__53720;
    wire N__53715;
    wire N__53714;
    wire N__53711;
    wire N__53710;
    wire N__53707;
    wire N__53706;
    wire N__53703;
    wire N__53700;
    wire N__53697;
    wire N__53694;
    wire N__53691;
    wire N__53688;
    wire N__53679;
    wire N__53678;
    wire N__53677;
    wire N__53674;
    wire N__53671;
    wire N__53668;
    wire N__53665;
    wire N__53658;
    wire N__53655;
    wire N__53652;
    wire N__53649;
    wire N__53646;
    wire N__53643;
    wire N__53640;
    wire N__53637;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53625;
    wire N__53622;
    wire N__53621;
    wire N__53618;
    wire N__53615;
    wire N__53612;
    wire N__53607;
    wire N__53606;
    wire N__53605;
    wire N__53602;
    wire N__53599;
    wire N__53596;
    wire N__53595;
    wire N__53594;
    wire N__53591;
    wire N__53588;
    wire N__53585;
    wire N__53580;
    wire N__53577;
    wire N__53568;
    wire N__53565;
    wire N__53562;
    wire N__53561;
    wire N__53558;
    wire N__53555;
    wire N__53550;
    wire N__53549;
    wire N__53548;
    wire N__53545;
    wire N__53542;
    wire N__53539;
    wire N__53536;
    wire N__53535;
    wire N__53532;
    wire N__53527;
    wire N__53524;
    wire N__53519;
    wire N__53514;
    wire N__53511;
    wire N__53510;
    wire N__53507;
    wire N__53504;
    wire N__53503;
    wire N__53498;
    wire N__53495;
    wire N__53494;
    wire N__53489;
    wire N__53486;
    wire N__53483;
    wire N__53480;
    wire N__53475;
    wire N__53472;
    wire N__53471;
    wire N__53470;
    wire N__53467;
    wire N__53462;
    wire N__53459;
    wire N__53456;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53446;
    wire N__53439;
    wire N__53436;
    wire N__53433;
    wire N__53432;
    wire N__53431;
    wire N__53430;
    wire N__53427;
    wire N__53424;
    wire N__53419;
    wire N__53416;
    wire N__53413;
    wire N__53406;
    wire N__53405;
    wire N__53404;
    wire N__53401;
    wire N__53396;
    wire N__53393;
    wire N__53388;
    wire N__53385;
    wire N__53382;
    wire N__53379;
    wire N__53376;
    wire N__53373;
    wire N__53370;
    wire N__53367;
    wire N__53364;
    wire N__53363;
    wire N__53362;
    wire N__53361;
    wire N__53360;
    wire N__53355;
    wire N__53352;
    wire N__53349;
    wire N__53346;
    wire N__53343;
    wire N__53340;
    wire N__53337;
    wire N__53334;
    wire N__53331;
    wire N__53328;
    wire N__53319;
    wire N__53318;
    wire N__53315;
    wire N__53312;
    wire N__53311;
    wire N__53308;
    wire N__53303;
    wire N__53300;
    wire N__53295;
    wire N__53292;
    wire N__53289;
    wire N__53286;
    wire N__53283;
    wire N__53280;
    wire N__53277;
    wire N__53274;
    wire N__53273;
    wire N__53268;
    wire N__53265;
    wire N__53262;
    wire N__53259;
    wire N__53256;
    wire N__53253;
    wire N__53250;
    wire N__53247;
    wire N__53244;
    wire N__53241;
    wire N__53238;
    wire N__53237;
    wire N__53234;
    wire N__53231;
    wire N__53226;
    wire N__53225;
    wire N__53222;
    wire N__53221;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53211;
    wire N__53208;
    wire N__53207;
    wire N__53204;
    wire N__53201;
    wire N__53198;
    wire N__53195;
    wire N__53192;
    wire N__53189;
    wire N__53178;
    wire N__53175;
    wire N__53174;
    wire N__53171;
    wire N__53168;
    wire N__53165;
    wire N__53162;
    wire N__53159;
    wire N__53154;
    wire N__53153;
    wire N__53150;
    wire N__53147;
    wire N__53142;
    wire N__53139;
    wire N__53136;
    wire N__53133;
    wire N__53130;
    wire N__53129;
    wire N__53126;
    wire N__53125;
    wire N__53122;
    wire N__53121;
    wire N__53118;
    wire N__53115;
    wire N__53110;
    wire N__53103;
    wire N__53100;
    wire N__53099;
    wire N__53098;
    wire N__53097;
    wire N__53096;
    wire N__53093;
    wire N__53088;
    wire N__53085;
    wire N__53082;
    wire N__53077;
    wire N__53070;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53054;
    wire N__53051;
    wire N__53048;
    wire N__53045;
    wire N__53044;
    wire N__53039;
    wire N__53036;
    wire N__53031;
    wire N__53028;
    wire N__53027;
    wire N__53024;
    wire N__53023;
    wire N__53022;
    wire N__53021;
    wire N__53018;
    wire N__53017;
    wire N__53014;
    wire N__53011;
    wire N__53006;
    wire N__53001;
    wire N__52992;
    wire N__52989;
    wire N__52988;
    wire N__52985;
    wire N__52982;
    wire N__52977;
    wire N__52976;
    wire N__52973;
    wire N__52970;
    wire N__52967;
    wire N__52964;
    wire N__52961;
    wire N__52956;
    wire N__52955;
    wire N__52952;
    wire N__52949;
    wire N__52948;
    wire N__52947;
    wire N__52944;
    wire N__52937;
    wire N__52932;
    wire N__52929;
    wire N__52926;
    wire N__52923;
    wire N__52920;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52910;
    wire N__52907;
    wire N__52904;
    wire N__52901;
    wire N__52898;
    wire N__52895;
    wire N__52890;
    wire N__52887;
    wire N__52884;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52876;
    wire N__52873;
    wire N__52870;
    wire N__52863;
    wire N__52860;
    wire N__52859;
    wire N__52856;
    wire N__52853;
    wire N__52850;
    wire N__52845;
    wire N__52842;
    wire N__52841;
    wire N__52836;
    wire N__52833;
    wire N__52832;
    wire N__52831;
    wire N__52830;
    wire N__52827;
    wire N__52824;
    wire N__52823;
    wire N__52818;
    wire N__52815;
    wire N__52812;
    wire N__52809;
    wire N__52806;
    wire N__52805;
    wire N__52802;
    wire N__52799;
    wire N__52796;
    wire N__52793;
    wire N__52790;
    wire N__52779;
    wire N__52776;
    wire N__52773;
    wire N__52772;
    wire N__52769;
    wire N__52766;
    wire N__52761;
    wire N__52758;
    wire N__52757;
    wire N__52756;
    wire N__52753;
    wire N__52750;
    wire N__52747;
    wire N__52744;
    wire N__52743;
    wire N__52740;
    wire N__52737;
    wire N__52734;
    wire N__52731;
    wire N__52722;
    wire N__52721;
    wire N__52718;
    wire N__52715;
    wire N__52712;
    wire N__52707;
    wire N__52706;
    wire N__52705;
    wire N__52698;
    wire N__52695;
    wire N__52692;
    wire N__52689;
    wire N__52686;
    wire N__52683;
    wire N__52682;
    wire N__52681;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52653;
    wire N__52652;
    wire N__52651;
    wire N__52648;
    wire N__52645;
    wire N__52642;
    wire N__52637;
    wire N__52634;
    wire N__52631;
    wire N__52626;
    wire N__52623;
    wire N__52622;
    wire N__52621;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52605;
    wire N__52604;
    wire N__52601;
    wire N__52598;
    wire N__52595;
    wire N__52592;
    wire N__52589;
    wire N__52586;
    wire N__52581;
    wire N__52578;
    wire N__52575;
    wire N__52572;
    wire N__52569;
    wire N__52566;
    wire N__52563;
    wire N__52560;
    wire N__52557;
    wire N__52554;
    wire N__52551;
    wire N__52548;
    wire N__52545;
    wire N__52544;
    wire N__52543;
    wire N__52542;
    wire N__52539;
    wire N__52532;
    wire N__52529;
    wire N__52524;
    wire N__52523;
    wire N__52520;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52510;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52500;
    wire N__52497;
    wire N__52494;
    wire N__52489;
    wire N__52482;
    wire N__52481;
    wire N__52478;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52453;
    wire N__52448;
    wire N__52443;
    wire N__52440;
    wire N__52437;
    wire N__52434;
    wire N__52433;
    wire N__52430;
    wire N__52427;
    wire N__52426;
    wire N__52421;
    wire N__52418;
    wire N__52415;
    wire N__52410;
    wire N__52407;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52397;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52389;
    wire N__52386;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52355;
    wire N__52354;
    wire N__52351;
    wire N__52350;
    wire N__52349;
    wire N__52346;
    wire N__52343;
    wire N__52340;
    wire N__52335;
    wire N__52332;
    wire N__52329;
    wire N__52324;
    wire N__52321;
    wire N__52314;
    wire N__52311;
    wire N__52310;
    wire N__52305;
    wire N__52302;
    wire N__52299;
    wire N__52296;
    wire N__52295;
    wire N__52292;
    wire N__52291;
    wire N__52288;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52276;
    wire N__52269;
    wire N__52268;
    wire N__52265;
    wire N__52262;
    wire N__52261;
    wire N__52260;
    wire N__52259;
    wire N__52256;
    wire N__52253;
    wire N__52250;
    wire N__52245;
    wire N__52236;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52221;
    wire N__52218;
    wire N__52215;
    wire N__52214;
    wire N__52211;
    wire N__52208;
    wire N__52203;
    wire N__52200;
    wire N__52199;
    wire N__52196;
    wire N__52193;
    wire N__52192;
    wire N__52187;
    wire N__52184;
    wire N__52181;
    wire N__52178;
    wire N__52175;
    wire N__52170;
    wire N__52167;
    wire N__52166;
    wire N__52163;
    wire N__52162;
    wire N__52159;
    wire N__52158;
    wire N__52155;
    wire N__52154;
    wire N__52153;
    wire N__52150;
    wire N__52149;
    wire N__52144;
    wire N__52141;
    wire N__52136;
    wire N__52131;
    wire N__52122;
    wire N__52121;
    wire N__52120;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52107;
    wire N__52106;
    wire N__52105;
    wire N__52104;
    wire N__52103;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52088;
    wire N__52079;
    wire N__52072;
    wire N__52065;
    wire N__52064;
    wire N__52063;
    wire N__52062;
    wire N__52061;
    wire N__52060;
    wire N__52059;
    wire N__52056;
    wire N__52053;
    wire N__52052;
    wire N__52049;
    wire N__52044;
    wire N__52039;
    wire N__52036;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52022;
    wire N__52011;
    wire N__52008;
    wire N__52005;
    wire N__52002;
    wire N__51999;
    wire N__51996;
    wire N__51995;
    wire N__51992;
    wire N__51989;
    wire N__51984;
    wire N__51983;
    wire N__51978;
    wire N__51975;
    wire N__51974;
    wire N__51969;
    wire N__51966;
    wire N__51965;
    wire N__51960;
    wire N__51957;
    wire N__51954;
    wire N__51953;
    wire N__51950;
    wire N__51947;
    wire N__51942;
    wire N__51939;
    wire N__51938;
    wire N__51935;
    wire N__51932;
    wire N__51931;
    wire N__51926;
    wire N__51923;
    wire N__51920;
    wire N__51917;
    wire N__51914;
    wire N__51911;
    wire N__51906;
    wire N__51905;
    wire N__51902;
    wire N__51901;
    wire N__51900;
    wire N__51899;
    wire N__51898;
    wire N__51897;
    wire N__51894;
    wire N__51889;
    wire N__51886;
    wire N__51881;
    wire N__51878;
    wire N__51873;
    wire N__51864;
    wire N__51861;
    wire N__51860;
    wire N__51859;
    wire N__51858;
    wire N__51857;
    wire N__51856;
    wire N__51855;
    wire N__51852;
    wire N__51851;
    wire N__51850;
    wire N__51847;
    wire N__51842;
    wire N__51839;
    wire N__51838;
    wire N__51837;
    wire N__51836;
    wire N__51831;
    wire N__51828;
    wire N__51825;
    wire N__51822;
    wire N__51821;
    wire N__51814;
    wire N__51811;
    wire N__51806;
    wire N__51801;
    wire N__51796;
    wire N__51793;
    wire N__51790;
    wire N__51787;
    wire N__51782;
    wire N__51777;
    wire N__51774;
    wire N__51769;
    wire N__51766;
    wire N__51759;
    wire N__51758;
    wire N__51753;
    wire N__51750;
    wire N__51749;
    wire N__51748;
    wire N__51747;
    wire N__51746;
    wire N__51745;
    wire N__51742;
    wire N__51737;
    wire N__51734;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51720;
    wire N__51711;
    wire N__51708;
    wire N__51707;
    wire N__51704;
    wire N__51701;
    wire N__51698;
    wire N__51697;
    wire N__51696;
    wire N__51695;
    wire N__51694;
    wire N__51693;
    wire N__51690;
    wire N__51687;
    wire N__51686;
    wire N__51685;
    wire N__51684;
    wire N__51679;
    wire N__51676;
    wire N__51673;
    wire N__51670;
    wire N__51665;
    wire N__51662;
    wire N__51657;
    wire N__51654;
    wire N__51651;
    wire N__51646;
    wire N__51643;
    wire N__51632;
    wire N__51627;
    wire N__51624;
    wire N__51623;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51591;
    wire N__51590;
    wire N__51587;
    wire N__51586;
    wire N__51583;
    wire N__51580;
    wire N__51575;
    wire N__51572;
    wire N__51569;
    wire N__51564;
    wire N__51561;
    wire N__51560;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51552;
    wire N__51551;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51541;
    wire N__51538;
    wire N__51533;
    wire N__51522;
    wire N__51521;
    wire N__51520;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51510;
    wire N__51509;
    wire N__51506;
    wire N__51503;
    wire N__51500;
    wire N__51495;
    wire N__51492;
    wire N__51483;
    wire N__51480;
    wire N__51479;
    wire N__51474;
    wire N__51471;
    wire N__51468;
    wire N__51465;
    wire N__51464;
    wire N__51459;
    wire N__51456;
    wire N__51453;
    wire N__51450;
    wire N__51447;
    wire N__51444;
    wire N__51441;
    wire N__51438;
    wire N__51437;
    wire N__51434;
    wire N__51431;
    wire N__51428;
    wire N__51425;
    wire N__51420;
    wire N__51417;
    wire N__51414;
    wire N__51411;
    wire N__51408;
    wire N__51405;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51393;
    wire N__51390;
    wire N__51387;
    wire N__51384;
    wire N__51381;
    wire N__51378;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51370;
    wire N__51367;
    wire N__51364;
    wire N__51361;
    wire N__51358;
    wire N__51355;
    wire N__51348;
    wire N__51347;
    wire N__51344;
    wire N__51341;
    wire N__51340;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51326;
    wire N__51321;
    wire N__51318;
    wire N__51317;
    wire N__51314;
    wire N__51311;
    wire N__51306;
    wire N__51305;
    wire N__51302;
    wire N__51299;
    wire N__51294;
    wire N__51291;
    wire N__51288;
    wire N__51287;
    wire N__51284;
    wire N__51281;
    wire N__51276;
    wire N__51275;
    wire N__51272;
    wire N__51269;
    wire N__51264;
    wire N__51261;
    wire N__51258;
    wire N__51255;
    wire N__51252;
    wire N__51249;
    wire N__51248;
    wire N__51245;
    wire N__51242;
    wire N__51239;
    wire N__51234;
    wire N__51231;
    wire N__51230;
    wire N__51227;
    wire N__51224;
    wire N__51221;
    wire N__51218;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51192;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51180;
    wire N__51177;
    wire N__51176;
    wire N__51173;
    wire N__51170;
    wire N__51165;
    wire N__51164;
    wire N__51161;
    wire N__51158;
    wire N__51153;
    wire N__51150;
    wire N__51149;
    wire N__51146;
    wire N__51143;
    wire N__51138;
    wire N__51137;
    wire N__51134;
    wire N__51131;
    wire N__51126;
    wire N__51123;
    wire N__51122;
    wire N__51119;
    wire N__51116;
    wire N__51111;
    wire N__51110;
    wire N__51107;
    wire N__51104;
    wire N__51099;
    wire N__51096;
    wire N__51095;
    wire N__51092;
    wire N__51089;
    wire N__51088;
    wire N__51083;
    wire N__51080;
    wire N__51077;
    wire N__51074;
    wire N__51069;
    wire N__51066;
    wire N__51065;
    wire N__51062;
    wire N__51059;
    wire N__51054;
    wire N__51053;
    wire N__51050;
    wire N__51047;
    wire N__51042;
    wire N__51039;
    wire N__51038;
    wire N__51035;
    wire N__51032;
    wire N__51027;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51015;
    wire N__51012;
    wire N__51011;
    wire N__51008;
    wire N__51005;
    wire N__51000;
    wire N__50999;
    wire N__50996;
    wire N__50993;
    wire N__50988;
    wire N__50985;
    wire N__50982;
    wire N__50979;
    wire N__50976;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50964;
    wire N__50961;
    wire N__50958;
    wire N__50955;
    wire N__50952;
    wire N__50949;
    wire N__50946;
    wire N__50945;
    wire N__50942;
    wire N__50939;
    wire N__50934;
    wire N__50933;
    wire N__50930;
    wire N__50927;
    wire N__50922;
    wire N__50919;
    wire N__50918;
    wire N__50915;
    wire N__50912;
    wire N__50907;
    wire N__50906;
    wire N__50903;
    wire N__50900;
    wire N__50895;
    wire N__50892;
    wire N__50891;
    wire N__50888;
    wire N__50885;
    wire N__50880;
    wire N__50879;
    wire N__50876;
    wire N__50873;
    wire N__50868;
    wire N__50865;
    wire N__50864;
    wire N__50861;
    wire N__50858;
    wire N__50853;
    wire N__50852;
    wire N__50849;
    wire N__50846;
    wire N__50841;
    wire N__50838;
    wire N__50835;
    wire N__50832;
    wire N__50831;
    wire N__50828;
    wire N__50825;
    wire N__50820;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50812;
    wire N__50809;
    wire N__50804;
    wire N__50799;
    wire N__50796;
    wire N__50795;
    wire N__50792;
    wire N__50789;
    wire N__50786;
    wire N__50781;
    wire N__50778;
    wire N__50775;
    wire N__50772;
    wire N__50769;
    wire N__50766;
    wire N__50763;
    wire N__50760;
    wire N__50757;
    wire N__50754;
    wire N__50751;
    wire N__50748;
    wire N__50745;
    wire N__50742;
    wire N__50739;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50718;
    wire N__50715;
    wire N__50714;
    wire N__50711;
    wire N__50708;
    wire N__50707;
    wire N__50704;
    wire N__50701;
    wire N__50698;
    wire N__50691;
    wire N__50688;
    wire N__50685;
    wire N__50682;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50665;
    wire N__50662;
    wire N__50659;
    wire N__50656;
    wire N__50649;
    wire N__50646;
    wire N__50645;
    wire N__50642;
    wire N__50639;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50622;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50612;
    wire N__50609;
    wire N__50608;
    wire N__50605;
    wire N__50602;
    wire N__50599;
    wire N__50598;
    wire N__50595;
    wire N__50590;
    wire N__50587;
    wire N__50580;
    wire N__50579;
    wire N__50578;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50556;
    wire N__50553;
    wire N__50544;
    wire N__50541;
    wire N__50540;
    wire N__50537;
    wire N__50534;
    wire N__50529;
    wire N__50526;
    wire N__50523;
    wire N__50522;
    wire N__50521;
    wire N__50518;
    wire N__50515;
    wire N__50512;
    wire N__50511;
    wire N__50506;
    wire N__50503;
    wire N__50500;
    wire N__50497;
    wire N__50492;
    wire N__50487;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50478;
    wire N__50473;
    wire N__50470;
    wire N__50469;
    wire N__50462;
    wire N__50459;
    wire N__50454;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50442;
    wire N__50439;
    wire N__50438;
    wire N__50435;
    wire N__50434;
    wire N__50431;
    wire N__50430;
    wire N__50421;
    wire N__50418;
    wire N__50417;
    wire N__50414;
    wire N__50411;
    wire N__50408;
    wire N__50405;
    wire N__50402;
    wire N__50399;
    wire N__50394;
    wire N__50393;
    wire N__50390;
    wire N__50389;
    wire N__50388;
    wire N__50385;
    wire N__50380;
    wire N__50377;
    wire N__50376;
    wire N__50375;
    wire N__50372;
    wire N__50369;
    wire N__50366;
    wire N__50361;
    wire N__50358;
    wire N__50355;
    wire N__50350;
    wire N__50343;
    wire N__50342;
    wire N__50339;
    wire N__50338;
    wire N__50337;
    wire N__50334;
    wire N__50331;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50313;
    wire N__50310;
    wire N__50307;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50297;
    wire N__50294;
    wire N__50291;
    wire N__50288;
    wire N__50283;
    wire N__50280;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50268;
    wire N__50265;
    wire N__50262;
    wire N__50259;
    wire N__50256;
    wire N__50253;
    wire N__50252;
    wire N__50251;
    wire N__50250;
    wire N__50247;
    wire N__50242;
    wire N__50239;
    wire N__50234;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50217;
    wire N__50216;
    wire N__50213;
    wire N__50210;
    wire N__50207;
    wire N__50204;
    wire N__50199;
    wire N__50198;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50190;
    wire N__50187;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50173;
    wire N__50166;
    wire N__50163;
    wire N__50160;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50139;
    wire N__50138;
    wire N__50137;
    wire N__50134;
    wire N__50129;
    wire N__50128;
    wire N__50127;
    wire N__50126;
    wire N__50121;
    wire N__50118;
    wire N__50115;
    wire N__50112;
    wire N__50109;
    wire N__50104;
    wire N__50097;
    wire N__50096;
    wire N__50091;
    wire N__50088;
    wire N__50085;
    wire N__50082;
    wire N__50081;
    wire N__50080;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50068;
    wire N__50063;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50048;
    wire N__50045;
    wire N__50042;
    wire N__50037;
    wire N__50036;
    wire N__50033;
    wire N__50032;
    wire N__50029;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50015;
    wire N__50012;
    wire N__50011;
    wire N__50006;
    wire N__50003;
    wire N__50000;
    wire N__49995;
    wire N__49992;
    wire N__49989;
    wire N__49986;
    wire N__49983;
    wire N__49980;
    wire N__49977;
    wire N__49976;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49959;
    wire N__49958;
    wire N__49955;
    wire N__49952;
    wire N__49949;
    wire N__49944;
    wire N__49941;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49933;
    wire N__49930;
    wire N__49927;
    wire N__49924;
    wire N__49921;
    wire N__49916;
    wire N__49911;
    wire N__49910;
    wire N__49907;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49895;
    wire N__49894;
    wire N__49887;
    wire N__49884;
    wire N__49883;
    wire N__49880;
    wire N__49879;
    wire N__49876;
    wire N__49873;
    wire N__49870;
    wire N__49867;
    wire N__49860;
    wire N__49859;
    wire N__49858;
    wire N__49855;
    wire N__49852;
    wire N__49849;
    wire N__49846;
    wire N__49843;
    wire N__49840;
    wire N__49835;
    wire N__49830;
    wire N__49827;
    wire N__49824;
    wire N__49823;
    wire N__49820;
    wire N__49817;
    wire N__49816;
    wire N__49813;
    wire N__49808;
    wire N__49805;
    wire N__49802;
    wire N__49797;
    wire N__49794;
    wire N__49793;
    wire N__49790;
    wire N__49787;
    wire N__49782;
    wire N__49781;
    wire N__49778;
    wire N__49775;
    wire N__49772;
    wire N__49769;
    wire N__49766;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49754;
    wire N__49751;
    wire N__49748;
    wire N__49743;
    wire N__49740;
    wire N__49739;
    wire N__49736;
    wire N__49733;
    wire N__49732;
    wire N__49729;
    wire N__49724;
    wire N__49719;
    wire N__49716;
    wire N__49713;
    wire N__49712;
    wire N__49711;
    wire N__49708;
    wire N__49705;
    wire N__49702;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49688;
    wire N__49687;
    wire N__49686;
    wire N__49683;
    wire N__49682;
    wire N__49679;
    wire N__49676;
    wire N__49673;
    wire N__49670;
    wire N__49667;
    wire N__49656;
    wire N__49655;
    wire N__49652;
    wire N__49649;
    wire N__49648;
    wire N__49647;
    wire N__49644;
    wire N__49641;
    wire N__49638;
    wire N__49635;
    wire N__49628;
    wire N__49625;
    wire N__49620;
    wire N__49617;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49609;
    wire N__49606;
    wire N__49601;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49587;
    wire N__49584;
    wire N__49581;
    wire N__49580;
    wire N__49577;
    wire N__49574;
    wire N__49569;
    wire N__49568;
    wire N__49565;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49548;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49538;
    wire N__49535;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49519;
    wire N__49514;
    wire N__49511;
    wire N__49508;
    wire N__49505;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49495;
    wire N__49490;
    wire N__49485;
    wire N__49484;
    wire N__49481;
    wire N__49478;
    wire N__49475;
    wire N__49472;
    wire N__49467;
    wire N__49464;
    wire N__49463;
    wire N__49460;
    wire N__49457;
    wire N__49452;
    wire N__49449;
    wire N__49446;
    wire N__49443;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49430;
    wire N__49429;
    wire N__49428;
    wire N__49425;
    wire N__49424;
    wire N__49421;
    wire N__49418;
    wire N__49415;
    wire N__49406;
    wire N__49403;
    wire N__49400;
    wire N__49395;
    wire N__49386;
    wire N__49383;
    wire N__49380;
    wire N__49379;
    wire N__49376;
    wire N__49373;
    wire N__49370;
    wire N__49365;
    wire N__49364;
    wire N__49361;
    wire N__49358;
    wire N__49353;
    wire N__49350;
    wire N__49347;
    wire N__49344;
    wire N__49341;
    wire N__49338;
    wire N__49335;
    wire N__49332;
    wire N__49329;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49310;
    wire N__49309;
    wire N__49306;
    wire N__49303;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49287;
    wire N__49284;
    wire N__49281;
    wire N__49278;
    wire N__49277;
    wire N__49276;
    wire N__49275;
    wire N__49274;
    wire N__49273;
    wire N__49272;
    wire N__49271;
    wire N__49270;
    wire N__49269;
    wire N__49268;
    wire N__49265;
    wire N__49264;
    wire N__49263;
    wire N__49262;
    wire N__49255;
    wire N__49250;
    wire N__49247;
    wire N__49238;
    wire N__49237;
    wire N__49236;
    wire N__49233;
    wire N__49228;
    wire N__49225;
    wire N__49216;
    wire N__49211;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49195;
    wire N__49190;
    wire N__49185;
    wire N__49184;
    wire N__49181;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49173;
    wire N__49168;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49160;
    wire N__49157;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49136;
    wire N__49125;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49117;
    wire N__49116;
    wire N__49115;
    wire N__49112;
    wire N__49111;
    wire N__49108;
    wire N__49105;
    wire N__49096;
    wire N__49095;
    wire N__49094;
    wire N__49093;
    wire N__49092;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49082;
    wire N__49079;
    wire N__49074;
    wire N__49073;
    wire N__49072;
    wire N__49071;
    wire N__49070;
    wire N__49067;
    wire N__49064;
    wire N__49061;
    wire N__49056;
    wire N__49051;
    wire N__49050;
    wire N__49047;
    wire N__49040;
    wire N__49035;
    wire N__49028;
    wire N__49025;
    wire N__49020;
    wire N__49015;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48978;
    wire N__48975;
    wire N__48974;
    wire N__48973;
    wire N__48966;
    wire N__48965;
    wire N__48962;
    wire N__48959;
    wire N__48958;
    wire N__48953;
    wire N__48950;
    wire N__48947;
    wire N__48944;
    wire N__48941;
    wire N__48936;
    wire N__48933;
    wire N__48930;
    wire N__48927;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48917;
    wire N__48914;
    wire N__48911;
    wire N__48906;
    wire N__48905;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48897;
    wire N__48894;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48874;
    wire N__48869;
    wire N__48866;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48850;
    wire N__48849;
    wire N__48846;
    wire N__48845;
    wire N__48842;
    wire N__48839;
    wire N__48838;
    wire N__48835;
    wire N__48834;
    wire N__48829;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48815;
    wire N__48810;
    wire N__48801;
    wire N__48800;
    wire N__48797;
    wire N__48796;
    wire N__48793;
    wire N__48788;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48771;
    wire N__48768;
    wire N__48765;
    wire N__48762;
    wire N__48759;
    wire N__48756;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48746;
    wire N__48743;
    wire N__48738;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48726;
    wire N__48723;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48713;
    wire N__48708;
    wire N__48707;
    wire N__48704;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48681;
    wire N__48680;
    wire N__48677;
    wire N__48674;
    wire N__48669;
    wire N__48666;
    wire N__48663;
    wire N__48662;
    wire N__48661;
    wire N__48660;
    wire N__48657;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48636;
    wire N__48633;
    wire N__48630;
    wire N__48627;
    wire N__48624;
    wire N__48621;
    wire N__48618;
    wire N__48615;
    wire N__48612;
    wire N__48609;
    wire N__48608;
    wire N__48603;
    wire N__48600;
    wire N__48599;
    wire N__48596;
    wire N__48593;
    wire N__48592;
    wire N__48591;
    wire N__48586;
    wire N__48581;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48561;
    wire N__48558;
    wire N__48557;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48543;
    wire N__48540;
    wire N__48539;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48531;
    wire N__48528;
    wire N__48525;
    wire N__48522;
    wire N__48519;
    wire N__48516;
    wire N__48509;
    wire N__48508;
    wire N__48507;
    wire N__48502;
    wire N__48497;
    wire N__48492;
    wire N__48491;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48473;
    wire N__48470;
    wire N__48467;
    wire N__48462;
    wire N__48459;
    wire N__48454;
    wire N__48447;
    wire N__48444;
    wire N__48443;
    wire N__48440;
    wire N__48437;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48408;
    wire N__48405;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48395;
    wire N__48392;
    wire N__48389;
    wire N__48386;
    wire N__48383;
    wire N__48380;
    wire N__48377;
    wire N__48372;
    wire N__48369;
    wire N__48366;
    wire N__48363;
    wire N__48360;
    wire N__48359;
    wire N__48358;
    wire N__48355;
    wire N__48350;
    wire N__48345;
    wire N__48344;
    wire N__48341;
    wire N__48338;
    wire N__48335;
    wire N__48332;
    wire N__48329;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48312;
    wire N__48309;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48299;
    wire N__48294;
    wire N__48293;
    wire N__48290;
    wire N__48289;
    wire N__48284;
    wire N__48283;
    wire N__48282;
    wire N__48281;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48267;
    wire N__48264;
    wire N__48261;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48240;
    wire N__48239;
    wire N__48238;
    wire N__48235;
    wire N__48228;
    wire N__48225;
    wire N__48222;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48212;
    wire N__48207;
    wire N__48204;
    wire N__48201;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48191;
    wire N__48190;
    wire N__48187;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48169;
    wire N__48164;
    wire N__48161;
    wire N__48158;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48128;
    wire N__48127;
    wire N__48126;
    wire N__48125;
    wire N__48124;
    wire N__48123;
    wire N__48120;
    wire N__48117;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48084;
    wire N__48075;
    wire N__48070;
    wire N__48063;
    wire N__48060;
    wire N__48059;
    wire N__48058;
    wire N__48057;
    wire N__48056;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48032;
    wire N__48023;
    wire N__48018;
    wire N__48015;
    wire N__48014;
    wire N__48013;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__47999;
    wire N__47996;
    wire N__47991;
    wire N__47990;
    wire N__47989;
    wire N__47986;
    wire N__47983;
    wire N__47980;
    wire N__47975;
    wire N__47972;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47952;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47940;
    wire N__47937;
    wire N__47936;
    wire N__47933;
    wire N__47932;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47916;
    wire N__47913;
    wire N__47910;
    wire N__47907;
    wire N__47906;
    wire N__47903;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47891;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47840;
    wire N__47837;
    wire N__47834;
    wire N__47829;
    wire N__47826;
    wire N__47825;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47815;
    wire N__47808;
    wire N__47805;
    wire N__47804;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47794;
    wire N__47791;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47768;
    wire N__47767;
    wire N__47764;
    wire N__47761;
    wire N__47758;
    wire N__47751;
    wire N__47748;
    wire N__47747;
    wire N__47746;
    wire N__47743;
    wire N__47740;
    wire N__47737;
    wire N__47730;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47684;
    wire N__47683;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47646;
    wire N__47645;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47630;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47613;
    wire N__47610;
    wire N__47609;
    wire N__47606;
    wire N__47603;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47589;
    wire N__47586;
    wire N__47583;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47552;
    wire N__47547;
    wire N__47544;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47536;
    wire N__47533;
    wire N__47532;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47478;
    wire N__47475;
    wire N__47474;
    wire N__47471;
    wire N__47468;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47436;
    wire N__47433;
    wire N__47432;
    wire N__47427;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47417;
    wire N__47412;
    wire N__47409;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47378;
    wire N__47375;
    wire N__47374;
    wire N__47369;
    wire N__47366;
    wire N__47361;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47264;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47237;
    wire N__47234;
    wire N__47233;
    wire N__47230;
    wire N__47225;
    wire N__47220;
    wire N__47219;
    wire N__47216;
    wire N__47213;
    wire N__47208;
    wire N__47207;
    wire N__47204;
    wire N__47201;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47168;
    wire N__47165;
    wire N__47164;
    wire N__47161;
    wire N__47158;
    wire N__47155;
    wire N__47152;
    wire N__47145;
    wire N__47142;
    wire N__47141;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47117;
    wire N__47114;
    wire N__47111;
    wire N__47106;
    wire N__47103;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47082;
    wire N__47079;
    wire N__47078;
    wire N__47073;
    wire N__47070;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47037;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47025;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47003;
    wire N__46998;
    wire N__46995;
    wire N__46994;
    wire N__46991;
    wire N__46990;
    wire N__46987;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46975;
    wire N__46968;
    wire N__46967;
    wire N__46964;
    wire N__46961;
    wire N__46958;
    wire N__46955;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46941;
    wire N__46940;
    wire N__46937;
    wire N__46936;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46919;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46897;
    wire N__46892;
    wire N__46889;
    wire N__46886;
    wire N__46875;
    wire N__46872;
    wire N__46869;
    wire N__46868;
    wire N__46865;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46839;
    wire N__46836;
    wire N__46835;
    wire N__46832;
    wire N__46829;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46809;
    wire N__46804;
    wire N__46801;
    wire N__46794;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46786;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46765;
    wire N__46758;
    wire N__46755;
    wire N__46752;
    wire N__46749;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46743;
    wire N__46742;
    wire N__46741;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46726;
    wire N__46721;
    wire N__46720;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46706;
    wire N__46703;
    wire N__46698;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46667;
    wire N__46666;
    wire N__46665;
    wire N__46662;
    wire N__46659;
    wire N__46654;
    wire N__46647;
    wire N__46646;
    wire N__46645;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46626;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46618;
    wire N__46615;
    wire N__46612;
    wire N__46609;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46595;
    wire N__46592;
    wire N__46589;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46569;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46557;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46530;
    wire N__46529;
    wire N__46528;
    wire N__46525;
    wire N__46524;
    wire N__46521;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46491;
    wire N__46490;
    wire N__46487;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46445;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46424;
    wire N__46423;
    wire N__46420;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46404;
    wire N__46401;
    wire N__46392;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46328;
    wire N__46327;
    wire N__46324;
    wire N__46323;
    wire N__46320;
    wire N__46313;
    wire N__46308;
    wire N__46307;
    wire N__46304;
    wire N__46301;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46293;
    wire N__46290;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46269;
    wire N__46266;
    wire N__46265;
    wire N__46262;
    wire N__46259;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46205;
    wire N__46204;
    wire N__46203;
    wire N__46202;
    wire N__46201;
    wire N__46200;
    wire N__46199;
    wire N__46198;
    wire N__46197;
    wire N__46196;
    wire N__46195;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46188;
    wire N__46187;
    wire N__46186;
    wire N__46185;
    wire N__46184;
    wire N__46183;
    wire N__46182;
    wire N__46181;
    wire N__46170;
    wire N__46163;
    wire N__46154;
    wire N__46149;
    wire N__46148;
    wire N__46145;
    wire N__46142;
    wire N__46129;
    wire N__46124;
    wire N__46119;
    wire N__46116;
    wire N__46109;
    wire N__46106;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46073;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46058;
    wire N__46055;
    wire N__46054;
    wire N__46053;
    wire N__46050;
    wire N__46049;
    wire N__46048;
    wire N__46047;
    wire N__46046;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46038;
    wire N__46033;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46028;
    wire N__46027;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46019;
    wire N__46016;
    wire N__46005;
    wire N__45998;
    wire N__45995;
    wire N__45992;
    wire N__45991;
    wire N__45988;
    wire N__45987;
    wire N__45986;
    wire N__45985;
    wire N__45982;
    wire N__45975;
    wire N__45966;
    wire N__45963;
    wire N__45958;
    wire N__45955;
    wire N__45944;
    wire N__45941;
    wire N__45938;
    wire N__45933;
    wire N__45926;
    wire N__45915;
    wire N__45912;
    wire N__45911;
    wire N__45910;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45906;
    wire N__45905;
    wire N__45904;
    wire N__45903;
    wire N__45902;
    wire N__45901;
    wire N__45900;
    wire N__45899;
    wire N__45898;
    wire N__45897;
    wire N__45896;
    wire N__45895;
    wire N__45894;
    wire N__45887;
    wire N__45874;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45862;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45837;
    wire N__45836;
    wire N__45835;
    wire N__45834;
    wire N__45833;
    wire N__45826;
    wire N__45823;
    wire N__45820;
    wire N__45815;
    wire N__45810;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45796;
    wire N__45791;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45758;
    wire N__45757;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45738;
    wire N__45737;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45720;
    wire N__45719;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45681;
    wire N__45680;
    wire N__45679;
    wire N__45676;
    wire N__45673;
    wire N__45670;
    wire N__45663;
    wire N__45660;
    wire N__45659;
    wire N__45658;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45633;
    wire N__45632;
    wire N__45631;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45612;
    wire N__45611;
    wire N__45608;
    wire N__45605;
    wire N__45602;
    wire N__45601;
    wire N__45596;
    wire N__45593;
    wire N__45588;
    wire N__45587;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45558;
    wire N__45557;
    wire N__45556;
    wire N__45555;
    wire N__45554;
    wire N__45553;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45521;
    wire N__45516;
    wire N__45513;
    wire N__45512;
    wire N__45503;
    wire N__45494;
    wire N__45491;
    wire N__45486;
    wire N__45477;
    wire N__45474;
    wire N__45473;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45453;
    wire N__45452;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45432;
    wire N__45431;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45411;
    wire N__45408;
    wire N__45407;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45387;
    wire N__45386;
    wire N__45385;
    wire N__45382;
    wire N__45379;
    wire N__45376;
    wire N__45373;
    wire N__45366;
    wire N__45365;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45345;
    wire N__45342;
    wire N__45341;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45283;
    wire N__45278;
    wire N__45275;
    wire N__45270;
    wire N__45267;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45259;
    wire N__45254;
    wire N__45251;
    wire N__45246;
    wire N__45243;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45235;
    wire N__45230;
    wire N__45227;
    wire N__45222;
    wire N__45221;
    wire N__45220;
    wire N__45219;
    wire N__45218;
    wire N__45217;
    wire N__45216;
    wire N__45215;
    wire N__45214;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45210;
    wire N__45209;
    wire N__45208;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45152;
    wire N__45145;
    wire N__45136;
    wire N__45127;
    wire N__45122;
    wire N__45121;
    wire N__45116;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45083;
    wire N__45082;
    wire N__45079;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45041;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45026;
    wire N__45023;
    wire N__45018;
    wire N__45015;
    wire N__45014;
    wire N__45011;
    wire N__45008;
    wire N__45007;
    wire N__45002;
    wire N__44999;
    wire N__44994;
    wire N__44991;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44983;
    wire N__44978;
    wire N__44975;
    wire N__44970;
    wire N__44967;
    wire N__44966;
    wire N__44963;
    wire N__44960;
    wire N__44959;
    wire N__44954;
    wire N__44951;
    wire N__44946;
    wire N__44943;
    wire N__44942;
    wire N__44939;
    wire N__44936;
    wire N__44935;
    wire N__44930;
    wire N__44927;
    wire N__44922;
    wire N__44919;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44907;
    wire N__44906;
    wire N__44903;
    wire N__44900;
    wire N__44895;
    wire N__44892;
    wire N__44891;
    wire N__44888;
    wire N__44885;
    wire N__44884;
    wire N__44879;
    wire N__44876;
    wire N__44871;
    wire N__44868;
    wire N__44867;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44852;
    wire N__44849;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44828;
    wire N__44827;
    wire N__44826;
    wire N__44825;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44801;
    wire N__44792;
    wire N__44787;
    wire N__44784;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44776;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44762;
    wire N__44757;
    wire N__44754;
    wire N__44753;
    wire N__44750;
    wire N__44747;
    wire N__44742;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44730;
    wire N__44727;
    wire N__44726;
    wire N__44723;
    wire N__44720;
    wire N__44719;
    wire N__44714;
    wire N__44711;
    wire N__44706;
    wire N__44703;
    wire N__44702;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44687;
    wire N__44684;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44648;
    wire N__44647;
    wire N__44646;
    wire N__44645;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44621;
    wire N__44612;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44597;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44589;
    wire N__44586;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44547;
    wire N__44544;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44518;
    wire N__44511;
    wire N__44508;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44498;
    wire N__44497;
    wire N__44496;
    wire N__44493;
    wire N__44486;
    wire N__44481;
    wire N__44478;
    wire N__44477;
    wire N__44476;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44464;
    wire N__44457;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44449;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44346;
    wire N__44345;
    wire N__44344;
    wire N__44339;
    wire N__44336;
    wire N__44335;
    wire N__44332;
    wire N__44327;
    wire N__44324;
    wire N__44319;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44296;
    wire N__44293;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44270;
    wire N__44269;
    wire N__44264;
    wire N__44261;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44238;
    wire N__44237;
    wire N__44234;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44186;
    wire N__44181;
    wire N__44180;
    wire N__44177;
    wire N__44174;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44157;
    wire N__44154;
    wire N__44153;
    wire N__44150;
    wire N__44147;
    wire N__44142;
    wire N__44141;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44131;
    wire N__44128;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44112;
    wire N__44111;
    wire N__44110;
    wire N__44107;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44060;
    wire N__44057;
    wire N__44054;
    wire N__44049;
    wire N__44048;
    wire N__44047;
    wire N__44040;
    wire N__44037;
    wire N__44036;
    wire N__44033;
    wire N__44030;
    wire N__44027;
    wire N__44024;
    wire N__44019;
    wire N__44016;
    wire N__44015;
    wire N__44012;
    wire N__44011;
    wire N__44008;
    wire N__44005;
    wire N__44002;
    wire N__43999;
    wire N__43992;
    wire N__43989;
    wire N__43988;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43976;
    wire N__43971;
    wire N__43970;
    wire N__43969;
    wire N__43966;
    wire N__43961;
    wire N__43958;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43934;
    wire N__43931;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43915;
    wire N__43912;
    wire N__43905;
    wire N__43902;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43892;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43877;
    wire N__43876;
    wire N__43873;
    wire N__43868;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43847;
    wire N__43846;
    wire N__43845;
    wire N__43838;
    wire N__43837;
    wire N__43836;
    wire N__43833;
    wire N__43832;
    wire N__43831;
    wire N__43830;
    wire N__43827;
    wire N__43822;
    wire N__43819;
    wire N__43814;
    wire N__43811;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43792;
    wire N__43789;
    wire N__43782;
    wire N__43779;
    wire N__43778;
    wire N__43777;
    wire N__43776;
    wire N__43773;
    wire N__43766;
    wire N__43761;
    wire N__43758;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43721;
    wire N__43720;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43712;
    wire N__43709;
    wire N__43706;
    wire N__43703;
    wire N__43696;
    wire N__43689;
    wire N__43686;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43676;
    wire N__43675;
    wire N__43668;
    wire N__43665;
    wire N__43664;
    wire N__43661;
    wire N__43658;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43646;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43626;
    wire N__43625;
    wire N__43624;
    wire N__43621;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43595;
    wire N__43594;
    wire N__43593;
    wire N__43592;
    wire N__43591;
    wire N__43590;
    wire N__43589;
    wire N__43588;
    wire N__43587;
    wire N__43586;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43544;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43528;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43500;
    wire N__43499;
    wire N__43498;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43479;
    wire N__43478;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43458;
    wire N__43455;
    wire N__43454;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43427;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43407;
    wire N__43406;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43386;
    wire N__43383;
    wire N__43382;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43352;
    wire N__43351;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43339;
    wire N__43334;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43316;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43298;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43283;
    wire N__43282;
    wire N__43281;
    wire N__43280;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43256;
    wire N__43247;
    wire N__43242;
    wire N__43239;
    wire N__43238;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43228;
    wire N__43225;
    wire N__43218;
    wire N__43215;
    wire N__43214;
    wire N__43211;
    wire N__43208;
    wire N__43207;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43191;
    wire N__43190;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43173;
    wire N__43172;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43152;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43131;
    wire N__43130;
    wire N__43129;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43113;
    wire N__43112;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43092;
    wire N__43091;
    wire N__43090;
    wire N__43089;
    wire N__43088;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43064;
    wire N__43055;
    wire N__43050;
    wire N__43047;
    wire N__43046;
    wire N__43045;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43020;
    wire N__43019;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42972;
    wire N__42969;
    wire N__42966;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42945;
    wire N__42944;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42908;
    wire N__42905;
    wire N__42900;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42885;
    wire N__42882;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42842;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42824;
    wire N__42821;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42809;
    wire N__42808;
    wire N__42807;
    wire N__42804;
    wire N__42803;
    wire N__42802;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42747;
    wire N__42746;
    wire N__42743;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42729;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42721;
    wire N__42720;
    wire N__42717;
    wire N__42712;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42697;
    wire N__42692;
    wire N__42689;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42659;
    wire N__42658;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42639;
    wire N__42638;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42623;
    wire N__42620;
    wire N__42615;
    wire N__42614;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42599;
    wire N__42596;
    wire N__42591;
    wire N__42590;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42572;
    wire N__42569;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42533;
    wire N__42528;
    wire N__42525;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42510;
    wire N__42507;
    wire N__42506;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42492;
    wire N__42489;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42474;
    wire N__42471;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42449;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42435;
    wire N__42432;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42414;
    wire N__42411;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42393;
    wire N__42390;
    wire N__42389;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42376;
    wire N__42371;
    wire N__42366;
    wire N__42365;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42347;
    wire N__42342;
    wire N__42341;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42326;
    wire N__42323;
    wire N__42318;
    wire N__42315;
    wire N__42314;
    wire N__42313;
    wire N__42310;
    wire N__42307;
    wire N__42304;
    wire N__42301;
    wire N__42296;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42267;
    wire N__42264;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42252;
    wire N__42249;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42237;
    wire N__42234;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42222;
    wire N__42219;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42207;
    wire N__42204;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42168;
    wire N__42165;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42150;
    wire N__42147;
    wire N__42146;
    wire N__42145;
    wire N__42144;
    wire N__42137;
    wire N__42134;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42119;
    wire N__42118;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42101;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42074;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42060;
    wire N__42057;
    wire N__42056;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42042;
    wire N__42039;
    wire N__42038;
    wire N__42037;
    wire N__42034;
    wire N__42033;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42019;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42005;
    wire N__42002;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41966;
    wire N__41965;
    wire N__41962;
    wire N__41957;
    wire N__41952;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41942;
    wire N__41939;
    wire N__41934;
    wire N__41931;
    wire N__41930;
    wire N__41929;
    wire N__41926;
    wire N__41921;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41900;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41813;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41792;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41770;
    wire N__41763;
    wire N__41762;
    wire N__41759;
    wire N__41758;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41729;
    wire N__41728;
    wire N__41725;
    wire N__41720;
    wire N__41719;
    wire N__41714;
    wire N__41713;
    wire N__41710;
    wire N__41707;
    wire N__41704;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41687;
    wire N__41684;
    wire N__41681;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41576;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41505;
    wire N__41504;
    wire N__41501;
    wire N__41498;
    wire N__41493;
    wire N__41492;
    wire N__41491;
    wire N__41490;
    wire N__41487;
    wire N__41480;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41465;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41430;
    wire N__41427;
    wire N__41426;
    wire N__41421;
    wire N__41418;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41357;
    wire N__41356;
    wire N__41353;
    wire N__41348;
    wire N__41343;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41319;
    wire N__41316;
    wire N__41315;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41300;
    wire N__41297;
    wire N__41292;
    wire N__41289;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41281;
    wire N__41276;
    wire N__41273;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41261;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41228;
    wire N__41225;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41208;
    wire N__41205;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41167;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41151;
    wire N__41150;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41142;
    wire N__41139;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41125;
    wire N__41118;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41110;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41091;
    wire N__41088;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41080;
    wire N__41075;
    wire N__41072;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41057;
    wire N__41054;
    wire N__41051;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41034;
    wire N__41031;
    wire N__41030;
    wire N__41029;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41013;
    wire N__41010;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41002;
    wire N__40997;
    wire N__40994;
    wire N__40989;
    wire N__40986;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40962;
    wire N__40959;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40951;
    wire N__40946;
    wire N__40943;
    wire N__40938;
    wire N__40935;
    wire N__40934;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40917;
    wire N__40916;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40898;
    wire N__40895;
    wire N__40890;
    wire N__40887;
    wire N__40886;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40866;
    wire N__40865;
    wire N__40864;
    wire N__40861;
    wire N__40856;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40844;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40824;
    wire N__40823;
    wire N__40822;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40808;
    wire N__40807;
    wire N__40806;
    wire N__40805;
    wire N__40804;
    wire N__40803;
    wire N__40802;
    wire N__40801;
    wire N__40800;
    wire N__40799;
    wire N__40794;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40758;
    wire N__40753;
    wire N__40744;
    wire N__40735;
    wire N__40730;
    wire N__40727;
    wire N__40716;
    wire N__40713;
    wire N__40712;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40667;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40647;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40639;
    wire N__40634;
    wire N__40631;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40599;
    wire N__40598;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40554;
    wire N__40553;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40538;
    wire N__40535;
    wire N__40530;
    wire N__40527;
    wire N__40526;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40509;
    wire N__40508;
    wire N__40507;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40481;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40461;
    wire N__40460;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40426;
    wire N__40421;
    wire N__40418;
    wire N__40413;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40405;
    wire N__40400;
    wire N__40397;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40365;
    wire N__40364;
    wire N__40363;
    wire N__40360;
    wire N__40355;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40343;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40323;
    wire N__40322;
    wire N__40321;
    wire N__40318;
    wire N__40313;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40301;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40284;
    wire N__40281;
    wire N__40280;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40260;
    wire N__40257;
    wire N__40256;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40227;
    wire N__40224;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40216;
    wire N__40211;
    wire N__40208;
    wire N__40203;
    wire N__40202;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40184;
    wire N__40179;
    wire N__40176;
    wire N__40175;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40158;
    wire N__40155;
    wire N__40154;
    wire N__40153;
    wire N__40152;
    wire N__40151;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40127;
    wire N__40118;
    wire N__40113;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40105;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40086;
    wire N__40083;
    wire N__40082;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40065;
    wire N__40064;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40049;
    wire N__40046;
    wire N__40041;
    wire N__40038;
    wire N__40037;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40020;
    wire N__40019;
    wire N__40016;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__39998;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39974;
    wire N__39973;
    wire N__39972;
    wire N__39971;
    wire N__39970;
    wire N__39969;
    wire N__39968;
    wire N__39967;
    wire N__39966;
    wire N__39965;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39957;
    wire N__39956;
    wire N__39955;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39910;
    wire N__39905;
    wire N__39896;
    wire N__39887;
    wire N__39884;
    wire N__39875;
    wire N__39864;
    wire N__39863;
    wire N__39862;
    wire N__39861;
    wire N__39860;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39836;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39767;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39750;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39738;
    wire N__39737;
    wire N__39734;
    wire N__39731;
    wire N__39726;
    wire N__39723;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39708;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39652;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39624;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39612;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39597;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39585;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39566;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39549;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39534;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39522;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39510;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39498;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39483;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39455;
    wire N__39452;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39440;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39428;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39402;
    wire N__39401;
    wire N__39400;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39362;
    wire N__39361;
    wire N__39358;
    wire N__39353;
    wire N__39350;
    wire N__39347;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39329;
    wire N__39328;
    wire N__39327;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39311;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39299;
    wire N__39296;
    wire N__39295;
    wire N__39290;
    wire N__39289;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39277;
    wire N__39274;
    wire N__39269;
    wire N__39264;
    wire N__39261;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39249;
    wire N__39246;
    wire N__39245;
    wire N__39242;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39224;
    wire N__39219;
    wire N__39216;
    wire N__39215;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39191;
    wire N__39186;
    wire N__39183;
    wire N__39182;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39159;
    wire N__39156;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39134;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39116;
    wire N__39113;
    wire N__39112;
    wire N__39109;
    wire N__39104;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39089;
    wire N__39088;
    wire N__39085;
    wire N__39080;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39063;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39047;
    wire N__39042;
    wire N__39041;
    wire N__39040;
    wire N__39037;
    wire N__39032;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39022;
    wire N__39019;
    wire N__39014;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38993;
    wire N__38988;
    wire N__38985;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38973;
    wire N__38972;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38917;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38899;
    wire N__38896;
    wire N__38889;
    wire N__38886;
    wire N__38885;
    wire N__38882;
    wire N__38881;
    wire N__38878;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38762;
    wire N__38761;
    wire N__38760;
    wire N__38759;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38735;
    wire N__38726;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38708;
    wire N__38707;
    wire N__38706;
    wire N__38705;
    wire N__38704;
    wire N__38703;
    wire N__38702;
    wire N__38701;
    wire N__38700;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38692;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38652;
    wire N__38649;
    wire N__38640;
    wire N__38631;
    wire N__38628;
    wire N__38621;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38423;
    wire N__38422;
    wire N__38419;
    wire N__38414;
    wire N__38409;
    wire N__38408;
    wire N__38403;
    wire N__38400;
    wire N__38399;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38367;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38352;
    wire N__38349;
    wire N__38348;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38336;
    wire N__38335;
    wire N__38332;
    wire N__38327;
    wire N__38324;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38304;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38290;
    wire N__38289;
    wire N__38284;
    wire N__38279;
    wire N__38276;
    wire N__38271;
    wire N__38268;
    wire N__38267;
    wire N__38266;
    wire N__38263;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38238;
    wire N__38235;
    wire N__38234;
    wire N__38231;
    wire N__38230;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38218;
    wire N__38211;
    wire N__38210;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38202;
    wire N__38199;
    wire N__38194;
    wire N__38191;
    wire N__38184;
    wire N__38181;
    wire N__38180;
    wire N__38179;
    wire N__38174;
    wire N__38171;
    wire N__38166;
    wire N__38165;
    wire N__38160;
    wire N__38159;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38139;
    wire N__38136;
    wire N__38135;
    wire N__38132;
    wire N__38131;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38119;
    wire N__38112;
    wire N__38109;
    wire N__38108;
    wire N__38107;
    wire N__38104;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38094;
    wire N__38089;
    wire N__38086;
    wire N__38079;
    wire N__38078;
    wire N__38077;
    wire N__38076;
    wire N__38071;
    wire N__38066;
    wire N__38061;
    wire N__38060;
    wire N__38059;
    wire N__38058;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38040;
    wire N__38039;
    wire N__38034;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38022;
    wire N__38021;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38009;
    wire N__38008;
    wire N__38005;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37986;
    wire N__37983;
    wire N__37982;
    wire N__37977;
    wire N__37976;
    wire N__37975;
    wire N__37972;
    wire N__37967;
    wire N__37962;
    wire N__37959;
    wire N__37958;
    wire N__37957;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37945;
    wire N__37938;
    wire N__37935;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37927;
    wire N__37922;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37907;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37886;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37872;
    wire N__37869;
    wire N__37864;
    wire N__37859;
    wire N__37856;
    wire N__37851;
    wire N__37850;
    wire N__37847;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37823;
    wire N__37822;
    wire N__37821;
    wire N__37818;
    wire N__37813;
    wire N__37810;
    wire N__37805;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37784;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37773;
    wire N__37770;
    wire N__37765;
    wire N__37762;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37718;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37710;
    wire N__37705;
    wire N__37700;
    wire N__37695;
    wire N__37694;
    wire N__37693;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37671;
    wire N__37670;
    wire N__37667;
    wire N__37666;
    wire N__37665;
    wire N__37660;
    wire N__37655;
    wire N__37650;
    wire N__37649;
    wire N__37648;
    wire N__37647;
    wire N__37646;
    wire N__37643;
    wire N__37642;
    wire N__37639;
    wire N__37634;
    wire N__37627;
    wire N__37624;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37598;
    wire N__37597;
    wire N__37596;
    wire N__37595;
    wire N__37594;
    wire N__37593;
    wire N__37592;
    wire N__37589;
    wire N__37588;
    wire N__37587;
    wire N__37586;
    wire N__37583;
    wire N__37582;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37558;
    wire N__37551;
    wire N__37548;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37526;
    wire N__37523;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37512;
    wire N__37505;
    wire N__37502;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37485;
    wire N__37482;
    wire N__37481;
    wire N__37480;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37469;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37452;
    wire N__37443;
    wire N__37440;
    wire N__37439;
    wire N__37438;
    wire N__37437;
    wire N__37436;
    wire N__37435;
    wire N__37434;
    wire N__37431;
    wire N__37430;
    wire N__37423;
    wire N__37418;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37403;
    wire N__37400;
    wire N__37389;
    wire N__37386;
    wire N__37385;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37365;
    wire N__37364;
    wire N__37361;
    wire N__37360;
    wire N__37357;
    wire N__37352;
    wire N__37347;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37335;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37323;
    wire N__37320;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37305;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37256;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37224;
    wire N__37223;
    wire N__37218;
    wire N__37215;
    wire N__37214;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37182;
    wire N__37181;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37167;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37155;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37092;
    wire N__37091;
    wire N__37090;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37075;
    wire N__37068;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37056;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37044;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37029;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37014;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37002;
    wire N__36999;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36984;
    wire N__36981;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36969;
    wire N__36966;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36951;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36915;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36891;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36874;
    wire N__36869;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36843;
    wire N__36842;
    wire N__36841;
    wire N__36840;
    wire N__36835;
    wire N__36830;
    wire N__36825;
    wire N__36824;
    wire N__36821;
    wire N__36820;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36804;
    wire N__36803;
    wire N__36800;
    wire N__36799;
    wire N__36798;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36777;
    wire N__36774;
    wire N__36773;
    wire N__36770;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36748;
    wire N__36741;
    wire N__36740;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36723;
    wire N__36722;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36710;
    wire N__36705;
    wire N__36704;
    wire N__36703;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36691;
    wire N__36684;
    wire N__36683;
    wire N__36682;
    wire N__36681;
    wire N__36676;
    wire N__36671;
    wire N__36668;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36654;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36639;
    wire N__36638;
    wire N__36637;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36619;
    wire N__36612;
    wire N__36609;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36601;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36555;
    wire N__36550;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36534;
    wire N__36531;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36516;
    wire N__36515;
    wire N__36510;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36495;
    wire N__36494;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36479;
    wire N__36474;
    wire N__36471;
    wire N__36470;
    wire N__36467;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36444;
    wire N__36443;
    wire N__36442;
    wire N__36439;
    wire N__36436;
    wire N__36433;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36419;
    wire N__36418;
    wire N__36415;
    wire N__36410;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36398;
    wire N__36395;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36362;
    wire N__36359;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36309;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36297;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36282;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36251;
    wire N__36250;
    wire N__36249;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36197;
    wire N__36192;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36170;
    wire N__36165;
    wire N__36162;
    wire N__36161;
    wire N__36156;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36141;
    wire N__36138;
    wire N__36137;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36099;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36087;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36075;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36063;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36051;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36024;
    wire N__36023;
    wire N__36022;
    wire N__36021;
    wire N__36016;
    wire N__36011;
    wire N__36006;
    wire N__36005;
    wire N__36002;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35979;
    wire N__35978;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35963;
    wire N__35958;
    wire N__35957;
    wire N__35956;
    wire N__35953;
    wire N__35948;
    wire N__35943;
    wire N__35942;
    wire N__35941;
    wire N__35934;
    wire N__35931;
    wire N__35930;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35876;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35837;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35810;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35798;
    wire N__35795;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35764;
    wire N__35761;
    wire N__35756;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35738;
    wire N__35735;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35670;
    wire N__35667;
    wire N__35664;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35565;
    wire N__35562;
    wire N__35561;
    wire N__35556;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35529;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35514;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35502;
    wire N__35499;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35484;
    wire N__35481;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35466;
    wire N__35463;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35426;
    wire N__35425;
    wire N__35422;
    wire N__35417;
    wire N__35412;
    wire N__35411;
    wire N__35410;
    wire N__35405;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35352;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35311;
    wire N__35306;
    wire N__35303;
    wire N__35298;
    wire N__35295;
    wire N__35294;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35271;
    wire N__35268;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35256;
    wire N__35253;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35241;
    wire N__35238;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35226;
    wire N__35223;
    wire N__35222;
    wire N__35219;
    wire N__35216;
    wire N__35213;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35193;
    wire N__35190;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35178;
    wire N__35175;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35163;
    wire N__35160;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35109;
    wire N__35106;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire VCCG0;
    wire CLK_c;
    wire tx_enable;
    wire GB_BUFFER_PIN_9_c_THRU_CO;
    wire \quad_counter0.n28_adj_4414 ;
    wire \quad_counter0.n26_adj_4415 ;
    wire \quad_counter0.n25_adj_4417_cascade_ ;
    wire \quad_counter0.n27_adj_4416 ;
    wire \c0.n32768 ;
    wire \c0.n32756 ;
    wire \c0.n8_adj_4498 ;
    wire \c0.n8_adj_4494 ;
    wire bfn_4_10_0_;
    wire \quad_counter0.b_delay_counter_1 ;
    wire \quad_counter0.n30001 ;
    wire \quad_counter0.b_delay_counter_2 ;
    wire \quad_counter0.n30002 ;
    wire \quad_counter0.b_delay_counter_3 ;
    wire \quad_counter0.n30003 ;
    wire \quad_counter0.b_delay_counter_4 ;
    wire \quad_counter0.n30004 ;
    wire \quad_counter0.b_delay_counter_5 ;
    wire \quad_counter0.n30005 ;
    wire \quad_counter0.b_delay_counter_6 ;
    wire \quad_counter0.n30006 ;
    wire \quad_counter0.b_delay_counter_7 ;
    wire \quad_counter0.n30007 ;
    wire \quad_counter0.n30008 ;
    wire \quad_counter0.b_delay_counter_8 ;
    wire bfn_4_11_0_;
    wire \quad_counter0.b_delay_counter_9 ;
    wire \quad_counter0.n30009 ;
    wire \quad_counter0.b_delay_counter_10 ;
    wire \quad_counter0.n30010 ;
    wire \quad_counter0.b_delay_counter_11 ;
    wire \quad_counter0.n30011 ;
    wire \quad_counter0.b_delay_counter_12 ;
    wire \quad_counter0.n30012 ;
    wire \quad_counter0.b_delay_counter_13 ;
    wire \quad_counter0.n30013 ;
    wire \quad_counter0.b_delay_counter_14 ;
    wire \quad_counter0.n30014 ;
    wire \quad_counter0.n30015 ;
    wire \quad_counter0.b_delay_counter_15 ;
    wire quadB_delayed;
    wire PIN_8_c;
    wire b_delay_counter_15__N_4237_cascade_;
    wire n17987;
    wire n19282;
    wire n187;
    wire b_delay_counter_15__N_4237;
    wire n19282_cascade_;
    wire b_delay_counter_0;
    wire n3_cascade_;
    wire tx_o;
    wire \c0.n32792 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.n32786 ;
    wire \c0.n32780 ;
    wire \c0.n32774 ;
    wire \c0.n32834 ;
    wire \c0.n3_adj_4636_cascade_ ;
    wire \c0.n32710 ;
    wire \c0.n32816 ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n32828 ;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.n32822 ;
    wire bfn_5_11_0_;
    wire \c0.tx.n30068 ;
    wire \c0.tx.n30069 ;
    wire \c0.tx.n30070 ;
    wire \c0.tx.n30071 ;
    wire \c0.tx.n30072 ;
    wire \c0.tx.n30073 ;
    wire \c0.tx.n30074 ;
    wire \c0.tx.n30075 ;
    wire bfn_5_12_0_;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.n32810 ;
    wire \c0.n32722 ;
    wire \c0.n32734 ;
    wire \c0.n32716 ;
    wire \c0.n14_adj_4792 ;
    wire \c0.n15_adj_4793_cascade_ ;
    wire \c0.n63_cascade_ ;
    wire \c0.n118_adj_4786 ;
    wire \c0.n6_adj_4532 ;
    wire \c0.n15_adj_4796 ;
    wire \c0.n18_adj_4794_cascade_ ;
    wire \c0.n20_adj_4795 ;
    wire \c0.n18086 ;
    wire \c0.n115 ;
    wire data_in_2_7;
    wire data_in_0_7;
    wire data_in_0_2;
    wire data_in_0_6;
    wire data_in_1_7;
    wire \c0.n10_adj_4531 ;
    wire LED_c;
    wire a_delay_counter_15__N_4220_cascade_;
    wire \c0.tx.r_Clock_Count_0 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx.r_Clock_Count_1 ;
    wire \c0.r_Clock_Count_2 ;
    wire \c0.r_Clock_Count_4 ;
    wire \c0.n8_adj_4652_cascade_ ;
    wire n22210_cascade_;
    wire \c0.tx.n19946 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire \c0.tx.r_Clock_Count_7 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire \c0.tx.r_Clock_Count_8 ;
    wire \c0.n47_adj_4651 ;
    wire \c0.n10_adj_4504_cascade_ ;
    wire \c0.n35 ;
    wire r_Bit_Index_2;
    wire \c0.n32762 ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.n17_adj_4788_cascade_ ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n16_adj_4787 ;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n32840 ;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n45_adj_4637_cascade_ ;
    wire \c0.n32714 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire \c0.n32804 ;
    wire \c0.n32712 ;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.n8_adj_4496 ;
    wire \c0.n32798 ;
    wire data_in_1_4;
    wire data_in_0_4;
    wire data_in_0_1;
    wire data_in_0_5;
    wire data_in_1_6;
    wire data_in_3_7;
    wire \c0.n17_adj_4791_cascade_ ;
    wire \c0.n16_adj_4790 ;
    wire \c0.n18094 ;
    wire data_in_1_5;
    wire data_in_0_0;
    wire data_in_1_0;
    wire data_in_0_3;
    wire data_in_2_4;
    wire data_in_2_1;
    wire data_in_1_1;
    wire n27744;
    wire n4_adj_4808;
    wire a_delay_counter_0;
    wire n39;
    wire bfn_7_9_0_;
    wire \quad_counter0.a_delay_counter_1 ;
    wire \quad_counter0.n30016 ;
    wire \quad_counter0.a_delay_counter_2 ;
    wire \quad_counter0.n30017 ;
    wire \quad_counter0.a_delay_counter_3 ;
    wire \quad_counter0.n30018 ;
    wire \quad_counter0.a_delay_counter_4 ;
    wire \quad_counter0.n30019 ;
    wire \quad_counter0.a_delay_counter_5 ;
    wire \quad_counter0.n30020 ;
    wire \quad_counter0.n30021 ;
    wire \quad_counter0.n30022 ;
    wire \quad_counter0.n30023 ;
    wire \quad_counter0.a_delay_counter_8 ;
    wire bfn_7_10_0_;
    wire \quad_counter0.n30024 ;
    wire \quad_counter0.n30025 ;
    wire \quad_counter0.a_delay_counter_11 ;
    wire \quad_counter0.n30026 ;
    wire \quad_counter0.n30027 ;
    wire \quad_counter0.n30028 ;
    wire \quad_counter0.n30029 ;
    wire \quad_counter0.n30030 ;
    wire a_delay_counter_15__N_4220;
    wire \c0.n19530 ;
    wire \quad_counter0.a_delay_counter_10 ;
    wire \quad_counter0.a_delay_counter_14 ;
    wire \quad_counter0.a_delay_counter_15 ;
    wire \quad_counter0.a_delay_counter_7 ;
    wire \quad_counter0.a_delay_counter_13 ;
    wire \quad_counter0.a_delay_counter_9 ;
    wire \quad_counter0.a_delay_counter_6 ;
    wire \quad_counter0.a_delay_counter_12 ;
    wire \quad_counter0.n28_adj_4410 ;
    wire \quad_counter0.n27_adj_4412 ;
    wire \quad_counter0.n26_adj_4411_cascade_ ;
    wire \quad_counter0.n25_adj_4413 ;
    wire \c0.tx.n4_cascade_ ;
    wire \c0.tx.n22211 ;
    wire n19493;
    wire PIN_7_c;
    wire n15010;
    wire quadA_delayed;
    wire r_SM_Main_2_adj_4818;
    wire \c0.tx.n36215_cascade_ ;
    wire \c0.n36218 ;
    wire \c0.tx.n19358 ;
    wire r_SM_Main_1_adj_4819;
    wire n35927;
    wire n19509;
    wire n9_cascade_;
    wire n22210;
    wire r_SM_Main_0;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n32718 ;
    wire \c0.n79_cascade_ ;
    wire \c0.n4_adj_4613_cascade_ ;
    wire \c0.n8 ;
    wire \c0.n10_cascade_ ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.n19820_cascade_ ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n27824 ;
    wire \c0.n16_adj_4797 ;
    wire \c0.n15_adj_4798_cascade_ ;
    wire \c0.n19546 ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.n33163 ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.n12_adj_4789 ;
    wire \c0.n35771 ;
    wire \c0.n35698_cascade_ ;
    wire data_in_1_2;
    wire \c0.n33263_cascade_ ;
    wire data_in_3_6;
    wire data_in_2_6;
    wire data_in_3_2;
    wire data_in_2_2;
    wire \c0.n33266 ;
    wire \c0.n63 ;
    wire \c0.n107 ;
    wire \c0.n14_adj_4784 ;
    wire \c0.n13_adj_4785 ;
    wire data_in_3_3;
    wire data_in_2_3;
    wire data_in_1_3;
    wire data_in_3_0;
    wire data_in_2_0;
    wire \c0.data_in_frame_4_6 ;
    wire data_in_3_4;
    wire \c0.data_in_frame_9_6 ;
    wire \c0.n8_adj_4508_cascade_ ;
    wire \c0.n33985_cascade_ ;
    wire \c0.data_in_frame_7_1 ;
    wire \c0.n33444 ;
    wire \c0.data_in_frame_5_0 ;
    wire \c0.data_in_frame_9_2 ;
    wire bfn_9_7_0_;
    wire \quad_counter1.n30046 ;
    wire \quad_counter1.n30047 ;
    wire \quad_counter1.n30048 ;
    wire \quad_counter1.n30049 ;
    wire \quad_counter1.n30050 ;
    wire \quad_counter1.n30051 ;
    wire \quad_counter1.n30052 ;
    wire \quad_counter1.n30053 ;
    wire bfn_9_8_0_;
    wire \quad_counter1.n30054 ;
    wire \quad_counter1.n30055 ;
    wire \quad_counter1.n30056 ;
    wire \quad_counter1.n30057 ;
    wire \quad_counter1.n30058 ;
    wire \quad_counter1.n30059 ;
    wire \quad_counter1.n30060 ;
    wire rx_i;
    wire \quad_counter0.n25_adj_4367_cascade_ ;
    wire \quad_counter0.n27_adj_4366 ;
    wire \quad_counter0.n28_adj_4364 ;
    wire \quad_counter0.n26_adj_4365 ;
    wire \quad_counter0.n19 ;
    wire \quad_counter0.n28_adj_4361_cascade_ ;
    wire \quad_counter0.n24_adj_4360 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire \quad_counter0.n18_adj_4353_cascade_ ;
    wire \quad_counter0.n7_cascade_ ;
    wire \quad_counter0.n34617_cascade_ ;
    wire \quad_counter0.n22_adj_4355_cascade_ ;
    wire \quad_counter0.n26_adj_4356 ;
    wire bfn_9_13_0_;
    wire \quad_counter0.n30347 ;
    wire \quad_counter0.n30348 ;
    wire \quad_counter0.n30349 ;
    wire \quad_counter0.n30350 ;
    wire \quad_counter0.n30351 ;
    wire \quad_counter0.n30352 ;
    wire \quad_counter0.n30353 ;
    wire \quad_counter0.n30354 ;
    wire bfn_9_14_0_;
    wire \quad_counter0.n30355 ;
    wire \quad_counter0.n30356 ;
    wire \quad_counter0.n30357 ;
    wire \quad_counter0.n30358 ;
    wire \quad_counter0.n30359 ;
    wire \quad_counter0.n30360 ;
    wire \quad_counter0.n30361 ;
    wire \quad_counter0.n30362 ;
    wire bfn_9_15_0_;
    wire \quad_counter0.n30363 ;
    wire \quad_counter0.n30364 ;
    wire \quad_counter0.n36144 ;
    wire \quad_counter0.n24_adj_4354 ;
    wire \quad_counter0.n3035 ;
    wire \c0.n93 ;
    wire \quad_counter0.n20_adj_4351 ;
    wire \quad_counter0.n22_adj_4350_cascade_ ;
    wire \quad_counter0.n16 ;
    wire \quad_counter0.n24_adj_4352 ;
    wire \c0.n11_adj_4614 ;
    wire \c0.FRAME_MATCHER_state_2 ;
    wire \c0.n3844 ;
    wire \c0.n6_adj_4618 ;
    wire \c0.n33215_cascade_ ;
    wire \c0.n6_adj_4616 ;
    wire \c0.n33263 ;
    wire \c0.n29676 ;
    wire \c0.n10800 ;
    wire \c0.data_out_frame_0__7__N_2568 ;
    wire \c0.n22387 ;
    wire \c0.n10800_cascade_ ;
    wire \c0.n4_adj_4615 ;
    wire \c0.FRAME_MATCHER_state_1 ;
    wire \c0.data_in_frame_7_0 ;
    wire \c0.data_in_frame_9_1 ;
    wire \c0.data_in_frame_2_3 ;
    wire \c0.n6_adj_4564 ;
    wire \c0.n5452_cascade_ ;
    wire \c0.data_in_frame_4_5 ;
    wire \c0.n19030_cascade_ ;
    wire n4;
    wire \c0.data_in_frame_11_2 ;
    wire \c0.n33985 ;
    wire \c0.n33714_cascade_ ;
    wire \c0.n18671 ;
    wire \c0.n10_adj_4769_cascade_ ;
    wire \c0.data_in_frame_4_4 ;
    wire \c0.n18330_cascade_ ;
    wire \c0.data_in_frame_6_5 ;
    wire \c0.n33997 ;
    wire \c0.n33997_cascade_ ;
    wire \c0.data_in_frame_10_7 ;
    wire \quad_counter0.A_delayed ;
    wire A_filtered;
    wire \c0.n33695 ;
    wire \c0.data_in_frame_11_0 ;
    wire \c0.n6_adj_4713 ;
    wire B_filtered;
    wire \quad_counter0.B_delayed ;
    wire \c0.n33714 ;
    wire \c0.n33923 ;
    wire \c0.n33982_cascade_ ;
    wire \c0.data_in_frame_10_5 ;
    wire a_delay_counter_15__N_4220_adj_4817;
    wire n39_adj_4816;
    wire \quad_counter1.a_delay_counter_13 ;
    wire \quad_counter1.a_delay_counter_2 ;
    wire \quad_counter1.a_delay_counter_1 ;
    wire \quad_counter1.a_delay_counter_5 ;
    wire \quad_counter1.a_delay_counter_9 ;
    wire a_delay_counter_0_adj_4811;
    wire \quad_counter1.a_delay_counter_3 ;
    wire \quad_counter1.a_delay_counter_4 ;
    wire \quad_counter1.a_delay_counter_14 ;
    wire \quad_counter1.a_delay_counter_7 ;
    wire \quad_counter1.a_delay_counter_12 ;
    wire \quad_counter1.a_delay_counter_15 ;
    wire \quad_counter1.n25_adj_4443 ;
    wire \quad_counter1.n27_adj_4442_cascade_ ;
    wire \quad_counter1.n28_adj_4440 ;
    wire n17985_cascade_;
    wire n19433;
    wire \quad_counter1.a_delay_counter_11 ;
    wire \quad_counter1.a_delay_counter_6 ;
    wire \quad_counter1.a_delay_counter_10 ;
    wire \quad_counter1.a_delay_counter_8 ;
    wire \quad_counter1.n26_adj_4441 ;
    wire bfn_10_9_0_;
    wire \quad_counter0.n30384 ;
    wire \quad_counter0.n30385 ;
    wire \quad_counter0.n30386 ;
    wire \quad_counter0.n30387 ;
    wire \quad_counter0.n30388 ;
    wire \quad_counter0.n30389 ;
    wire \quad_counter0.n30390 ;
    wire \quad_counter0.n30391 ;
    wire bfn_10_10_0_;
    wire \quad_counter0.n30392 ;
    wire \quad_counter0.n30393 ;
    wire \quad_counter0.n30394 ;
    wire \quad_counter0.n30395 ;
    wire \quad_counter0.n30396 ;
    wire \quad_counter0.n30397 ;
    wire \quad_counter0.n30398 ;
    wire \quad_counter0.n30399 ;
    wire bfn_10_11_0_;
    wire \quad_counter0.n30400 ;
    wire \quad_counter0.n30401 ;
    wire \quad_counter0.n30402 ;
    wire \quad_counter0.n30403 ;
    wire \quad_counter0.n3233 ;
    wire \quad_counter0.n36141 ;
    wire \quad_counter0.n26_adj_4358 ;
    wire \quad_counter0.n16_adj_4359 ;
    wire bfn_10_12_0_;
    wire \quad_counter0.n3119 ;
    wire \quad_counter0.n30365 ;
    wire \quad_counter0.n3118 ;
    wire \quad_counter0.n30366 ;
    wire \quad_counter0.n3216 ;
    wire \quad_counter0.n30367 ;
    wire \quad_counter0.n3116 ;
    wire \quad_counter0.n3215 ;
    wire \quad_counter0.n30368 ;
    wire \quad_counter0.n3115 ;
    wire \quad_counter0.n30369 ;
    wire \quad_counter0.n36143 ;
    wire \quad_counter0.n3213 ;
    wire \quad_counter0.n30370 ;
    wire \quad_counter0.n3113 ;
    wire \quad_counter0.n3212 ;
    wire \quad_counter0.n30371 ;
    wire \quad_counter0.n30372 ;
    wire \quad_counter0.n3112 ;
    wire \quad_counter0.n3211 ;
    wire bfn_10_13_0_;
    wire \quad_counter0.n3111 ;
    wire \quad_counter0.n3210 ;
    wire \quad_counter0.n30373 ;
    wire \quad_counter0.n3110 ;
    wire \quad_counter0.n3209 ;
    wire \quad_counter0.n30374 ;
    wire \quad_counter0.n3109 ;
    wire \quad_counter0.n3208 ;
    wire \quad_counter0.n30375 ;
    wire \quad_counter0.n3108 ;
    wire \quad_counter0.n3207 ;
    wire \quad_counter0.n30376 ;
    wire \quad_counter0.n3107 ;
    wire \quad_counter0.n3206 ;
    wire \quad_counter0.n30377 ;
    wire \quad_counter0.n3106 ;
    wire \quad_counter0.n3205 ;
    wire \quad_counter0.n30378 ;
    wire \quad_counter0.n3105 ;
    wire \quad_counter0.n3204 ;
    wire \quad_counter0.n30379 ;
    wire \quad_counter0.n30380 ;
    wire \quad_counter0.n3104 ;
    wire \quad_counter0.n3203 ;
    wire bfn_10_14_0_;
    wire \quad_counter0.n3103 ;
    wire \quad_counter0.n3202 ;
    wire \quad_counter0.n30381 ;
    wire \quad_counter0.n3102 ;
    wire \quad_counter0.n3201 ;
    wire \quad_counter0.n30382 ;
    wire \quad_counter0.n3101 ;
    wire \quad_counter0.n3134 ;
    wire \quad_counter0.n30383 ;
    wire \quad_counter0.n3200 ;
    wire \c0.n93_adj_4634 ;
    wire bfn_10_15_0_;
    wire \quad_counter0.n30330 ;
    wire \quad_counter0.n30331 ;
    wire \quad_counter0.n3016 ;
    wire \quad_counter0.n30332 ;
    wire \quad_counter0.n3015 ;
    wire \quad_counter0.n30333 ;
    wire \quad_counter0.n30334 ;
    wire \quad_counter0.n3013 ;
    wire \quad_counter0.n30335 ;
    wire \quad_counter0.n3012 ;
    wire \quad_counter0.n30336 ;
    wire \quad_counter0.n30337 ;
    wire \quad_counter0.n3011 ;
    wire bfn_10_16_0_;
    wire \quad_counter0.n3010 ;
    wire \quad_counter0.n30338 ;
    wire \quad_counter0.n3009 ;
    wire \quad_counter0.n30339 ;
    wire \quad_counter0.n3008 ;
    wire \quad_counter0.n30340 ;
    wire \quad_counter0.n3007 ;
    wire \quad_counter0.n30341 ;
    wire \quad_counter0.n3006 ;
    wire \quad_counter0.n30342 ;
    wire \quad_counter0.n3005 ;
    wire \quad_counter0.n30343 ;
    wire \quad_counter0.n3004 ;
    wire \quad_counter0.n30344 ;
    wire \quad_counter0.n30345 ;
    wire \quad_counter0.n3003 ;
    wire bfn_10_17_0_;
    wire \quad_counter0.n30346 ;
    wire \quad_counter0.n3002 ;
    wire data_in_2_5;
    wire \c0.n33473 ;
    wire \c0.n33451 ;
    wire \c0.n6_adj_4503_cascade_ ;
    wire \c0.data_in_frame_2_4 ;
    wire \c0.n19030 ;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.n33386 ;
    wire \c0.n33386_cascade_ ;
    wire \c0.data_in_frame_4_7 ;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.data_in_frame_3_1 ;
    wire \c0.n33720_cascade_ ;
    wire \c0.n17559_cascade_ ;
    wire \c0.data_in_frame_9_5 ;
    wire \c0.n18544_cascade_ ;
    wire \c0.n31505_cascade_ ;
    wire \c0.n4_adj_4548 ;
    wire \c0.n43_adj_4732_cascade_ ;
    wire \c0.n33778 ;
    wire \c0.n46_adj_4728 ;
    wire \c0.n47_adj_4729 ;
    wire \c0.n45_adj_4730_cascade_ ;
    wire \c0.n54 ;
    wire \c0.n17559 ;
    wire \c0.n48 ;
    wire \c0.n6_adj_4556_cascade_ ;
    wire \c0.n33404 ;
    wire \c0.n12_adj_4735_cascade_ ;
    wire \c0.n31526_cascade_ ;
    wire \c0.n33624 ;
    wire \c0.n5860 ;
    wire \c0.n33883 ;
    wire \c0.n44_adj_4731 ;
    wire \c0.n33800 ;
    wire \c0.data_in_frame_11_6 ;
    wire \c0.data_in_frame_9_4 ;
    wire \c0.n33641 ;
    wire \c0.data_in_frame_7_3 ;
    wire \c0.n31505 ;
    wire \c0.n33641_cascade_ ;
    wire \c0.n33836 ;
    wire \c0.n6_adj_4557 ;
    wire \c0.n33982 ;
    wire \c0.n18_adj_4725_cascade_ ;
    wire \c0.n33951 ;
    wire \c0.n16_adj_4726 ;
    wire \c0.n20_adj_4727_cascade_ ;
    wire \c0.data_in_frame_8_6 ;
    wire \c0.data_in_frame_8_4 ;
    wire \c0.n33723 ;
    wire \c0.n33723_cascade_ ;
    wire \c0.data_in_frame_12_7 ;
    wire \c0.data_in_frame_10_6 ;
    wire \c0.n6_adj_4539_cascade_ ;
    wire \c0.n19199_cascade_ ;
    wire \c0.data_in_frame_11_4 ;
    wire \c0.data_in_frame_11_3 ;
    wire PIN_13_c;
    wire quadB_delayed_adj_4813;
    wire \quad_counter1.n26_adj_4447_cascade_ ;
    wire n17983;
    wire \quad_counter1.n27_adj_4448 ;
    wire \quad_counter1.n25_adj_4449 ;
    wire \quad_counter1.n28_adj_4446 ;
    wire \quad_counter1.b_delay_counter_0 ;
    wire bfn_11_7_0_;
    wire \quad_counter1.b_delay_counter_1 ;
    wire \quad_counter1.n30031 ;
    wire \quad_counter1.b_delay_counter_2 ;
    wire \quad_counter1.n30032 ;
    wire \quad_counter1.b_delay_counter_3 ;
    wire \quad_counter1.n30033 ;
    wire \quad_counter1.b_delay_counter_4 ;
    wire \quad_counter1.n30034 ;
    wire \quad_counter1.b_delay_counter_5 ;
    wire \quad_counter1.n30035 ;
    wire \quad_counter1.b_delay_counter_6 ;
    wire \quad_counter1.n30036 ;
    wire \quad_counter1.b_delay_counter_7 ;
    wire \quad_counter1.n30037 ;
    wire \quad_counter1.n30038 ;
    wire \quad_counter1.b_delay_counter_8 ;
    wire bfn_11_8_0_;
    wire \quad_counter1.b_delay_counter_9 ;
    wire \quad_counter1.n30039 ;
    wire \quad_counter1.b_delay_counter_10 ;
    wire \quad_counter1.n30040 ;
    wire \quad_counter1.b_delay_counter_11 ;
    wire \quad_counter1.n30041 ;
    wire \quad_counter1.b_delay_counter_12 ;
    wire \quad_counter1.n30042 ;
    wire \quad_counter1.b_delay_counter_13 ;
    wire \quad_counter1.n30043 ;
    wire \quad_counter1.b_delay_counter_14 ;
    wire \quad_counter1.n30044 ;
    wire \quad_counter1.n30045 ;
    wire \quad_counter1.b_delay_counter_15 ;
    wire n19463;
    wire \quad_counter1.b_delay_counter_15__N_4237 ;
    wire \quad_counter0.n3219 ;
    wire \quad_counter0.n3218 ;
    wire \quad_counter0.n3217 ;
    wire \quad_counter0.n28297_cascade_ ;
    wire \quad_counter0.n3214 ;
    wire \quad_counter0.n10_adj_4357 ;
    wire \quad_counter0.n3019 ;
    wire \quad_counter0.n10_adj_4376_cascade_ ;
    wire \quad_counter0.n1847_cascade_ ;
    wire r_Bit_Index_1;
    wire r_Tx_Data_4;
    wire r_Bit_Index_0;
    wire \c0.n36167 ;
    wire \c0.n36170 ;
    wire \c0.n10_adj_4629 ;
    wire \quad_counter0.n3018 ;
    wire \quad_counter0.n3014 ;
    wire \quad_counter0.n3017 ;
    wire \quad_counter0.n28307 ;
    wire \quad_counter0.n10_adj_4349 ;
    wire r_Tx_Data_2;
    wire data_in_3_5;
    wire r_Tx_Data_1;
    wire \c0.n11057 ;
    wire bfn_11_14_0_;
    wire \quad_counter0.n30314 ;
    wire \quad_counter0.n30315 ;
    wire \quad_counter0.n30316 ;
    wire \quad_counter0.n30317 ;
    wire \quad_counter0.n30318 ;
    wire \quad_counter0.n30319 ;
    wire \quad_counter0.n30320 ;
    wire \quad_counter0.n30321 ;
    wire bfn_11_15_0_;
    wire \quad_counter0.n30322 ;
    wire \quad_counter0.n30323 ;
    wire \quad_counter0.n30324 ;
    wire \quad_counter0.n30325 ;
    wire \quad_counter0.n30326 ;
    wire \quad_counter0.n30327 ;
    wire \quad_counter0.n30328 ;
    wire \quad_counter0.n30329 ;
    wire bfn_11_16_0_;
    wire \quad_counter0.n36147 ;
    wire \quad_counter0.n2908 ;
    wire \quad_counter0.n2904 ;
    wire \quad_counter0.n2910 ;
    wire \quad_counter0.n2913 ;
    wire \quad_counter0.n2907 ;
    wire \quad_counter0.n2905 ;
    wire \quad_counter0.n2919 ;
    wire \quad_counter0.n36145 ;
    wire \quad_counter0.n2912 ;
    wire \quad_counter0.n2903 ;
    wire \quad_counter0.n20 ;
    wire \quad_counter0.n2909 ;
    wire \quad_counter0.n2911 ;
    wire \quad_counter0.n22_cascade_ ;
    wire \quad_counter0.n18 ;
    wire \quad_counter0.n2936 ;
    wire \quad_counter0.n2917 ;
    wire \quad_counter0.n2918 ;
    wire \quad_counter0.n2914 ;
    wire \quad_counter0.n28315 ;
    wire \quad_counter0.n2916 ;
    wire \quad_counter0.n2915 ;
    wire \quad_counter0.n10_adj_4348_cascade_ ;
    wire \quad_counter0.n2906 ;
    wire \quad_counter0.n13 ;
    wire \c0.n33454 ;
    wire \c0.n33720 ;
    wire \c0.n33341 ;
    wire \c0.n14_adj_4771 ;
    wire \c0.n13_adj_4773 ;
    wire \c0.n14_adj_4772_cascade_ ;
    wire \c0.n13_adj_4774 ;
    wire \c0.data_in_frame_8_5 ;
    wire \c0.n49 ;
    wire \c0.data_in_frame_11_1 ;
    wire \c0.n33476 ;
    wire \c0.n19102_cascade_ ;
    wire \c0.data_in_frame_11_5 ;
    wire \c0.data_out_frame_0__7__N_2744 ;
    wire \c0.n33650 ;
    wire \c0.n32325 ;
    wire \c0.n33311 ;
    wire \c0.n33311_cascade_ ;
    wire \c0.data_in_frame_0_4 ;
    wire \c0.data_in_frame_11_7 ;
    wire \c0.n33523 ;
    wire \c0.n18544 ;
    wire \c0.data_in_frame_7_5 ;
    wire \c0.n33954 ;
    wire \c0.n34003_cascade_ ;
    wire \c0.n33758 ;
    wire \c0.data_in_frame_15_5 ;
    wire \c0.n33781 ;
    wire \c0.n18847_cascade_ ;
    wire \c0.n10_adj_4708 ;
    wire \c0.data_in_frame_8_7 ;
    wire \c0.n19102 ;
    wire \c0.n33729 ;
    wire \c0.n33729_cascade_ ;
    wire \c0.n14_adj_4582 ;
    wire \c0.n34000 ;
    wire \c0.n19190 ;
    wire \c0.n15998 ;
    wire \c0.data_in_frame_7_2 ;
    wire \c0.data_in_frame_15_4 ;
    wire \c0.n33908_cascade_ ;
    wire \c0.n30_adj_4737 ;
    wire \c0.data_in_frame_15_0 ;
    wire \c0.data_in_frame_14_6 ;
    wire \c0.n17582 ;
    wire \c0.n18511 ;
    wire \c0.n33554 ;
    wire \c0.n33824_cascade_ ;
    wire \c0.n24_adj_4722_cascade_ ;
    wire \c0.n26_adj_4724_cascade_ ;
    wire \c0.n22_adj_4723 ;
    wire \c0.n33 ;
    wire \c0.n34_adj_4738 ;
    wire \c0.n32_adj_4739 ;
    wire \c0.data_in_frame_17_2 ;
    wire \c0.data_in_frame_17_4 ;
    wire \c0.data_in_frame_14_7 ;
    wire \quad_counter0.n28397_cascade_ ;
    wire bfn_12_7_0_;
    wire \quad_counter0.n1847 ;
    wire \quad_counter0.n30209 ;
    wire \quad_counter0.n30210 ;
    wire \quad_counter0.n30211 ;
    wire \quad_counter0.n30212 ;
    wire \quad_counter0.n30213 ;
    wire \quad_counter0.n36158 ;
    wire \quad_counter0.n30214 ;
    wire PIN_12_c;
    wire n17985;
    wire quadA_delayed_adj_4812;
    wire bfn_12_9_0_;
    wire \quad_counter0.n30404 ;
    wire \quad_counter0.n30405 ;
    wire \quad_counter0.n30406 ;
    wire \quad_counter0.n30407 ;
    wire \quad_counter0.n30408 ;
    wire \quad_counter0.n36140 ;
    wire \quad_counter0.n30409 ;
    wire \quad_counter0.n3313 ;
    wire \quad_counter0.n30410 ;
    wire \quad_counter0.n30411 ;
    wire \quad_counter0.n3312 ;
    wire bfn_12_10_0_;
    wire \quad_counter0.n3311 ;
    wire \quad_counter0.n30412 ;
    wire \quad_counter0.n3310 ;
    wire \quad_counter0.n30413 ;
    wire \quad_counter0.n3309 ;
    wire \quad_counter0.n30414 ;
    wire \quad_counter0.n3308 ;
    wire \quad_counter0.n30415 ;
    wire \quad_counter0.n3307 ;
    wire \quad_counter0.n30416 ;
    wire \quad_counter0.n3306 ;
    wire \quad_counter0.n30417 ;
    wire \quad_counter0.n3305 ;
    wire \quad_counter0.n30418 ;
    wire \quad_counter0.n30419 ;
    wire \quad_counter0.n3304 ;
    wire bfn_12_11_0_;
    wire \quad_counter0.n3303 ;
    wire \quad_counter0.n30420 ;
    wire \quad_counter0.n3302 ;
    wire \quad_counter0.n30421 ;
    wire \quad_counter0.n3301 ;
    wire \quad_counter0.n30422 ;
    wire \quad_counter0.n3300 ;
    wire \quad_counter0.n30423 ;
    wire \quad_counter0.n3299 ;
    wire \quad_counter0.n3332 ;
    wire \quad_counter0.n30424 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire \c0.n32730 ;
    wire bfn_12_13_0_;
    wire \quad_counter0.n30299 ;
    wire \quad_counter0.n30300 ;
    wire \quad_counter0.n30301 ;
    wire \quad_counter0.n30302 ;
    wire \quad_counter0.n30303 ;
    wire \quad_counter0.n30304 ;
    wire \quad_counter0.n30305 ;
    wire \quad_counter0.n30306 ;
    wire bfn_12_14_0_;
    wire \quad_counter0.n30307 ;
    wire \quad_counter0.n30308 ;
    wire \quad_counter0.n30309 ;
    wire \quad_counter0.n30310 ;
    wire \quad_counter0.n30311 ;
    wire \quad_counter0.n30312 ;
    wire \quad_counter0.n30313 ;
    wire \quad_counter0.n2813 ;
    wire \quad_counter0.n2811 ;
    wire \quad_counter0.n2810 ;
    wire \quad_counter0.n2807 ;
    wire \quad_counter0.n2808 ;
    wire \quad_counter0.n2812 ;
    wire \quad_counter0.n2805 ;
    wire \quad_counter0.n2804 ;
    wire \quad_counter0.n2806 ;
    wire \quad_counter0.n19_adj_4409_cascade_ ;
    wire \quad_counter0.n18_adj_4408 ;
    wire \quad_counter0.n2837 ;
    wire \quad_counter0.n2819 ;
    wire \quad_counter0.n2817 ;
    wire \quad_counter0.n2818 ;
    wire \quad_counter0.n28323_cascade_ ;
    wire \quad_counter0.n2814 ;
    wire \quad_counter0.n2816 ;
    wire \quad_counter0.n2815 ;
    wire \quad_counter0.n10_adj_4406_cascade_ ;
    wire \quad_counter0.n2809 ;
    wire \quad_counter0.n12_adj_4407 ;
    wire \c0.n32740 ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n33160 ;
    wire \c0.n19909_cascade_ ;
    wire \c0.data_out_frame_29_7_N_2879_2 ;
    wire \c0.n34017_cascade_ ;
    wire \c0.n29675_cascade_ ;
    wire \c0.n81_cascade_ ;
    wire \c0.n99 ;
    wire \c0.n3_adj_4636 ;
    wire \c0.n45_adj_4637 ;
    wire \c0.n29_adj_4776 ;
    wire \c0.n9_adj_4509 ;
    wire \c0.n34 ;
    wire \c0.n18330 ;
    wire \c0.n20_adj_4534 ;
    wire \c0.n28_adj_4777_cascade_ ;
    wire \c0.n32_adj_4778 ;
    wire \c0.n27710_cascade_ ;
    wire \c0.n35947_cascade_ ;
    wire \c0.n35808 ;
    wire \c0.n38_adj_4780_cascade_ ;
    wire \c0.n35804 ;
    wire \c0.n46_adj_4783_cascade_ ;
    wire \c0.data_in_frame_2_7 ;
    wire \c0.n39_adj_4781 ;
    wire \c0.n37_adj_4782 ;
    wire \c0.data_in_frame_0_5 ;
    wire \c0.n10_adj_4768 ;
    wire n18026;
    wire \c0.data_in_frame_6_6 ;
    wire \c0.data_out_frame_0__7__N_2747 ;
    wire \c0.n26_adj_4775 ;
    wire \c0.n33582 ;
    wire \c0.n33291_cascade_ ;
    wire \c0.n19_adj_4779 ;
    wire \c0.data_in_frame_2_6 ;
    wire \c0.data_in_frame_5_6 ;
    wire \c0.data_in_frame_6_7 ;
    wire \c0.n6_adj_4501_cascade_ ;
    wire \c0.data_in_frame_3_2 ;
    wire \c0.data_in_frame_5_5 ;
    wire \c0.n6_cascade_ ;
    wire \c0.n18141_cascade_ ;
    wire \c0.data_in_frame_3_3 ;
    wire \c0.n33927_cascade_ ;
    wire \c0.data_in_frame_10_2 ;
    wire \c0.n31439 ;
    wire \c0.data_in_frame_14_1 ;
    wire \c0.n2_adj_4741 ;
    wire \c0.n2_adj_4741_cascade_ ;
    wire \c0.n33283 ;
    wire \c0.data_in_frame_8_1 ;
    wire \c0.n33283_cascade_ ;
    wire \c0.n33871 ;
    wire \c0.data_in_frame_18_3 ;
    wire \c0.data_in_frame_14_5 ;
    wire \c0.data_in_frame_6_1 ;
    wire \c0.n18364 ;
    wire \c0.n33880_cascade_ ;
    wire \c0.data_in_frame_18_2 ;
    wire \c0.n12_adj_4716_cascade_ ;
    wire \c0.n33741 ;
    wire \c0.n18368 ;
    wire \c0.n33741_cascade_ ;
    wire \c0.n33880 ;
    wire \c0.data_in_frame_17_7 ;
    wire \c0.n33711 ;
    wire \c0.n5896 ;
    wire \c0.n34_adj_4718_cascade_ ;
    wire \c0.n37_adj_4720 ;
    wire \c0.n35_adj_4721 ;
    wire \c0.n38_adj_4719_cascade_ ;
    wire \c0.data_in_frame_16_1 ;
    wire \c0.n34003 ;
    wire \c0.n24_adj_4717 ;
    wire \c0.data_in_frame_18_0 ;
    wire \c0.n33371 ;
    wire \c0.n10_adj_4697 ;
    wire \c0.n33356 ;
    wire \c0.n18588_cascade_ ;
    wire \c0.n33789 ;
    wire \c0.n33789_cascade_ ;
    wire \c0.n19108_cascade_ ;
    wire \c0.n18431 ;
    wire \c0.n33886 ;
    wire \c0.data_in_frame_17_5 ;
    wire \c0.n8_adj_4745 ;
    wire \c0.n6242_cascade_ ;
    wire \c0.n33665_cascade_ ;
    wire \c0.data_in_frame_19_0 ;
    wire \c0.data_in_frame_20_0 ;
    wire \c0.n19199 ;
    wire \c0.n31589 ;
    wire \c0.n33514_cascade_ ;
    wire \c0.n19226 ;
    wire \c0.n12_adj_4696 ;
    wire \c0.n33717 ;
    wire \c0.data_in_frame_19_1 ;
    wire \c0.n33308 ;
    wire \c0.n33735 ;
    wire \c0.n33308_cascade_ ;
    wire \c0.n36 ;
    wire \c0.data_in_frame_19_7 ;
    wire \c0.n22_adj_4574 ;
    wire \c0.data_in_frame_20_1 ;
    wire \c0.n33945 ;
    wire \quad_counter0.n10_adj_4377 ;
    wire \quad_counter0.n1946_cascade_ ;
    wire \quad_counter0.n2019_cascade_ ;
    wire \quad_counter0.n1987 ;
    wire bfn_13_7_0_;
    wire \quad_counter0.n30215 ;
    wire \quad_counter0.n30216 ;
    wire \quad_counter0.n1917 ;
    wire \quad_counter0.n1984 ;
    wire \quad_counter0.n30217 ;
    wire \quad_counter0.n1916 ;
    wire \quad_counter0.n1983 ;
    wire \quad_counter0.n30218 ;
    wire \quad_counter0.n30219 ;
    wire \quad_counter0.n1914 ;
    wire \quad_counter0.n1981 ;
    wire \quad_counter0.n30220 ;
    wire \quad_counter0.n1913 ;
    wire \quad_counter0.n30221 ;
    wire \quad_counter0.n3316 ;
    wire \quad_counter0.n3315 ;
    wire \quad_counter0.n35311 ;
    wire \quad_counter0.n3317 ;
    wire \quad_counter0.n3314 ;
    wire \quad_counter0.n8_adj_4362 ;
    wire \quad_counter0.n8_adj_4369_cascade_ ;
    wire \quad_counter0.n3319 ;
    wire \quad_counter0.n3318 ;
    wire \quad_counter0.n7_adj_4363 ;
    wire \quad_counter0.n7_adj_4370 ;
    wire \quad_counter0.n18_adj_4368_cascade_ ;
    wire \quad_counter0.n34805 ;
    wire \quad_counter0.n7_adj_4395 ;
    wire \quad_counter0.n28331_cascade_ ;
    wire \quad_counter0.n10_adj_4402_cascade_ ;
    wire \quad_counter0.n16_adj_4403 ;
    wire \quad_counter0.n14_adj_4404 ;
    wire \quad_counter0.n18_adj_4405_cascade_ ;
    wire \quad_counter0.n2738 ;
    wire \quad_counter0.n2738_cascade_ ;
    wire \quad_counter0.n36149 ;
    wire \c0.n31012 ;
    wire \c0.n111 ;
    wire \c0.data_out_frame_0__7__N_2569_cascade_ ;
    wire \c0.n33170 ;
    wire r_SM_Main_2_N_3755_0;
    wire \c0.tx_active ;
    wire \c0.n35938 ;
    wire \c0.n6_adj_4638 ;
    wire \c0.n35339 ;
    wire \c0.n14779_cascade_ ;
    wire \c0.n6_adj_4617 ;
    wire \c0.n18115 ;
    wire \c0.n33166 ;
    wire \c0.n19820 ;
    wire \c0.n14779 ;
    wire \c0.data_out_frame_0__7__N_2569 ;
    wire \c0.n688 ;
    wire \c0.n118 ;
    wire \c0.n30958 ;
    wire \c0.n18100 ;
    wire \c0.n18100_cascade_ ;
    wire \c0.n18045 ;
    wire \c0.n4_adj_4537_cascade_ ;
    wire \c0.n18020_cascade_ ;
    wire \c0.n35757_cascade_ ;
    wire \c0.n79 ;
    wire \c0.n47_adj_4611_cascade_ ;
    wire \c0.n58 ;
    wire \c0.n4_adj_4612 ;
    wire data_in_3_1;
    wire \c0.n19909 ;
    wire \c0.n30862 ;
    wire \c0.n4_adj_4537 ;
    wire \c0.n30862_cascade_ ;
    wire \c0.n72 ;
    wire \c0.n29668 ;
    wire \c0.FRAME_MATCHER_state_0 ;
    wire \c0.n72_cascade_ ;
    wire \c0.n11851 ;
    wire \c0.data_out_frame_0__7__N_2570 ;
    wire \c0.n18675_cascade_ ;
    wire \c0.n5_adj_4545 ;
    wire \c0.n18667 ;
    wire \c0.n18667_cascade_ ;
    wire \c0.n33347 ;
    wire \c0.n18319 ;
    wire \c0.data_in_frame_0_0 ;
    wire \c0.data_in_frame_2_2 ;
    wire \c0.n35806 ;
    wire \c0.data_in_frame_0_6 ;
    wire \c0.n18354 ;
    wire \c0.n33326 ;
    wire \c0.n33804 ;
    wire \c0.n18354_cascade_ ;
    wire \c0.n31_adj_4766 ;
    wire \c0.n30_adj_4765 ;
    wire \c0.n29_adj_4767_cascade_ ;
    wire \c0.n33830 ;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.n33830_cascade_ ;
    wire \c0.n6_adj_4535 ;
    wire \c0.n18709 ;
    wire \c0.data_in_frame_7_4 ;
    wire \c0.data_in_frame_10_0 ;
    wire \c0.n8_adj_4555_cascade_ ;
    wire \c0.n7_adj_4554 ;
    wire \c0.n33441_cascade_ ;
    wire \c0.data_in_frame_7_7 ;
    wire \c0.n18141 ;
    wire \c0.data_in_frame_7_6 ;
    wire \c0.n6_adj_4733 ;
    wire \c0.n32298 ;
    wire \c0.data_in_frame_9_7 ;
    wire \c0.data_in_frame_10_1 ;
    wire \c0.n33698 ;
    wire \c0.n10_adj_4736 ;
    wire \c0.n33708 ;
    wire \c0.n33877 ;
    wire \c0.data_in_frame_4_2 ;
    wire \c0.data_in_frame_14_2 ;
    wire \c0.data_in_frame_8_0 ;
    wire \c0.data_in_frame_10_4 ;
    wire \c0.data_in_frame_12_5 ;
    wire \c0.n33874_cascade_ ;
    wire \c0.data_out_frame_0__7__N_2580 ;
    wire \c0.n5_adj_4742 ;
    wire \c0.n33288 ;
    wire \c0.n18705 ;
    wire \c0.data_in_frame_8_2 ;
    wire \c0.n18705_cascade_ ;
    wire \c0.n33291 ;
    wire \c0.n10_adj_4743 ;
    wire \c0.n33705 ;
    wire \c0.n10_adj_4744 ;
    wire \c0.data_in_frame_8_3 ;
    wire \c0.n33874 ;
    wire \c0.n19064 ;
    wire \c0.data_in_frame_13_2 ;
    wire \c0.data_in_frame_13_3 ;
    wire \c0.n18373_cascade_ ;
    wire \c0.n5965 ;
    wire \c0.n4_adj_4734 ;
    wire \c0.n5965_cascade_ ;
    wire \c0.data_in_frame_17_6 ;
    wire \c0.data_in_frame_10_3 ;
    wire \c0.n5996 ;
    wire \c0.n18290 ;
    wire \c0.data_in_frame_12_6 ;
    wire \c0.n18147 ;
    wire \c0.data_in_frame_12_0 ;
    wire \c0.n18_adj_4563 ;
    wire \c0.data_in_frame_19_4 ;
    wire \c0.n18582 ;
    wire \c0.data_in_frame_17_1 ;
    wire \c0.data_in_frame_12_3 ;
    wire \c0.n33545 ;
    wire \c0.n33545_cascade_ ;
    wire \c0.n35505_cascade_ ;
    wire \c0.data_in_frame_18_7 ;
    wire \c0.data_in_frame_18_6 ;
    wire \c0.n33852_cascade_ ;
    wire \c0.n33942 ;
    wire \c0.n10_adj_4575 ;
    wire \c0.n33647 ;
    wire \c0.n10_adj_4575_cascade_ ;
    wire \c0.n32302 ;
    wire \c0.n32390_cascade_ ;
    wire \c0.data_in_frame_23_0 ;
    wire bfn_14_5_0_;
    wire \quad_counter0.n30222 ;
    wire \quad_counter0.n30223 ;
    wire \quad_counter0.n30224 ;
    wire \quad_counter0.n30225 ;
    wire \quad_counter0.n30226 ;
    wire \quad_counter0.n30227 ;
    wire \quad_counter0.n30228 ;
    wire \quad_counter0.n30229 ;
    wire bfn_14_6_0_;
    wire \quad_counter0.n2087 ;
    wire \quad_counter0.n2119_cascade_ ;
    wire \quad_counter0.n1985 ;
    wire \quad_counter0.n1918 ;
    wire \quad_counter0.n2080 ;
    wire \quad_counter0.n1982 ;
    wire \quad_counter0.n1915 ;
    wire \quad_counter0.n2014_cascade_ ;
    wire \quad_counter0.n28371 ;
    wire \quad_counter0.n2012 ;
    wire \quad_counter0.n2013 ;
    wire \quad_counter0.n10_adj_4378_cascade_ ;
    wire \quad_counter0.n2019 ;
    wire \quad_counter0.n2045_cascade_ ;
    wire \quad_counter0.n2086 ;
    wire \quad_counter0.n9_adj_4379 ;
    wire \quad_counter0.n30_cascade_ ;
    wire \quad_counter0.n28291_cascade_ ;
    wire \quad_counter0.n10_cascade_ ;
    wire \quad_counter0.n21 ;
    wire \quad_counter0.n34759 ;
    wire \quad_counter0.n12 ;
    wire \quad_counter0.n30_adj_4371 ;
    wire \quad_counter0.n29_adj_4373 ;
    wire \quad_counter0.n28_adj_4372 ;
    wire \quad_counter0.n27_adj_4374 ;
    wire \quad_counter0.n2719 ;
    wire bfn_14_11_0_;
    wire \quad_counter0.n2718 ;
    wire \quad_counter0.n30285 ;
    wire \quad_counter0.n2717 ;
    wire \quad_counter0.n30286 ;
    wire \quad_counter0.n2716 ;
    wire \quad_counter0.n30287 ;
    wire \quad_counter0.n2715 ;
    wire \quad_counter0.n30288 ;
    wire \quad_counter0.n2714 ;
    wire \quad_counter0.n30289 ;
    wire \quad_counter0.n2713 ;
    wire \quad_counter0.n30290 ;
    wire \quad_counter0.n2712 ;
    wire \quad_counter0.n30291 ;
    wire \quad_counter0.n30292 ;
    wire \quad_counter0.n2711 ;
    wire bfn_14_12_0_;
    wire \quad_counter0.n2710 ;
    wire \quad_counter0.n30293 ;
    wire \quad_counter0.n2709 ;
    wire \quad_counter0.n30294 ;
    wire \quad_counter0.n2708 ;
    wire \quad_counter0.n30295 ;
    wire \quad_counter0.n2707 ;
    wire \quad_counter0.n30296 ;
    wire \quad_counter0.n2706 ;
    wire \quad_counter0.n30297 ;
    wire \quad_counter0.n30298 ;
    wire \quad_counter0.n2705 ;
    wire \quad_counter0.n12_adj_4396 ;
    wire \quad_counter0.n2441_cascade_ ;
    wire r_Tx_Data_6;
    wire \c0.tx_transmit_N_3651 ;
    wire bfn_14_14_0_;
    wire \c0.n30202 ;
    wire \c0.n30203 ;
    wire \c0.n30204 ;
    wire \c0.n30205 ;
    wire \c0.n30206 ;
    wire \c0.n30207 ;
    wire \c0.n30208 ;
    wire \c0.n19388 ;
    wire \c0.n29678 ;
    wire data_out_frame_29__7__N_1482_cascade_;
    wire n10_adj_4805;
    wire \c0.n17961 ;
    wire \c0.n29675 ;
    wire \c0.n78 ;
    wire \c0.data_out_frame_0__7__N_2571 ;
    wire \c0.data_out_frame_0_2 ;
    wire \c0.n35960_cascade_ ;
    wire \c0.n6_adj_4510_cascade_ ;
    wire \c0.data_out_frame_0_3 ;
    wire data_out_frame_5_2;
    wire data_out_frame_6_0;
    wire data_out_frame_7_0;
    wire \c0.n27710 ;
    wire \c0.n34190 ;
    wire \c0.data_out_frame_29_7_N_1483_0 ;
    wire \c0.n12_cascade_ ;
    wire \c0.data_out_frame_29_7_N_1483_1 ;
    wire \c0.n19297 ;
    wire \c0.n3315 ;
    wire \c0.n19297_cascade_ ;
    wire \c0.data_out_frame_29_7_N_1483_2 ;
    wire \c0.data_in_frame_14_0 ;
    wire \c0.n18663_cascade_ ;
    wire \c0.n33397_cascade_ ;
    wire \c0.n33604 ;
    wire \c0.data_in_frame_9_0 ;
    wire \c0.data_in_frame_0_2 ;
    wire \c0.data_in_frame_0_3 ;
    wire \c0.data_in_frame_0_1 ;
    wire \c0.n28 ;
    wire \c0.n32 ;
    wire \c0.data_in_frame_6_3 ;
    wire \c0.data_in_frame_4_0 ;
    wire \c0.n18663 ;
    wire \c0.n33344_cascade_ ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.n10_adj_4770_cascade_ ;
    wire \c0.n18314 ;
    wire \c0.data_in_frame_6_2 ;
    wire \c0.data_in_frame_4_3 ;
    wire \c0.data_in_frame_2_0 ;
    wire \c0.n33692 ;
    wire \c0.rx.n6_cascade_ ;
    wire \c0.rx.n35949_cascade_ ;
    wire n4_adj_4807;
    wire n4_adj_4807_cascade_;
    wire n18031;
    wire \c0.data_in_frame_5_2 ;
    wire \c0.data_in_frame_14_3 ;
    wire \c0.n6_adj_4546 ;
    wire \c0.data_in_frame_15_2 ;
    wire \c0.n33321 ;
    wire \c0.data_in_frame_3_7 ;
    wire \c0.data_in_frame_15_6 ;
    wire \c0.data_in_frame_12_1 ;
    wire \c0.n33843 ;
    wire \c0.n31_adj_4740 ;
    wire \c0.data_in_frame_15_7 ;
    wire \c0.data_in_frame_13_6 ;
    wire \c0.n6_adj_4715 ;
    wire \c0.n31480_cascade_ ;
    wire \c0.n33422 ;
    wire \c0.data_in_frame_13_5 ;
    wire \c0.n33610 ;
    wire \c0.n35077 ;
    wire \c0.data_in_frame_13_0 ;
    wire \c0.n12_adj_4714 ;
    wire \c0.n33913_cascade_ ;
    wire \c0.n18881 ;
    wire \c0.n18847 ;
    wire \c0.n16010_cascade_ ;
    wire \c0.n31526 ;
    wire \c0.n33591 ;
    wire \c0.n32241_cascade_ ;
    wire \c0.n16010 ;
    wire \c0.n18805 ;
    wire \c0.n34012 ;
    wire \c0.n18438 ;
    wire \c0.n33629 ;
    wire \c0.data_in_frame_28_4 ;
    wire \c0.n12_adj_4748_cascade_ ;
    wire \c0.n33517 ;
    wire \c0.n33517_cascade_ ;
    wire \c0.n33441 ;
    wire \c0.n33768 ;
    wire \c0.data_in_frame_12_4 ;
    wire \c0.n33768_cascade_ ;
    wire \c0.n33417 ;
    wire \c0.n6023 ;
    wire \c0.n6023_cascade_ ;
    wire \c0.data_in_frame_17_0 ;
    wire \c0.n33458 ;
    wire \c0.n19108 ;
    wire \c0.n10_adj_4709 ;
    wire \c0.n33621_cascade_ ;
    wire \c0.data_in_frame_16_7 ;
    wire \c0.data_in_frame_19_3 ;
    wire \c0.n12_adj_4712 ;
    wire \c0.n8_adj_4711_cascade_ ;
    wire \c0.n19060 ;
    wire \c0.n18578_cascade_ ;
    wire \c0.n15_adj_4746_cascade_ ;
    wire \c0.n14_adj_4578 ;
    wire \c0.n32087_cascade_ ;
    wire \c0.data_in_frame_26_5 ;
    wire \c0.n33966 ;
    wire \c0.data_in_frame_16_3 ;
    wire \c0.n33526 ;
    wire \c0.data_in_frame_18_5 ;
    wire \c0.n31651 ;
    wire \c0.n18559_cascade_ ;
    wire \c0.n33972 ;
    wire \c0.n33653 ;
    wire \c0.n15_adj_4664_cascade_ ;
    wire \c0.n14_adj_4663 ;
    wire \c0.n33939 ;
    wire \c0.data_in_frame_20_7 ;
    wire \c0.data_in_frame_20_6 ;
    wire \c0.data_in_frame_23_2 ;
    wire \c0.n18559 ;
    wire \c0.n6404_cascade_ ;
    wire \c0.n32390 ;
    wire \c0.data_in_frame_16_6 ;
    wire \quad_counter0.n2017 ;
    wire \quad_counter0.n2084 ;
    wire \quad_counter0.n2081 ;
    wire \quad_counter0.n2014 ;
    wire \quad_counter0.n2015 ;
    wire \quad_counter0.n2082 ;
    wire \quad_counter0.n1919 ;
    wire \quad_counter0.n1986 ;
    wire \quad_counter0.n1946 ;
    wire \quad_counter0.n2018 ;
    wire \quad_counter0.n2085 ;
    wire \quad_counter0.n2018_cascade_ ;
    wire \quad_counter0.n2016 ;
    wire \quad_counter0.n2083 ;
    wire \quad_counter0.n2045 ;
    wire \quad_counter0.n8_adj_4380_cascade_ ;
    wire \quad_counter0.n7_adj_4381 ;
    wire \quad_counter0.n35542_cascade_ ;
    wire bfn_15_9_0_;
    wire \quad_counter0.n3419 ;
    wire \quad_counter0.n30425 ;
    wire \quad_counter0.n3418 ;
    wire \quad_counter0.n30426 ;
    wire \quad_counter0.n3417 ;
    wire \quad_counter0.n30427 ;
    wire \quad_counter0.n3416 ;
    wire \quad_counter0.n30428 ;
    wire \quad_counter0.n3415 ;
    wire \quad_counter0.n30429 ;
    wire \quad_counter0.n3414 ;
    wire \quad_counter0.n36139 ;
    wire \quad_counter0.n30430 ;
    wire \quad_counter0.n3413 ;
    wire \quad_counter0.n30431 ;
    wire \quad_counter0.n30432 ;
    wire \quad_counter0.n3412 ;
    wire \quad_counter0.n3511 ;
    wire bfn_15_10_0_;
    wire \quad_counter0.n3411 ;
    wire \quad_counter0.n3510 ;
    wire \quad_counter0.n30433 ;
    wire \quad_counter0.n3410 ;
    wire \quad_counter0.n3509 ;
    wire \quad_counter0.n30434 ;
    wire \quad_counter0.n3409 ;
    wire \quad_counter0.n30435 ;
    wire \quad_counter0.n3408 ;
    wire \quad_counter0.n30436 ;
    wire \quad_counter0.n3407 ;
    wire \quad_counter0.n3506 ;
    wire \quad_counter0.n30437 ;
    wire \quad_counter0.n3406 ;
    wire \quad_counter0.n3505 ;
    wire \quad_counter0.n30438 ;
    wire \quad_counter0.n3405 ;
    wire \quad_counter0.n30439 ;
    wire \quad_counter0.n30440 ;
    wire \quad_counter0.n3404 ;
    wire \quad_counter0.n3503 ;
    wire bfn_15_11_0_;
    wire \quad_counter0.n3403 ;
    wire \quad_counter0.n30441 ;
    wire \quad_counter0.n3402 ;
    wire \quad_counter0.n30442 ;
    wire \quad_counter0.n3401 ;
    wire \quad_counter0.n30443 ;
    wire \quad_counter0.n3400 ;
    wire \quad_counter0.n30444 ;
    wire \quad_counter0.n3399 ;
    wire \quad_counter0.n30445 ;
    wire \quad_counter0.n3398 ;
    wire \quad_counter0.n3431 ;
    wire \quad_counter0.n30446 ;
    wire \quad_counter0.n3497 ;
    wire \quad_counter0.n36150 ;
    wire \quad_counter0.n2639 ;
    wire r_Tx_Data_3;
    wire data_out_frame_12_0;
    wire data_out_frame_13_0;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.n4_adj_4646 ;
    wire r_Tx_Data_7;
    wire n36084_cascade_;
    wire n10_adj_4804;
    wire r_Tx_Data_0;
    wire data_out_frame_10_1;
    wire data_out_frame_11_1;
    wire \c0.n35833 ;
    wire n35835;
    wire data_out_frame_9_0;
    wire \c0.n11 ;
    wire \c0.n36200_cascade_ ;
    wire data_out_frame_6_2;
    wire \c0.n5_adj_4511 ;
    wire \c0.n36209 ;
    wire data_out_frame_8_1;
    wire \c0.n36212_cascade_ ;
    wire n36092;
    wire n36088;
    wire n35820;
    wire \c0.n17959 ;
    wire \c0.n30906 ;
    wire \c0.n5024 ;
    wire n35991_cascade_;
    wire \c0.n11_adj_4626 ;
    wire \c0.rx.n28401_cascade_ ;
    wire n28381_cascade_;
    wire n1;
    wire data_out_frame_7_6;
    wire n35992;
    wire \c0.rx.r_SM_Main_2_N_3681_2_cascade_ ;
    wire \c0.rx.r_Bit_Index_0 ;
    wire \c0.rx.n34091_cascade_ ;
    wire \c0.rx.r_Bit_Index_1 ;
    wire \c0.rx.n28401 ;
    wire \c0.rx.n29888 ;
    wire \c0.rx.n34091 ;
    wire \c0.rx.n3821 ;
    wire \c0.rx.n29888_cascade_ ;
    wire \c0.rx.r_Bit_Index_2 ;
    wire \c0.data_in_frame_5_7 ;
    wire r_Rx_Data;
    wire \c0.rx.n35769_cascade_ ;
    wire \c0.rx.r_SM_Main_2_N_3687_0 ;
    wire \c0.rx.n35738 ;
    wire \c0.data_in_frame_3_4 ;
    wire \c0.rx.n33223_cascade_ ;
    wire \c0.rx.n35950 ;
    wire \c0.data_in_frame_13_1 ;
    wire \c0.n33233_cascade_ ;
    wire \c0.n63_adj_4633 ;
    wire \c0.n35633 ;
    wire \c0.n27708 ;
    wire \c0.data_in_frame_15_3 ;
    wire \c0.n18373 ;
    wire \c0.data_in_frame_23_7 ;
    wire \c0.n33813 ;
    wire \c0.data_in_frame_13_7 ;
    wire \c0.n14_adj_4538 ;
    wire \c0.n34727_cascade_ ;
    wire \c0.n29_adj_4761 ;
    wire \c0.data_in_frame_28_3 ;
    wire \c0.n34566 ;
    wire \c0.n24_adj_4760 ;
    wire \c0.data_in_frame_28_1 ;
    wire \c0.n17531_cascade_ ;
    wire \c0.n17545 ;
    wire \c0.n18588 ;
    wire \c0.data_in_frame_20_2 ;
    wire \c0.data_in_frame_16_0 ;
    wire \c0.n33601 ;
    wire \c0.n33827 ;
    wire \c0.n18974 ;
    wire \c0.n18974_cascade_ ;
    wire \c0.data_in_frame_18_1 ;
    wire \c0.data_in_frame_20_3 ;
    wire \c0.n6_adj_4661 ;
    wire \c0.data_in_frame_12_2 ;
    wire \c0.data_in_frame_15_1 ;
    wire \c0.n32087 ;
    wire \c0.n33864_cascade_ ;
    wire \c0.n33979 ;
    wire \c0.data_in_frame_14_4 ;
    wire \c0.n20_adj_4627 ;
    wire \c0.data_in_frame_20_5 ;
    wire \c0.n32357 ;
    wire \c0.n32026_cascade_ ;
    wire \c0.n16_adj_4667 ;
    wire \c0.n31940 ;
    wire \c0.n24_adj_4671 ;
    wire \c0.n32026 ;
    wire \c0.data_in_frame_16_2 ;
    wire \c0.n32241 ;
    wire \c0.n33618 ;
    wire \c0.n33618_cascade_ ;
    wire \c0.n6462 ;
    wire \c0.n22_adj_4670 ;
    wire \c0.n33514 ;
    wire \c0.n18166 ;
    wire \c0.n31417 ;
    wire \c0.n33833 ;
    wire \c0.n18487 ;
    wire \c0.n33621 ;
    wire \c0.n17702 ;
    wire \c0.n17702_cascade_ ;
    wire bfn_16_6_0_;
    wire \quad_counter0.n2119 ;
    wire \quad_counter0.n30230 ;
    wire \quad_counter0.n2118 ;
    wire \quad_counter0.n30231 ;
    wire \quad_counter0.n2117 ;
    wire \quad_counter0.n30232 ;
    wire \quad_counter0.n2116 ;
    wire \quad_counter0.n30233 ;
    wire \quad_counter0.n2115 ;
    wire \quad_counter0.n30234 ;
    wire \quad_counter0.n2114 ;
    wire \quad_counter0.n30235 ;
    wire \quad_counter0.n2113 ;
    wire \quad_counter0.n30236 ;
    wire \quad_counter0.n30237 ;
    wire \quad_counter0.n2112 ;
    wire bfn_16_7_0_;
    wire \quad_counter0.n2111 ;
    wire \quad_counter0.n30238 ;
    wire \quad_counter0.n2144 ;
    wire \quad_counter0.n36157 ;
    wire \quad_counter0.n10_adj_4389_cascade_ ;
    wire \quad_counter0.n14_adj_4418 ;
    wire \quad_counter0.n15_cascade_ ;
    wire \quad_counter0.n3512 ;
    wire \quad_counter0.n3513 ;
    wire \quad_counter0.n3507 ;
    wire \quad_counter0.n3500 ;
    wire \quad_counter0.n35976 ;
    wire \quad_counter0.n35977_cascade_ ;
    wire \quad_counter0.n33_adj_4346 ;
    wire \quad_counter0.n34205 ;
    wire \quad_counter0.n3508 ;
    wire \quad_counter0.n3501 ;
    wire \quad_counter0.n3504 ;
    wire \quad_counter0.n3499 ;
    wire \quad_counter0.n3502 ;
    wire \quad_counter0.n3498 ;
    wire \quad_counter0.n31_cascade_ ;
    wire \quad_counter0.n28_adj_4342 ;
    wire \quad_counter0.n34 ;
    wire \quad_counter0.n35978 ;
    wire bfn_16_12_0_;
    wire \quad_counter0.n3519 ;
    wire \quad_counter0.n30453 ;
    wire \quad_counter0.n3518 ;
    wire \quad_counter0.n30454 ;
    wire \quad_counter0.n12903 ;
    wire \quad_counter0.n3517 ;
    wire \quad_counter0.n9 ;
    wire \quad_counter0.n30455 ;
    wire \quad_counter0.n3516 ;
    wire \quad_counter0.n30456 ;
    wire \quad_counter0.n12904 ;
    wire \quad_counter0.n3515 ;
    wire \quad_counter0.n8_adj_4375 ;
    wire \quad_counter0.n30457 ;
    wire \quad_counter0.n12901 ;
    wire \quad_counter0.n3514 ;
    wire \quad_counter0.n30458 ;
    wire \quad_counter0.n10_adj_4347 ;
    wire \quad_counter0.n11 ;
    wire \quad_counter0.n28339_cascade_ ;
    wire \quad_counter0.n10_adj_4400 ;
    wire \quad_counter0.n10_adj_4399_cascade_ ;
    wire \quad_counter0.n16_adj_4401 ;
    wire \c0.n6_adj_4647_cascade_ ;
    wire \c0.n28313 ;
    wire data_out_frame_9_2;
    wire data_out_frame_8_2;
    wire \c0.n36206 ;
    wire n10;
    wire n10_adj_4806;
    wire \c0.n35963 ;
    wire data_out_frame_11_2;
    wire data_out_frame_10_2;
    wire \c0.n36203 ;
    wire data_out_frame_8_0;
    wire data_out_frame_9_7;
    wire \c0.n36194_cascade_ ;
    wire \c0.n11_adj_4655 ;
    wire n36094;
    wire \c0.n5 ;
    wire data_out_frame_7_3;
    wire data_out_frame_6_3;
    wire data_out_frame_12_6;
    wire \c0.n7_adj_4499 ;
    wire n35818;
    wire \c0.data_in_frame_4_1 ;
    wire \c0.data_in_frame_2_1 ;
    wire data_out_frame_13_6;
    wire \c0.rx.n19345_cascade_ ;
    wire \c0.rx.r_SM_Main_2_N_3681_2 ;
    wire \c0.rx.n17939 ;
    wire \c0.FRAME_MATCHER_rx_data_ready_prev ;
    wire rx_data_ready;
    wire r_Clock_Count_0;
    wire n226;
    wire bfn_16_21_0_;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n30061 ;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.n30062 ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.n30063 ;
    wire \c0.rx.n30064 ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.n30065 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.n30066 ;
    wire \c0.rx.n30067 ;
    wire \c0.rx.r_Clock_Count_7 ;
    wire n19327;
    wire n19940;
    wire \c0.n33241 ;
    wire \c0.data_in_frame_9_3 ;
    wire \c0.data_in_frame_6_0 ;
    wire data_in_frame_1_2;
    wire n36096;
    wire n10_adj_4820;
    wire \c0.n33506_cascade_ ;
    wire \c0.n33889 ;
    wire \c0.n12_adj_4710_cascade_ ;
    wire \c0.n32346 ;
    wire \c0.n18784_cascade_ ;
    wire \c0.n10_adj_4749 ;
    wire \c0.data_in_frame_23_6 ;
    wire \c0.n33726 ;
    wire \c0.n33329 ;
    wire \c0.n33726_cascade_ ;
    wire \c0.n15_adj_4747 ;
    wire \c0.n33532 ;
    wire \c0.data_in_frame_19_5 ;
    wire \c0.data_in_frame_23_3 ;
    wire \c0.n18784 ;
    wire \c0.data_in_frame_20_4 ;
    wire \c0.data_in_frame_22_5 ;
    wire \c0.n6_adj_4675 ;
    wire \c0.data_in_frame_29_6 ;
    wire \c0.data_in_frame_21_0 ;
    wire \c0.data_in_frame_29_0 ;
    wire \c0.n35181 ;
    wire \c0.data_in_frame_22_1 ;
    wire \c0.n33598 ;
    wire \c0.n33374_cascade_ ;
    wire \c0.data_in_frame_28_6 ;
    wire \c0.n38_adj_4701 ;
    wire \c0.n40_adj_4700 ;
    wire \c0.n39_adj_4702 ;
    wire \c0.n10_adj_4669 ;
    wire \c0.n35307 ;
    wire \c0.n16120_cascade_ ;
    wire \c0.data_in_frame_19_6 ;
    wire \c0.n6227 ;
    wire \c0.n31444 ;
    wire \c0.n41_adj_4704 ;
    wire \c0.n42_adj_4703 ;
    wire \c0.n33490_cascade_ ;
    wire \c0.n46 ;
    wire \c0.n25_cascade_ ;
    wire \c0.n31_cascade_ ;
    wire \c0.n18861 ;
    wire \c0.n33913 ;
    wire \c0.n33969 ;
    wire \c0.data_in_frame_16_5 ;
    wire \c0.n18228 ;
    wire \c0.n33957 ;
    wire \quad_counter1.n28257_cascade_ ;
    wire \quad_counter1.n10_adj_4472_cascade_ ;
    wire \quad_counter1.B_delayed ;
    wire \quad_counter1.A_delayed ;
    wire A_filtered_adj_4809;
    wire B_filtered_adj_4810;
    wire \quad_counter0.millisecond_counter_0 ;
    wire bfn_17_8_0_;
    wire \quad_counter0.millisecond_counter_1 ;
    wire \quad_counter0.n30140 ;
    wire \quad_counter0.millisecond_counter_2 ;
    wire \quad_counter0.n30141 ;
    wire \quad_counter0.millisecond_counter_3 ;
    wire \quad_counter0.n30142 ;
    wire \quad_counter0.millisecond_counter_4 ;
    wire \quad_counter0.n30143 ;
    wire \quad_counter0.millisecond_counter_5 ;
    wire \quad_counter0.n30144 ;
    wire \quad_counter0.millisecond_counter_6 ;
    wire \quad_counter0.n30145 ;
    wire \quad_counter0.millisecond_counter_7 ;
    wire \quad_counter0.n30146 ;
    wire \quad_counter0.n30147 ;
    wire \quad_counter0.millisecond_counter_8 ;
    wire bfn_17_9_0_;
    wire \quad_counter0.millisecond_counter_9 ;
    wire \quad_counter0.n30148 ;
    wire \quad_counter0.millisecond_counter_10 ;
    wire \quad_counter0.n30149 ;
    wire \quad_counter0.millisecond_counter_11 ;
    wire \quad_counter0.n30150 ;
    wire \quad_counter0.millisecond_counter_12 ;
    wire \quad_counter0.n30151 ;
    wire \quad_counter0.millisecond_counter_13 ;
    wire \quad_counter0.n30152 ;
    wire \quad_counter0.millisecond_counter_14 ;
    wire \quad_counter0.n30153 ;
    wire \quad_counter0.millisecond_counter_15 ;
    wire \quad_counter0.n30154 ;
    wire \quad_counter0.n30155 ;
    wire \quad_counter0.millisecond_counter_16 ;
    wire bfn_17_10_0_;
    wire \quad_counter0.millisecond_counter_17 ;
    wire \quad_counter0.n30156 ;
    wire \quad_counter0.n30157 ;
    wire \quad_counter0.n30158 ;
    wire \quad_counter0.n30159 ;
    wire \quad_counter0.n30160 ;
    wire \quad_counter0.millisecond_counter_22 ;
    wire \quad_counter0.n30161 ;
    wire \quad_counter0.millisecond_counter_23 ;
    wire \quad_counter0.n30162 ;
    wire \quad_counter0.n30163 ;
    wire \quad_counter0.millisecond_counter_24 ;
    wire bfn_17_11_0_;
    wire \quad_counter0.millisecond_counter_25 ;
    wire \quad_counter0.n30164 ;
    wire \quad_counter0.millisecond_counter_26 ;
    wire \quad_counter0.n30165 ;
    wire \quad_counter0.millisecond_counter_27 ;
    wire \quad_counter0.n30166 ;
    wire \quad_counter0.millisecond_counter_28 ;
    wire \quad_counter0.n30167 ;
    wire \quad_counter0.millisecond_counter_29 ;
    wire \quad_counter0.n30168 ;
    wire \quad_counter0.millisecond_counter_30 ;
    wire \quad_counter0.n30169 ;
    wire \quad_counter0.n30170 ;
    wire \quad_counter0.millisecond_counter_31 ;
    wire n34523;
    wire count_prev_0;
    wire \quad_counter0.n2619 ;
    wire bfn_17_13_0_;
    wire \quad_counter0.n2618 ;
    wire \quad_counter0.n30272 ;
    wire \quad_counter0.n2617 ;
    wire \quad_counter0.n30273 ;
    wire \quad_counter0.n2616 ;
    wire \quad_counter0.n30274 ;
    wire \quad_counter0.n2615 ;
    wire \quad_counter0.n30275 ;
    wire \quad_counter0.n2614 ;
    wire \quad_counter0.n30276 ;
    wire \quad_counter0.n2613 ;
    wire \quad_counter0.n30277 ;
    wire \quad_counter0.n2612 ;
    wire \quad_counter0.n30278 ;
    wire \quad_counter0.n30279 ;
    wire \quad_counter0.n2611 ;
    wire bfn_17_14_0_;
    wire \quad_counter0.n2610 ;
    wire \quad_counter0.n30280 ;
    wire \quad_counter0.n2609 ;
    wire \quad_counter0.n30281 ;
    wire \quad_counter0.n2608 ;
    wire \quad_counter0.n30282 ;
    wire \quad_counter0.n2607 ;
    wire \quad_counter0.n30283 ;
    wire \quad_counter0.n30284 ;
    wire \quad_counter0.n2606 ;
    wire data_out_frame_9_3;
    wire \c0.n36161_cascade_ ;
    wire \c0.n36164_cascade_ ;
    wire n36082;
    wire \c0.n5_adj_4515 ;
    wire \c0.n6_adj_4514 ;
    wire \c0.n35836_cascade_ ;
    wire n35838;
    wire data_out_frame_10_3;
    wire data_out_frame_8_3;
    wire data_out_frame_12_7;
    wire \c0.n36021 ;
    wire data_out_frame_11_0;
    wire data_out_frame_10_0;
    wire \c0.n36197 ;
    wire data_out_frame_13_7;
    wire \c0.n36191 ;
    wire data_out_frame_10_6;
    wire data_out_frame_11_6;
    wire data_out_frame_9_6;
    wire \c0.n36185_cascade_ ;
    wire \c0.n36188 ;
    wire data_out_frame_9_1;
    wire \c0.n33500 ;
    wire \c0.n18627 ;
    wire \c0.n18479 ;
    wire data_out_frame_11_7;
    wire data_out_frame_5_5;
    wire data_out_frame_7_2;
    wire \c0.data_in_frame_6_4 ;
    wire data_out_frame_6_5;
    wire data_out_frame_7_5;
    wire \c0.n36086 ;
    wire \c0.n5_adj_4619_cascade_ ;
    wire data_out_frame_6_6;
    wire \c0.n36012 ;
    wire \c0.n5_adj_4624 ;
    wire \c0.data_in_frame_0_7 ;
    wire data_out_frame_8_6;
    wire data_out_frame_5_6;
    wire bfn_17_22_0_;
    wire \quad_counter0.count_direction ;
    wire \quad_counter0.n30108 ;
    wire \quad_counter0.n30109 ;
    wire \quad_counter0.n30110 ;
    wire \quad_counter0.n30111 ;
    wire \quad_counter0.n30112 ;
    wire \quad_counter0.n30113 ;
    wire \quad_counter0.n30114 ;
    wire \quad_counter0.n30115 ;
    wire bfn_17_23_0_;
    wire \quad_counter0.n30116 ;
    wire \quad_counter0.n30117 ;
    wire \quad_counter0.n30118 ;
    wire \quad_counter0.n30119 ;
    wire \quad_counter0.n30120 ;
    wire \quad_counter0.n30121 ;
    wire \quad_counter0.n30122 ;
    wire \quad_counter0.n30123 ;
    wire bfn_17_24_0_;
    wire \quad_counter0.n30124 ;
    wire \quad_counter0.n30125 ;
    wire \quad_counter0.n30126 ;
    wire n2326;
    wire \quad_counter0.n30127 ;
    wire \quad_counter0.n30128 ;
    wire encoder0_position_21;
    wire n2324;
    wire \quad_counter0.n30129 ;
    wire n2323;
    wire \quad_counter0.n30130 ;
    wire \quad_counter0.n30131 ;
    wire bfn_17_25_0_;
    wire \quad_counter0.n30132 ;
    wire \quad_counter0.n30133 ;
    wire \quad_counter0.n30134 ;
    wire n2318;
    wire \quad_counter0.n30135 ;
    wire \quad_counter0.n30136 ;
    wire n2316;
    wire \quad_counter0.n30137 ;
    wire \quad_counter0.n30138 ;
    wire \quad_counter0.n30139 ;
    wire \quad_counter0.n2300 ;
    wire bfn_17_26_0_;
    wire \c0.n12_adj_4759 ;
    wire \c0.n34841 ;
    wire \c0.n6_adj_4666 ;
    wire \c0.n32366 ;
    wire \c0.data_in_frame_21_7 ;
    wire \c0.data_in_frame_21_6 ;
    wire \c0.data_in_frame_24_1 ;
    wire \c0.n33662 ;
    wire \c0.n36530_cascade_ ;
    wire \c0.n32431_cascade_ ;
    wire \c0.n32431 ;
    wire \c0.data_in_frame_29_4 ;
    wire \c0.data_in_frame_17_3 ;
    wire \c0.n18011 ;
    wire \c0.data_in_frame_23_4 ;
    wire \c0.data_in_frame_16_4 ;
    wire \c0.data_in_frame_18_4 ;
    wire \c0.n18415 ;
    wire \c0.n29 ;
    wire \quad_counter1.n2936_cascade_ ;
    wire \quad_counter1.n28263 ;
    wire \quad_counter1.n10_adj_4458_cascade_ ;
    wire \quad_counter1.n20 ;
    wire \quad_counter1.n13_cascade_ ;
    wire \quad_counter1.n22 ;
    wire bfn_18_3_0_;
    wire \quad_counter1.n30580 ;
    wire \quad_counter1.n30581 ;
    wire \quad_counter1.n30582 ;
    wire \quad_counter1.n30583 ;
    wire \quad_counter1.n30584 ;
    wire \quad_counter1.n36159 ;
    wire \quad_counter1.n30585 ;
    wire \quad_counter1.n30586 ;
    wire \quad_counter1.n30587 ;
    wire bfn_18_4_0_;
    wire \quad_counter1.n30588 ;
    wire \quad_counter1.n30589 ;
    wire \quad_counter1.n30590 ;
    wire \quad_counter1.n30591 ;
    wire \quad_counter1.n30592 ;
    wire \quad_counter1.n30593 ;
    wire \quad_counter1.n30594 ;
    wire \quad_counter1.n30595 ;
    wire bfn_18_5_0_;
    wire \quad_counter1.n2936 ;
    wire \quad_counter1.n30596 ;
    wire \quad_counter1.n18_adj_4459 ;
    wire \quad_counter1.n16_adj_4473 ;
    wire \quad_counter1.n22_adj_4474 ;
    wire \quad_counter1.n24_adj_4476_cascade_ ;
    wire \quad_counter1.n20_adj_4475 ;
    wire \quad_counter1.n3035_cascade_ ;
    wire \quad_counter0.n28365 ;
    wire \quad_counter0.n10_adj_4382_cascade_ ;
    wire \quad_counter0.n7_adj_4383_cascade_ ;
    wire \quad_counter0.n2243_cascade_ ;
    wire \quad_counter0.millisecond_counter_21 ;
    wire bfn_18_9_0_;
    wire \quad_counter0.n2219 ;
    wire \quad_counter0.n30239 ;
    wire \quad_counter0.n2218 ;
    wire \quad_counter0.n30240 ;
    wire \quad_counter0.n2217 ;
    wire \quad_counter0.n30241 ;
    wire \quad_counter0.n2216 ;
    wire \quad_counter0.n30242 ;
    wire \quad_counter0.n2215 ;
    wire \quad_counter0.n30243 ;
    wire \quad_counter0.n2214 ;
    wire \quad_counter0.n36155 ;
    wire \quad_counter0.n30244 ;
    wire \quad_counter0.n2213 ;
    wire \quad_counter0.n30245 ;
    wire \quad_counter0.n30246 ;
    wire \quad_counter0.n2212 ;
    wire bfn_18_10_0_;
    wire \quad_counter0.n2211 ;
    wire \quad_counter0.n30247 ;
    wire \quad_counter0.n2210 ;
    wire \quad_counter0.n2243 ;
    wire \quad_counter0.n30248 ;
    wire \quad_counter0.n7_adj_4393 ;
    wire \quad_counter0.n2342_adj_4384_cascade_ ;
    wire \quad_counter0.n28361 ;
    wire \quad_counter0.n8_adj_4390 ;
    wire \quad_counter0.millisecond_counter_20 ;
    wire bfn_18_11_0_;
    wire \quad_counter0.n2319_adj_4385 ;
    wire \quad_counter0.n30249 ;
    wire \quad_counter0.n2318_adj_4386 ;
    wire \quad_counter0.n30250 ;
    wire \quad_counter0.n2317_adj_4387 ;
    wire \quad_counter0.n30251 ;
    wire \quad_counter0.n2316_adj_4391 ;
    wire \quad_counter0.n30252 ;
    wire \quad_counter0.n2315_adj_4392 ;
    wire \quad_counter0.n30253 ;
    wire \quad_counter0.n2314_adj_4388 ;
    wire \quad_counter0.n36154 ;
    wire \quad_counter0.n30254 ;
    wire \quad_counter0.n2313 ;
    wire \quad_counter0.n30255 ;
    wire \quad_counter0.n30256 ;
    wire \quad_counter0.n2312 ;
    wire bfn_18_12_0_;
    wire \quad_counter0.n2311 ;
    wire \quad_counter0.n30257 ;
    wire \quad_counter0.n2310 ;
    wire \quad_counter0.n30258 ;
    wire \quad_counter0.n2309 ;
    wire \quad_counter0.n2342_adj_4384 ;
    wire \quad_counter0.n30259 ;
    wire \quad_counter0.millisecond_counter_19 ;
    wire bfn_18_13_0_;
    wire \quad_counter0.n2419 ;
    wire \quad_counter0.n30260 ;
    wire \quad_counter0.n2418 ;
    wire \quad_counter0.n30261 ;
    wire \quad_counter0.n30262 ;
    wire \quad_counter0.n2416 ;
    wire \quad_counter0.n30263 ;
    wire \quad_counter0.n2415 ;
    wire \quad_counter0.n30264 ;
    wire \quad_counter0.n36153 ;
    wire \quad_counter0.n30265 ;
    wire \quad_counter0.n2413 ;
    wire \quad_counter0.n30266 ;
    wire \quad_counter0.n30267 ;
    wire \quad_counter0.n2412 ;
    wire bfn_18_14_0_;
    wire \quad_counter0.n2411 ;
    wire \quad_counter0.n30268 ;
    wire \quad_counter0.n2410 ;
    wire \quad_counter0.n30269 ;
    wire \quad_counter0.n2409 ;
    wire \quad_counter0.n30270 ;
    wire \quad_counter0.n2408 ;
    wire \quad_counter0.n2441 ;
    wire \quad_counter0.n30271 ;
    wire \quad_counter0.millisecond_counter_18 ;
    wire \quad_counter0.n2519 ;
    wire \quad_counter0.n2513 ;
    wire \quad_counter0.n2512 ;
    wire \quad_counter0.n2511 ;
    wire \quad_counter0.n2509 ;
    wire \quad_counter0.n2508 ;
    wire \quad_counter0.n2507 ;
    wire \quad_counter0.n14 ;
    wire \quad_counter0.n2540 ;
    wire \quad_counter0.n2540_cascade_ ;
    wire \quad_counter0.n36151 ;
    wire \quad_counter0.n2517 ;
    wire \quad_counter0.n2518 ;
    wire \quad_counter0.n28345 ;
    wire \quad_counter0.n2514 ;
    wire \quad_counter0.n2516 ;
    wire \quad_counter0.n2515 ;
    wire \quad_counter0.n10_adj_4397_cascade_ ;
    wire \quad_counter0.n2510 ;
    wire \quad_counter0.n9_adj_4398 ;
    wire bfn_18_16_0_;
    wire \quad_counter1.count_direction ;
    wire n2279;
    wire \quad_counter1.n30076 ;
    wire \quad_counter1.n30077 ;
    wire \quad_counter1.n30078 ;
    wire \quad_counter1.n30079 ;
    wire \quad_counter1.n30080 ;
    wire \quad_counter1.n30081 ;
    wire \quad_counter1.n30082 ;
    wire \quad_counter1.n30083 ;
    wire n2272;
    wire bfn_18_17_0_;
    wire \quad_counter1.n30084 ;
    wire \quad_counter1.n30085 ;
    wire n2269;
    wire \quad_counter1.n30086 ;
    wire \quad_counter1.n30087 ;
    wire \quad_counter1.n30088 ;
    wire \quad_counter1.n30089 ;
    wire \quad_counter1.n30090 ;
    wire \quad_counter1.n30091 ;
    wire bfn_18_18_0_;
    wire \quad_counter1.n30092 ;
    wire \quad_counter1.n30093 ;
    wire \quad_counter1.n30094 ;
    wire n2260;
    wire \quad_counter1.n30095 ;
    wire \quad_counter1.n30096 ;
    wire \quad_counter1.n30097 ;
    wire \quad_counter1.n30098 ;
    wire \quad_counter1.n30099 ;
    wire n2256;
    wire bfn_18_19_0_;
    wire \quad_counter1.n30100 ;
    wire \quad_counter1.n30101 ;
    wire n2253;
    wire \quad_counter1.n30102 ;
    wire \quad_counter1.n30103 ;
    wire \quad_counter1.n30104 ;
    wire \quad_counter1.n30105 ;
    wire \quad_counter1.n30106 ;
    wire \quad_counter1.n30107 ;
    wire \quad_counter1.n2230 ;
    wire bfn_18_20_0_;
    wire data_in_frame_1_6;
    wire n2252;
    wire n2257;
    wire data_out_frame_8_7;
    wire data_in_frame_1_3;
    wire n2251;
    wire \c0.data_out_frame_0_4 ;
    wire \c0.n36173_cascade_ ;
    wire \c0.n35814_cascade_ ;
    wire r_SM_Main_1;
    wire \c0.rx.r_SM_Main_0 ;
    wire data_out_frame_7_4;
    wire \c0.n5_adj_4707 ;
    wire n2345;
    wire n2342;
    wire n2339;
    wire \c0.data_in_frame_5_3 ;
    wire n2262;
    wire n2255;
    wire data_out_frame_11_4;
    wire data_out_frame_10_4;
    wire \c0.n35813 ;
    wire \c0.n35964 ;
    wire n2325;
    wire \c0.n33407 ;
    wire n2331;
    wire \c0.n27862 ;
    wire \c0.n18084 ;
    wire \c0.data_in_frame_25_7 ;
    wire \c0.n33_adj_4764 ;
    wire \c0.n28_adj_4762_cascade_ ;
    wire n2249;
    wire \c0.n35314 ;
    wire \c0.n25_adj_4758 ;
    wire \c0.n31_adj_4763 ;
    wire \c0.data_in_frame_22_7 ;
    wire \c0.n31374 ;
    wire \c0.n33864 ;
    wire \c0.n18961_cascade_ ;
    wire \c0.n14_adj_4668 ;
    wire \c0.n33665 ;
    wire \c0.n32263 ;
    wire \c0.n32263_cascade_ ;
    wire \c0.n33576 ;
    wire \c0.data_in_frame_19_2 ;
    wire \c0.n6215 ;
    wire \c0.n33576_cascade_ ;
    wire \c0.n33577_cascade_ ;
    wire \c0.n33638 ;
    wire \c0.n14_adj_4757 ;
    wire \c0.data_in_frame_25_5 ;
    wire \c0.n30_adj_4706 ;
    wire \c0.n33632 ;
    wire \c0.n18405 ;
    wire \c0.data_in_frame_25_6 ;
    wire \c0.n13 ;
    wire \c0.n33994 ;
    wire \c0.n32294_cascade_ ;
    wire \c0.n37 ;
    wire \c0.n18961 ;
    wire \c0.data_in_frame_23_1 ;
    wire \c0.n33577 ;
    wire \c0.data_in_frame_23_5 ;
    wire \c0.n8_adj_4622 ;
    wire \c0.n7_adj_4662 ;
    wire \c0.n32316 ;
    wire \c0.n32316_cascade_ ;
    wire \c0.n31451 ;
    wire \c0.n21_adj_4659 ;
    wire \c0.n19_adj_4658_cascade_ ;
    wire \c0.n20_adj_4656 ;
    wire \c0.n5_adj_4660_cascade_ ;
    wire \c0.n16118 ;
    wire \c0.n33792 ;
    wire \c0.data_in_frame_24_3 ;
    wire \c0.n34006 ;
    wire \c0.data_in_frame_28_5 ;
    wire \c0.n10_adj_4755 ;
    wire \c0.data_in_frame_22_0 ;
    wire \c0.n35142 ;
    wire \c0.n35787 ;
    wire \c0.data_in_frame_26_1 ;
    wire \c0.n33991 ;
    wire \c0.n33858 ;
    wire \c0.n10_adj_4673_cascade_ ;
    wire \c0.n32310 ;
    wire \quad_counter1.n2919 ;
    wire bfn_19_2_0_;
    wire \quad_counter1.n2918 ;
    wire \quad_counter1.n30564 ;
    wire \quad_counter1.n2917 ;
    wire \quad_counter1.n30565 ;
    wire \quad_counter1.n2916 ;
    wire \quad_counter1.n30566 ;
    wire \quad_counter1.n2915 ;
    wire \quad_counter1.n30567 ;
    wire \quad_counter1.n2914 ;
    wire \quad_counter1.n30568 ;
    wire \quad_counter1.n2913 ;
    wire \quad_counter1.n30569 ;
    wire \quad_counter1.n2912 ;
    wire \quad_counter1.n30570 ;
    wire \quad_counter1.n30571 ;
    wire \quad_counter1.n2911 ;
    wire bfn_19_3_0_;
    wire \quad_counter1.n2910 ;
    wire \quad_counter1.n30572 ;
    wire \quad_counter1.n2909 ;
    wire \quad_counter1.n30573 ;
    wire \quad_counter1.n2908 ;
    wire \quad_counter1.n30574 ;
    wire \quad_counter1.n2907 ;
    wire \quad_counter1.n30575 ;
    wire \quad_counter1.n2906 ;
    wire \quad_counter1.n30576 ;
    wire \quad_counter1.n2905 ;
    wire \quad_counter1.n30577 ;
    wire \quad_counter1.n2904 ;
    wire \quad_counter1.n30578 ;
    wire \quad_counter1.n30579 ;
    wire bfn_19_4_0_;
    wire \quad_counter1.n2903 ;
    wire bfn_19_5_0_;
    wire \quad_counter1.n3019 ;
    wire \quad_counter1.n30597 ;
    wire \quad_counter1.n3018 ;
    wire \quad_counter1.n30598 ;
    wire \quad_counter1.n3017 ;
    wire \quad_counter1.n30599 ;
    wire \quad_counter1.n3016 ;
    wire \quad_counter1.n30600 ;
    wire \quad_counter1.n3015 ;
    wire \quad_counter1.n30601 ;
    wire \quad_counter1.n3014 ;
    wire \quad_counter1.n36156 ;
    wire \quad_counter1.n30602 ;
    wire \quad_counter1.n3013 ;
    wire \quad_counter1.n30603 ;
    wire \quad_counter1.n30604 ;
    wire \quad_counter1.n3012 ;
    wire bfn_19_6_0_;
    wire \quad_counter1.n3011 ;
    wire \quad_counter1.n30605 ;
    wire \quad_counter1.n3010 ;
    wire \quad_counter1.n30606 ;
    wire \quad_counter1.n3009 ;
    wire \quad_counter1.n30607 ;
    wire \quad_counter1.n3008 ;
    wire \quad_counter1.n30608 ;
    wire \quad_counter1.n3007 ;
    wire \quad_counter1.n30609 ;
    wire \quad_counter1.n3006 ;
    wire \quad_counter1.n30610 ;
    wire \quad_counter1.n3005 ;
    wire \quad_counter1.n30611 ;
    wire \quad_counter1.n30612 ;
    wire \quad_counter1.n3004 ;
    wire bfn_19_7_0_;
    wire \quad_counter1.n3003 ;
    wire \quad_counter1.n30613 ;
    wire \quad_counter1.n3002 ;
    wire \quad_counter1.n3035 ;
    wire \quad_counter1.n30614 ;
    wire \quad_counter1.n18_adj_4479_cascade_ ;
    wire \quad_counter1.n24_adj_4480 ;
    wire \quad_counter1.n19_adj_4485 ;
    wire \quad_counter1.n26_adj_4484_cascade_ ;
    wire bfn_19_11_0_;
    wire \quad_counter1.n30634 ;
    wire \quad_counter1.n30635 ;
    wire \quad_counter1.n30636 ;
    wire \quad_counter1.n30637 ;
    wire \quad_counter1.n30638 ;
    wire \quad_counter1.n30639 ;
    wire \quad_counter1.n30640 ;
    wire \quad_counter1.n30641 ;
    wire bfn_19_12_0_;
    wire \quad_counter1.n30642 ;
    wire \quad_counter1.n30643 ;
    wire \quad_counter1.n30644 ;
    wire \quad_counter1.n30645 ;
    wire \quad_counter1.n30646 ;
    wire \quad_counter1.n30647 ;
    wire \quad_counter1.n30648 ;
    wire \quad_counter1.n30649 ;
    wire bfn_19_13_0_;
    wire \quad_counter1.n30650 ;
    wire \quad_counter1.n30651 ;
    wire \quad_counter1.n30652 ;
    wire \quad_counter1.n30653 ;
    wire \quad_counter1.n36148 ;
    wire \quad_counter1.n24_adj_4487 ;
    wire \quad_counter1.n16_adj_4486 ;
    wire \quad_counter1.n28_adj_4488 ;
    wire \quad_counter1.n3233 ;
    wire n2278;
    wire data_out_frame_12_3;
    wire \c0.n11_adj_4517 ;
    wire n2264;
    wire n2276;
    wire \c0.n11_adj_4507 ;
    wire data_out_frame_12_1;
    wire data_out_frame_11_5;
    wire \c0.n36179_cascade_ ;
    wire data_out_frame_9_5;
    wire \c0.n36182_cascade_ ;
    wire n36098_cascade_;
    wire n2270;
    wire n2268;
    wire n2266;
    wire data_out_frame_8_5;
    wire \c0.n18357_cascade_ ;
    wire data_out_frame_10_7;
    wire n2263;
    wire n2265;
    wire n2258;
    wire \c0.n18689_cascade_ ;
    wire \c0.n38_adj_4568_cascade_ ;
    wire n2250;
    wire \c0.n43_adj_4569 ;
    wire n2254;
    wire \c0.data_in_frame_21_5 ;
    wire \c0.data_in_frame_5_1 ;
    wire encoder1_position_23;
    wire \c0.n33400 ;
    wire n2261;
    wire encoder1_position_25;
    wire encoder1_position_15;
    wire \c0.n11_adj_4576 ;
    wire data_out_frame_12_4;
    wire data_out_frame_5_3;
    wire data_in_frame_1_1;
    wire data_out_frame_5_4;
    wire encoder1_position_24;
    wire data_out_frame_12_5;
    wire \c0.n11_adj_4621 ;
    wire data_out_frame_13_5;
    wire data_out_frame_6_4;
    wire n2344;
    wire data_out_frame_13_4;
    wire n2327;
    wire n2314;
    wire n2338;
    wire \c0.n35140 ;
    wire \c0.n12_adj_4536 ;
    wire \c0.data_in_frame_5_4 ;
    wire n2332;
    wire \c0.n12_adj_4526 ;
    wire \c0.data_in_frame_13_4 ;
    wire n2330;
    wire \c0.data_in_frame_24_2 ;
    wire n2335;
    wire n2337;
    wire data_out_frame_8_4;
    wire \c0.n35812 ;
    wire data_out_frame_9_4;
    wire \c0.n18568 ;
    wire \c0.n35416 ;
    wire n2315;
    wire \c0.data_in_frame_27_7 ;
    wire \c0.data_in_frame_25_4 ;
    wire \c0.n33594 ;
    wire \c0.data_in_frame_24_4 ;
    wire \c0.n34009 ;
    wire \c0.n34009_cascade_ ;
    wire \c0.n31355 ;
    wire \c0.data_in_frame_27_0 ;
    wire \c0.data_in_frame_26_6 ;
    wire \c0.n33374 ;
    wire \c0.data_in_frame_26_4 ;
    wire \c0.data_in_frame_22_2 ;
    wire \c0.n33849 ;
    wire \c0.n18193 ;
    wire \c0.n33775 ;
    wire \c0.n33350 ;
    wire \c0.n32339 ;
    wire \c0.n8_adj_4540 ;
    wire \c0.n18596 ;
    wire \c0.n16120 ;
    wire \c0.n6_adj_4756 ;
    wire \c0.data_in_frame_27_2 ;
    wire \c0.n31784 ;
    wire \c0.n17_adj_4753 ;
    wire \c0.n4_adj_4751_cascade_ ;
    wire \c0.n20_adj_4754 ;
    wire \c0.data_in_frame_29_7 ;
    wire \c0.data_in_frame_27_6 ;
    wire \c0.n33463 ;
    wire \c0.n35250 ;
    wire \c0.data_in_frame_26_0 ;
    wire \c0.n33846 ;
    wire \c0.n33490 ;
    wire \c0.n33816 ;
    wire \c0.data_in_frame_28_7 ;
    wire \c0.n33976 ;
    wire \c0.n16_adj_4750_cascade_ ;
    wire \c0.n18_adj_4752 ;
    wire \c0.data_in_frame_27_4 ;
    wire \quad_counter1.n36131 ;
    wire \quad_counter1.n19_cascade_ ;
    wire \quad_counter1.n2837 ;
    wire \quad_counter1.n28267_cascade_ ;
    wire \quad_counter1.n10_adj_4455_cascade_ ;
    wire \quad_counter1.n12_adj_4456 ;
    wire \quad_counter1.n2819 ;
    wire bfn_20_4_0_;
    wire \quad_counter1.n2818 ;
    wire \quad_counter1.n30549 ;
    wire \quad_counter1.n2817 ;
    wire \quad_counter1.n30550 ;
    wire \quad_counter1.n2816 ;
    wire \quad_counter1.n30551 ;
    wire \quad_counter1.n2815 ;
    wire \quad_counter1.n30552 ;
    wire \quad_counter1.n2814 ;
    wire \quad_counter1.n30553 ;
    wire \quad_counter1.n30554 ;
    wire \quad_counter1.n2812 ;
    wire \quad_counter1.n30555 ;
    wire \quad_counter1.n30556 ;
    wire bfn_20_5_0_;
    wire \quad_counter1.n30557 ;
    wire \quad_counter1.n2809 ;
    wire \quad_counter1.n30558 ;
    wire \quad_counter1.n2808 ;
    wire \quad_counter1.n30559 ;
    wire \quad_counter1.n30560 ;
    wire \quad_counter1.n2806 ;
    wire \quad_counter1.n30561 ;
    wire \quad_counter1.n2805 ;
    wire \quad_counter1.n30562 ;
    wire \quad_counter1.n30563 ;
    wire \quad_counter1.n2804 ;
    wire \quad_counter1.n26_adj_4482 ;
    wire \quad_counter1.n3134_cascade_ ;
    wire \quad_counter1.n8_adj_4477 ;
    wire \quad_counter1.n7_adj_4478 ;
    wire \quad_counter1.n34587_cascade_ ;
    wire \quad_counter1.n22_adj_4481 ;
    wire bfn_20_8_0_;
    wire \quad_counter1.n3119 ;
    wire \quad_counter1.n30615 ;
    wire \quad_counter1.n3118 ;
    wire \quad_counter1.n30616 ;
    wire \quad_counter1.n3117 ;
    wire \quad_counter1.n3216 ;
    wire \quad_counter1.n30617 ;
    wire \quad_counter1.n3116 ;
    wire \quad_counter1.n3215 ;
    wire \quad_counter1.n30618 ;
    wire \quad_counter1.n3115 ;
    wire \quad_counter1.n30619 ;
    wire \quad_counter1.n3114 ;
    wire \quad_counter1.n36152 ;
    wire \quad_counter1.n3213 ;
    wire \quad_counter1.n30620 ;
    wire \quad_counter1.n3113 ;
    wire \quad_counter1.n3212 ;
    wire \quad_counter1.n30621 ;
    wire \quad_counter1.n30622 ;
    wire \quad_counter1.n3112 ;
    wire \quad_counter1.n3211 ;
    wire bfn_20_9_0_;
    wire \quad_counter1.n3111 ;
    wire \quad_counter1.n3210 ;
    wire \quad_counter1.n30623 ;
    wire \quad_counter1.n3110 ;
    wire \quad_counter1.n3209 ;
    wire \quad_counter1.n30624 ;
    wire \quad_counter1.n3109 ;
    wire \quad_counter1.n3208 ;
    wire \quad_counter1.n30625 ;
    wire \quad_counter1.n3108 ;
    wire \quad_counter1.n3207 ;
    wire \quad_counter1.n30626 ;
    wire \quad_counter1.n3107 ;
    wire \quad_counter1.n3206 ;
    wire \quad_counter1.n30627 ;
    wire \quad_counter1.n3106 ;
    wire \quad_counter1.n3205 ;
    wire \quad_counter1.n30628 ;
    wire \quad_counter1.n3105 ;
    wire \quad_counter1.n3204 ;
    wire \quad_counter1.n30629 ;
    wire \quad_counter1.n30630 ;
    wire \quad_counter1.n3104 ;
    wire \quad_counter1.n3203 ;
    wire bfn_20_10_0_;
    wire \quad_counter1.n3103 ;
    wire \quad_counter1.n3202 ;
    wire \quad_counter1.n30631 ;
    wire \quad_counter1.n3102 ;
    wire \quad_counter1.n3201 ;
    wire \quad_counter1.n30632 ;
    wire \quad_counter1.n3101 ;
    wire \quad_counter1.n3134 ;
    wire \quad_counter1.n30633 ;
    wire \quad_counter1.n3200 ;
    wire \quad_counter0.n3117 ;
    wire \quad_counter0.n3114 ;
    wire \quad_counter0.n8 ;
    wire \quad_counter0.n2417 ;
    wire \quad_counter0.n2414 ;
    wire \quad_counter0.n8_adj_4394 ;
    wire \c0.n4_adj_4623 ;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.n32750 ;
    wire \quad_counter1.n8 ;
    wire \quad_counter1.n8_adj_4444 ;
    wire \quad_counter1.n35309_cascade_ ;
    wire \quad_counter1.n7 ;
    wire n10_adj_4821;
    wire byte_transmit_counter_5;
    wire n14821;
    wire r_Tx_Data_5;
    wire \quad_counter1.n35603 ;
    wire \c0.n35824 ;
    wire \c0.n26_adj_4625_cascade_ ;
    wire n35826;
    wire n2274;
    wire data_out_frame_7_1;
    wire \c0.n5_adj_4505_cascade_ ;
    wire \c0.n35830_cascade_ ;
    wire n35832;
    wire data_out_frame_10_5;
    wire \c0.n36016_cascade_ ;
    wire \c0.n35827_cascade_ ;
    wire n35829;
    wire n2271;
    wire data_out_frame_5_0;
    wire n2259;
    wire data_out_frame_7_7;
    wire \c0.n5_adj_4653 ;
    wire encoder1_position_22;
    wire data_out_frame_5_7;
    wire data_out_frame_5_1;
    wire \c0.n36090 ;
    wire data_out_frame_6_7;
    wire encoder0_position_1;
    wire \c0.n33503_cascade_ ;
    wire \c0.n47 ;
    wire \c0.n41_adj_4571_cascade_ ;
    wire \c0.n30_cascade_ ;
    wire \c0.n39_adj_4567 ;
    wire \c0.n45_adj_4572 ;
    wire \c0.n33314_cascade_ ;
    wire \c0.n18124 ;
    wire \c0.n24_cascade_ ;
    wire encoder0_position_19;
    wire \c0.n18 ;
    wire encoder0_position_20;
    wire \c0.n33765 ;
    wire \c0.n33765_cascade_ ;
    wire \c0.n26_adj_4559 ;
    wire \c0.n33493 ;
    wire \c0.n33493_cascade_ ;
    wire \c0.n33749 ;
    wire control_mode_1;
    wire encoder1_position_26;
    wire \c0.n33432_cascade_ ;
    wire n2248;
    wire data_out_frame_6_1;
    wire control_mode_2;
    wire control_mode_3;
    wire \c0.data_out_frame_29__7__N_738_cascade_ ;
    wire \c0.n33389 ;
    wire \c0.n22 ;
    wire \c0.n33579_cascade_ ;
    wire n2343;
    wire control_mode_7;
    wire data_in_frame_1_5;
    wire encoder0_position_10;
    wire n2328;
    wire \c0.n10_adj_4547 ;
    wire control_mode_6;
    wire \c0.n33414 ;
    wire n2322;
    wire encoder0_position_23;
    wire n2336;
    wire n2329;
    wire \c0.data_in_frame_22_4 ;
    wire \c0.data_in_frame_29_2 ;
    wire \c0.data_in_frame_29_1 ;
    wire encoder0_position_8;
    wire n2341;
    wire \c0.data_in_frame_26_3 ;
    wire \c0.data_in_frame_25_3 ;
    wire n2320;
    wire encoder0_position_25;
    wire \c0.n33233 ;
    wire \c0.data_in_frame_22_3 ;
    wire \c0.data_in_frame_28_2 ;
    wire \c0.data_in_frame_27_5 ;
    wire \c0.n9_adj_4631 ;
    wire \c0.data_in_frame_28_0 ;
    wire rx_data_6;
    wire \c0.n33539 ;
    wire \c0.n33933 ;
    wire \c0.data_in_frame_27_1 ;
    wire \c0.data_in_frame_21_1 ;
    wire \c0.data_in_frame_21_2 ;
    wire \c0.n33948 ;
    wire \c0.n33467 ;
    wire \c0.data_in_frame_27_3 ;
    wire \c0.n33678 ;
    wire \c0.data_in_frame_29_5 ;
    wire \c0.n12_adj_4518 ;
    wire \c0.data_in_frame_29_3 ;
    wire \c0.n18971 ;
    wire \c0.n33551 ;
    wire \c0.n32433 ;
    wire \c0.n33762 ;
    wire \c0.data_in_frame_25_0 ;
    wire \c0.n32259 ;
    wire \c0.data_in_frame_22_6 ;
    wire \c0.n32320 ;
    wire \c0.n33563 ;
    wire \c0.data_in_frame_25_2 ;
    wire \c0.n33988_cascade_ ;
    wire \c0.n33536 ;
    wire \c0.data_in_frame_24_7 ;
    wire rx_data_1;
    wire \c0.data_in_frame_25_1 ;
    wire rx_data_5;
    wire \c0.n35211 ;
    wire \c0.data_in_frame_24_5 ;
    wire \c0.n33988 ;
    wire \c0.n33930_cascade_ ;
    wire \c0.n32341 ;
    wire \c0.n10_adj_4674 ;
    wire \quad_counter1.n2811 ;
    wire \quad_counter1.n2807 ;
    wire \quad_counter1.n2810 ;
    wire \quad_counter1.n2813 ;
    wire \quad_counter1.n18_adj_4457 ;
    wire \quad_counter1.n28269_cascade_ ;
    wire \quad_counter1.n10_adj_4468_cascade_ ;
    wire \quad_counter1.n36130 ;
    wire \quad_counter1.n2719 ;
    wire bfn_21_5_0_;
    wire \quad_counter1.n2718 ;
    wire \quad_counter1.n30535 ;
    wire \quad_counter1.n2717 ;
    wire \quad_counter1.n30536 ;
    wire \quad_counter1.n2716 ;
    wire \quad_counter1.n30537 ;
    wire \quad_counter1.n2715 ;
    wire \quad_counter1.n30538 ;
    wire \quad_counter1.n2714 ;
    wire \quad_counter1.n30539 ;
    wire \quad_counter1.n30540 ;
    wire \quad_counter1.n2712 ;
    wire \quad_counter1.n30541 ;
    wire \quad_counter1.n30542 ;
    wire bfn_21_6_0_;
    wire \quad_counter1.n30543 ;
    wire \quad_counter1.n30544 ;
    wire \quad_counter1.n30545 ;
    wire \quad_counter1.n30546 ;
    wire \quad_counter1.n30547 ;
    wire \quad_counter1.n30548 ;
    wire \quad_counter1.n14_cascade_ ;
    wire \quad_counter1.n28273_cascade_ ;
    wire \quad_counter1.n10_adj_4450_cascade_ ;
    wire \quad_counter1.n9_adj_4451 ;
    wire bfn_21_9_0_;
    wire \quad_counter1.n30510 ;
    wire \quad_counter1.n30511 ;
    wire \quad_counter1.n30512 ;
    wire \quad_counter1.n30513 ;
    wire \quad_counter1.n30514 ;
    wire \quad_counter1.n30515 ;
    wire \quad_counter1.n30516 ;
    wire \quad_counter1.n30517 ;
    wire bfn_21_10_0_;
    wire \quad_counter1.n30518 ;
    wire \quad_counter1.n30519 ;
    wire \quad_counter1.n30520 ;
    wire \quad_counter1.n30521 ;
    wire \quad_counter1.n36134 ;
    wire \quad_counter1.n12 ;
    wire \quad_counter1.n2441 ;
    wire n34871;
    wire count_prev_0_adj_4815;
    wire n34871_cascade_;
    wire \quad_counter1.n18_cascade_ ;
    wire \quad_counter1.n7_adj_4425 ;
    wire \quad_counter1.n8_adj_4424_cascade_ ;
    wire \quad_counter1.n25 ;
    wire \quad_counter1.n26 ;
    wire \quad_counter1.n28 ;
    wire \quad_counter1.n27 ;
    wire \quad_counter1.n3332_cascade_ ;
    wire n2275;
    wire n2277;
    wire \c0.n26_adj_4516 ;
    wire encoder0_position_7;
    wire encoder1_position_8;
    wire encoder0_position_6;
    wire \c0.n33615 ;
    wire \c0.n12_adj_4553_cascade_ ;
    wire data_out_frame_13_3;
    wire data_out_frame_29_6;
    wire n2267;
    wire data_in_frame_1_0;
    wire encoder1_position_13;
    wire encoder1_position_12;
    wire \c0.n18232_cascade_ ;
    wire n2273;
    wire count_enable_adj_4814;
    wire \c0.n33902 ;
    wire \c0.data_out_frame_29__7__N_976_cascade_ ;
    wire \c0.n33772 ;
    wire \c0.n42_adj_4570 ;
    wire \c0.n33305 ;
    wire \c0.data_out_frame_29__7__N_740 ;
    wire \c0.n18689 ;
    wire \c0.n6_adj_4560 ;
    wire \c0.n18523 ;
    wire \c0.n35113_cascade_ ;
    wire \c0.n31401 ;
    wire \c0.n12_adj_4561_cascade_ ;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.n18092 ;
    wire \c0.rx.n33168 ;
    wire r_SM_Main_2;
    wire \c0.rx.n34953 ;
    wire encoder0_position_31;
    wire encoder0_position_30;
    wire control_mode_5;
    wire encoder0_position_22;
    wire \c0.n18199 ;
    wire encoder1_position_20;
    wire \c0.data_out_frame_29__7__N_756 ;
    wire \c0.data_out_frame_29__7__N_734 ;
    wire \c0.n33425_cascade_ ;
    wire encoder0_position_18;
    wire n35693;
    wire control_mode_4;
    wire encoder1_position_27;
    wire encoder0_position_9;
    wire \c0.n17510 ;
    wire \c0.n33393 ;
    wire \c0.n33280 ;
    wire encoder1_position_28;
    wire \c0.n33496 ;
    wire \c0.n33496_cascade_ ;
    wire encoder1_position_14;
    wire \c0.n6_adj_4544_cascade_ ;
    wire n36176;
    wire n36099;
    wire data_in_frame_1_7;
    wire n2334;
    wire encoder0_position_11;
    wire n2340;
    wire n2333;
    wire encoder1_position_29;
    wire \c0.n18214 ;
    wire encoder1_position_17;
    wire encoder0_position_13;
    wire \c0.n33896 ;
    wire \c0.n33896_cascade_ ;
    wire \c0.n6_adj_4541 ;
    wire \c0.n18892 ;
    wire \c0.n33360_cascade_ ;
    wire \c0.n18181 ;
    wire \c0.n18740 ;
    wire encoder0_position_12;
    wire encoder1_position_16;
    wire encoder0_position_27;
    wire \c0.n33807 ;
    wire \c0.n6_adj_4566_cascade_ ;
    wire encoder0_position_29;
    wire \c0.n18572 ;
    wire rx_data_3;
    wire \c0.data_in_frame_21_3 ;
    wire \c0.n27890 ;
    wire \c0.n33224 ;
    wire \c0.n12_adj_4519 ;
    wire \c0.n33224_cascade_ ;
    wire \c0.data_in_frame_21_4 ;
    wire \c0.n9_adj_4628 ;
    wire n2321;
    wire encoder0_position_24;
    wire \c0.n9 ;
    wire rx_data_0;
    wire rx_data_2;
    wire \c0.n9_adj_4530 ;
    wire rx_data_7;
    wire \c0.n33257 ;
    wire \c0.data_in_frame_26_7 ;
    wire \c0.data_in_frame_26_2 ;
    wire \c0.data_in_frame_24_0 ;
    wire \c0.n17627 ;
    wire \c0.n31545 ;
    wire \c0.n31545_cascade_ ;
    wire \c0.n18578 ;
    wire \c0.data_in_frame_24_6 ;
    wire \c0.n20_adj_4698 ;
    wire \c0.n19_adj_4699_cascade_ ;
    wire \c0.n33819 ;
    wire \c0.n32_adj_4705 ;
    wire \quad_counter1.n2713 ;
    wire \quad_counter1.n2705 ;
    wire \quad_counter1.n2707 ;
    wire \quad_counter1.n2709 ;
    wire \quad_counter1.n2708 ;
    wire \quad_counter1.n16_adj_4469_cascade_ ;
    wire \quad_counter1.n2711 ;
    wire \quad_counter1.n2706 ;
    wire \quad_counter1.n14_adj_4470 ;
    wire \quad_counter1.n18_adj_4471_cascade_ ;
    wire \quad_counter1.n2710 ;
    wire \quad_counter1.n2738 ;
    wire \quad_counter1.n3219 ;
    wire \quad_counter1.n3218 ;
    wire \quad_counter1.n3214 ;
    wire \quad_counter1.n28243_cascade_ ;
    wire \quad_counter1.n3217 ;
    wire \quad_counter1.n10_adj_4483 ;
    wire \quad_counter1.n10_cascade_ ;
    wire \quad_counter1.n16_cascade_ ;
    wire \quad_counter1.n2639 ;
    wire \quad_counter1.n2639_cascade_ ;
    wire \quad_counter1.n36132 ;
    wire data_out_frame_11_3;
    wire bfn_22_7_0_;
    wire \quad_counter1.n30171 ;
    wire \quad_counter1.millisecond_counter_2 ;
    wire \quad_counter1.n30172 ;
    wire \quad_counter1.n30173 ;
    wire \quad_counter1.millisecond_counter_4 ;
    wire \quad_counter1.n30174 ;
    wire \quad_counter1.n30175 ;
    wire \quad_counter1.millisecond_counter_6 ;
    wire \quad_counter1.n30176 ;
    wire \quad_counter1.n30177 ;
    wire \quad_counter1.n30178 ;
    wire bfn_22_8_0_;
    wire \quad_counter1.n30179 ;
    wire \quad_counter1.n30180 ;
    wire \quad_counter1.millisecond_counter_11 ;
    wire \quad_counter1.n30181 ;
    wire \quad_counter1.millisecond_counter_12 ;
    wire \quad_counter1.n30182 ;
    wire \quad_counter1.millisecond_counter_13 ;
    wire \quad_counter1.n30183 ;
    wire \quad_counter1.millisecond_counter_14 ;
    wire \quad_counter1.n30184 ;
    wire \quad_counter1.millisecond_counter_15 ;
    wire \quad_counter1.n30185 ;
    wire \quad_counter1.n30186 ;
    wire \quad_counter1.millisecond_counter_16 ;
    wire bfn_22_9_0_;
    wire \quad_counter1.n30187 ;
    wire \quad_counter1.n30188 ;
    wire \quad_counter1.n30189 ;
    wire \quad_counter1.n30190 ;
    wire \quad_counter1.n30191 ;
    wire \quad_counter1.n30192 ;
    wire \quad_counter1.n30193 ;
    wire \quad_counter1.n30194 ;
    wire bfn_22_10_0_;
    wire \quad_counter1.n30195 ;
    wire \quad_counter1.n30196 ;
    wire \quad_counter1.n30197 ;
    wire \quad_counter1.n30198 ;
    wire \quad_counter1.n30199 ;
    wire \quad_counter1.n30200 ;
    wire \quad_counter1.n30201 ;
    wire bfn_22_11_0_;
    wire \quad_counter1.n30447 ;
    wire \quad_counter1.n30448 ;
    wire \quad_counter1.n12936 ;
    wire \quad_counter1.n30449 ;
    wire \quad_counter1.n30450 ;
    wire \quad_counter1.n12935 ;
    wire \quad_counter1.n8_adj_4453 ;
    wire \quad_counter1.n30451 ;
    wire \quad_counter1.n12934 ;
    wire \quad_counter1.n30452 ;
    wire \quad_counter1.n9_adj_4452 ;
    wire \quad_counter1.n35987 ;
    wire \quad_counter1.n10_adj_4454 ;
    wire \quad_counter1.n31_adj_4461_cascade_ ;
    wire \quad_counter1.n35986 ;
    wire \quad_counter1.n34_adj_4465_cascade_ ;
    wire \quad_counter1.millisecond_counter_3 ;
    wire \quad_counter1.n34207_cascade_ ;
    wire \quad_counter1.millisecond_counter_0 ;
    wire \quad_counter1.millisecond_counter_1 ;
    wire \quad_counter1.millisecond_counter_7 ;
    wire \quad_counter1.n34519_cascade_ ;
    wire \quad_counter1.millisecond_counter_5 ;
    wire \quad_counter1.n12_adj_4467 ;
    wire \quad_counter1.millisecond_counter_10 ;
    wire bfn_22_13_0_;
    wire \quad_counter1.n3319 ;
    wire \quad_counter1.n30654 ;
    wire \quad_counter1.n3318 ;
    wire \quad_counter1.n30655 ;
    wire \quad_counter1.n3317 ;
    wire \quad_counter1.n30656 ;
    wire \quad_counter1.n3316 ;
    wire \quad_counter1.n30657 ;
    wire \quad_counter1.n3315 ;
    wire \quad_counter1.n30658 ;
    wire \quad_counter1.n3314 ;
    wire \quad_counter1.n36146 ;
    wire \quad_counter1.n30659 ;
    wire \quad_counter1.n3313 ;
    wire \quad_counter1.n30660 ;
    wire \quad_counter1.n30661 ;
    wire \quad_counter1.n3312 ;
    wire bfn_22_14_0_;
    wire \quad_counter1.n3311 ;
    wire \quad_counter1.n30662 ;
    wire \quad_counter1.n3310 ;
    wire \quad_counter1.n30663 ;
    wire \quad_counter1.n3309 ;
    wire \quad_counter1.n30664 ;
    wire \quad_counter1.n3308 ;
    wire \quad_counter1.n30665 ;
    wire \quad_counter1.n3307 ;
    wire \quad_counter1.n30666 ;
    wire \quad_counter1.n3306 ;
    wire \quad_counter1.n30667 ;
    wire \quad_counter1.n3305 ;
    wire \quad_counter1.n30668 ;
    wire \quad_counter1.n30669 ;
    wire \quad_counter1.n3304 ;
    wire bfn_22_15_0_;
    wire \quad_counter1.n3303 ;
    wire \quad_counter1.n30670 ;
    wire \quad_counter1.n3302 ;
    wire \quad_counter1.n30671 ;
    wire \quad_counter1.n3301 ;
    wire \quad_counter1.n30672 ;
    wire \quad_counter1.n3300 ;
    wire \quad_counter1.n30673 ;
    wire \quad_counter1.n3299 ;
    wire \quad_counter1.n3332 ;
    wire \quad_counter1.n30674 ;
    wire \quad_counter1.n35050 ;
    wire \quad_counter1.n33_adj_4466 ;
    wire \c0.n35821 ;
    wire n35823;
    wire data_out_frame_28_3;
    wire encoder0_position_2;
    wire encoder0_position_17;
    wire encoder1_position_19;
    wire control_mode_0;
    wire \c0.n35113 ;
    wire encoder1_position_10;
    wire \c0.n33755 ;
    wire \c0.n31446_cascade_ ;
    wire encoder1_position_9;
    wire rx_data_4;
    wire \c0.n33249 ;
    wire data_in_frame_1_4;
    wire \c0.n26_adj_4654 ;
    wire encoder1_position_3;
    wire encoder1_position_11;
    wire \c0.n31673 ;
    wire \c0.n33425 ;
    wire \c0.data_out_frame_29__7__N_658_cascade_ ;
    wire encoder1_position_21;
    wire encoder0_position_3;
    wire \c0.n18218 ;
    wire encoder0_position_4;
    wire \c0.n18469_cascade_ ;
    wire \c0.n33681 ;
    wire \c0.n18241_cascade_ ;
    wire \c0.n10_adj_4528 ;
    wire \c0.n14_adj_4527_cascade_ ;
    wire \c0.n31511_cascade_ ;
    wire FRAME_MATCHER_state_31_N_2976_2;
    wire encoder1_position_1;
    wire data_out_frame_29__7__N_1482;
    wire data_out_frame_13_1;
    wire \c0.n33579 ;
    wire encoder1_position_4;
    wire \c0.n6_adj_4558_cascade_ ;
    wire encoder0_position_14;
    wire encoder1_position_5;
    wire \c0.n18499_cascade_ ;
    wire \c0.n33569_cascade_ ;
    wire encoder1_position_31;
    wire encoder0_position_0;
    wire \c0.n6_adj_4565 ;
    wire \c0.n33897 ;
    wire \c0.n31429 ;
    wire encoder1_position_2;
    wire \c0.n33897_cascade_ ;
    wire \c0.n33732 ;
    wire \c0.n33892 ;
    wire encoder0_position_15;
    wire \c0.n18895 ;
    wire encoder0_position_16;
    wire encoder1_position_18;
    wire \c0.n33353 ;
    wire \c0.n33318 ;
    wire encoder1_position_30;
    wire \c0.n33487 ;
    wire n2317;
    wire encoder0_position_28;
    wire count_enable;
    wire n2319;
    wire encoder0_position_26;
    wire \c0.n9_adj_4493 ;
    wire \quad_counter1.millisecond_counter_17 ;
    wire \quad_counter1.n28271_cascade_ ;
    wire \quad_counter1.n10_adj_4423_cascade_ ;
    wire \quad_counter1.n11 ;
    wire \quad_counter1.millisecond_counter_18 ;
    wire \quad_counter1.n2619 ;
    wire bfn_23_7_0_;
    wire \quad_counter1.n2519 ;
    wire \quad_counter1.n2618 ;
    wire \quad_counter1.n30522 ;
    wire \quad_counter1.n2518 ;
    wire \quad_counter1.n2617 ;
    wire \quad_counter1.n30523 ;
    wire \quad_counter1.n2517 ;
    wire \quad_counter1.n2616 ;
    wire \quad_counter1.n30524 ;
    wire \quad_counter1.n2516 ;
    wire \quad_counter1.n2615 ;
    wire \quad_counter1.n30525 ;
    wire \quad_counter1.n2515 ;
    wire \quad_counter1.n2614 ;
    wire \quad_counter1.n30526 ;
    wire \quad_counter1.n2514 ;
    wire \quad_counter1.n2613 ;
    wire \quad_counter1.n30527 ;
    wire \quad_counter1.n2513 ;
    wire \quad_counter1.n2612 ;
    wire \quad_counter1.n30528 ;
    wire \quad_counter1.n30529 ;
    wire \quad_counter1.n2512 ;
    wire \quad_counter1.n2611 ;
    wire bfn_23_8_0_;
    wire \quad_counter1.n2511 ;
    wire \quad_counter1.n2610 ;
    wire \quad_counter1.n30530 ;
    wire \quad_counter1.n2510 ;
    wire \quad_counter1.n2609 ;
    wire \quad_counter1.n30531 ;
    wire \quad_counter1.n2509 ;
    wire \quad_counter1.n2608 ;
    wire \quad_counter1.n30532 ;
    wire \quad_counter1.n2508 ;
    wire \quad_counter1.n2607 ;
    wire \quad_counter1.n30533 ;
    wire \quad_counter1.n2507 ;
    wire \quad_counter1.n30534 ;
    wire \quad_counter1.n2606 ;
    wire \quad_counter1.n2540 ;
    wire \quad_counter1.n36133 ;
    wire bfn_23_9_0_;
    wire \quad_counter1.n30499 ;
    wire \quad_counter1.n2417 ;
    wire \quad_counter1.n30500 ;
    wire \quad_counter1.n2416 ;
    wire \quad_counter1.n30501 ;
    wire \quad_counter1.n2415 ;
    wire \quad_counter1.n30502 ;
    wire \quad_counter1.n2414 ;
    wire \quad_counter1.n30503 ;
    wire \quad_counter1.n2413 ;
    wire \quad_counter1.n30504 ;
    wire \quad_counter1.n2412 ;
    wire \quad_counter1.n30505 ;
    wire \quad_counter1.n30506 ;
    wire \quad_counter1.n2411 ;
    wire bfn_23_10_0_;
    wire \quad_counter1.n2410 ;
    wire \quad_counter1.n30507 ;
    wire \quad_counter1.n2409 ;
    wire \quad_counter1.n30508 ;
    wire \quad_counter1.n30509 ;
    wire \quad_counter1.n2408 ;
    wire \quad_counter1.millisecond_counter_19 ;
    wire \quad_counter1.n2418 ;
    wire \quad_counter1.n2419 ;
    wire \quad_counter1.n7_adj_4445 ;
    wire \quad_counter1.n36135 ;
    wire \quad_counter1.n28_adj_4460 ;
    wire \quad_counter1.millisecond_counter_20 ;
    wire \quad_counter1.n28277_cascade_ ;
    wire \quad_counter1.n10_adj_4437_cascade_ ;
    wire \quad_counter1.n7_adj_4439_cascade_ ;
    wire \quad_counter1.n2342 ;
    wire \quad_counter1.millisecond_counter_9 ;
    wire bfn_23_12_0_;
    wire \quad_counter1.n3419 ;
    wire \quad_counter1.n30675 ;
    wire \quad_counter1.n3418 ;
    wire \quad_counter1.n30676 ;
    wire \quad_counter1.n3417 ;
    wire \quad_counter1.n30677 ;
    wire \quad_counter1.n3416 ;
    wire \quad_counter1.n30678 ;
    wire \quad_counter1.n3415 ;
    wire \quad_counter1.n30679 ;
    wire \quad_counter1.n3414 ;
    wire \quad_counter1.n3513 ;
    wire \quad_counter1.n30680 ;
    wire \quad_counter1.n3512 ;
    wire \quad_counter1.n30681 ;
    wire \quad_counter1.n30682 ;
    wire \quad_counter1.n3412 ;
    wire bfn_23_13_0_;
    wire \quad_counter1.n3510 ;
    wire \quad_counter1.n30683 ;
    wire \quad_counter1.n3410 ;
    wire \quad_counter1.n30684 ;
    wire \quad_counter1.n3409 ;
    wire \quad_counter1.n3508 ;
    wire \quad_counter1.n30685 ;
    wire \quad_counter1.n3408 ;
    wire \quad_counter1.n3507 ;
    wire \quad_counter1.n30686 ;
    wire \quad_counter1.n30687 ;
    wire \quad_counter1.n3406 ;
    wire \quad_counter1.n30688 ;
    wire \quad_counter1.n3504 ;
    wire \quad_counter1.n30689 ;
    wire \quad_counter1.n30690 ;
    wire \quad_counter1.n3404 ;
    wire \quad_counter1.n3503 ;
    wire bfn_23_14_0_;
    wire \quad_counter1.n3403 ;
    wire \quad_counter1.n3502 ;
    wire \quad_counter1.n30691 ;
    wire \quad_counter1.n3402 ;
    wire \quad_counter1.n3501 ;
    wire \quad_counter1.n30692 ;
    wire \quad_counter1.n3401 ;
    wire \quad_counter1.n3500 ;
    wire \quad_counter1.n30693 ;
    wire \quad_counter1.n3400 ;
    wire \quad_counter1.n3499 ;
    wire \quad_counter1.n30694 ;
    wire \quad_counter1.n3399 ;
    wire \quad_counter1.n3498 ;
    wire \quad_counter1.n30695 ;
    wire \quad_counter1.n3398 ;
    wire \quad_counter1.n30696 ;
    wire \quad_counter1.n3506 ;
    wire \quad_counter1.n3511 ;
    wire \quad_counter1.n3497_cascade_ ;
    wire \quad_counter1.n3505 ;
    wire \quad_counter1.n30_adj_4463 ;
    wire \quad_counter1.n12_adj_4464_cascade_ ;
    wire \quad_counter1.n35985 ;
    wire \quad_counter1.n3407 ;
    wire \quad_counter1.n3405 ;
    wire \quad_counter1.n3411 ;
    wire \quad_counter1.n3413 ;
    wire \quad_counter1.n30_adj_4426 ;
    wire \quad_counter1.n28_adj_4427 ;
    wire \quad_counter1.n29_adj_4428_cascade_ ;
    wire \quad_counter1.n27_adj_4429 ;
    wire \quad_counter1.n3431 ;
    wire \quad_counter1.n3431_cascade_ ;
    wire \quad_counter1.n36142 ;
    wire \quad_counter1.millisecond_counter_8 ;
    wire \quad_counter1.n3519 ;
    wire \quad_counter1.n3514 ;
    wire \quad_counter1.n3517 ;
    wire \quad_counter1.n28415_cascade_ ;
    wire \quad_counter1.n3518 ;
    wire \quad_counter1.n3515 ;
    wire \quad_counter1.n3509 ;
    wire \quad_counter1.n10_adj_4462_cascade_ ;
    wire \quad_counter1.n3516 ;
    wire \quad_counter1.n21 ;
    wire data_out_frame_13_2;
    wire data_out_frame_12_2;
    wire \c0.n11_adj_4513 ;
    wire \c0.n9_adj_4552 ;
    wire \c0.n31299 ;
    wire \c0.n31299_cascade_ ;
    wire \c0.data_out_frame_28_6 ;
    wire \c0.n32238 ;
    wire \c0.n32238_cascade_ ;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.byte_transmit_counter_2 ;
    wire data_out_frame_21_0;
    wire \c0.n14078_cascade_ ;
    wire data_out_frame_17_0;
    wire \c0.n41_adj_4642_cascade_ ;
    wire \c0.n43_adj_4641 ;
    wire \c0.n40_adj_4643 ;
    wire \c0.n39_adj_4644 ;
    wire \c0.n50_cascade_ ;
    wire \c0.n45_adj_4645 ;
    wire \c0.n18083 ;
    wire \c0.n17669 ;
    wire n17453;
    wire n36101;
    wire n26_cascade_;
    wire byte_transmit_counter_4;
    wire n36102;
    wire \c0.n17570 ;
    wire \c0.n14_adj_4522_cascade_ ;
    wire \c0.n9_adj_4524_cascade_ ;
    wire \c0.data_out_frame_29_4 ;
    wire \c0.n33795 ;
    wire \c0.n42_adj_4640 ;
    wire \c0.n18469 ;
    wire \c0.n161 ;
    wire bfn_24_1_0_;
    wire \c0.n29970 ;
    wire \c0.n29970_THRU_CRY_0_THRU_CO ;
    wire \c0.n29970_THRU_CRY_1_THRU_CO ;
    wire \c0.n29970_THRU_CRY_2_THRU_CO ;
    wire \c0.n29970_THRU_CRY_3_THRU_CO ;
    wire \c0.n29970_THRU_CRY_4_THRU_CO ;
    wire \c0.n29970_THRU_CRY_5_THRU_CO ;
    wire \c0.n29970_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire bfn_24_2_0_;
    wire \c0.n3_adj_4579 ;
    wire \c0.n29971 ;
    wire \c0.n29971_THRU_CRY_0_THRU_CO ;
    wire \c0.n29971_THRU_CRY_1_THRU_CO ;
    wire \c0.n29971_THRU_CRY_2_THRU_CO ;
    wire \c0.n29971_THRU_CRY_3_THRU_CO ;
    wire \c0.n29971_THRU_CRY_4_THRU_CO ;
    wire \c0.n29971_THRU_CRY_5_THRU_CO ;
    wire \c0.n29971_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire bfn_24_3_0_;
    wire \c0.n3_adj_4580 ;
    wire \c0.n29972 ;
    wire \c0.n29972_THRU_CRY_0_THRU_CO ;
    wire \c0.n29972_THRU_CRY_1_THRU_CO ;
    wire \c0.n29972_THRU_CRY_2_THRU_CO ;
    wire \c0.n29972_THRU_CRY_3_THRU_CO ;
    wire \c0.n29972_THRU_CRY_4_THRU_CO ;
    wire \c0.n29972_THRU_CRY_5_THRU_CO ;
    wire \c0.n29972_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire bfn_24_4_0_;
    wire \c0.n3_adj_4581 ;
    wire \c0.n29973 ;
    wire \c0.n29973_THRU_CRY_0_THRU_CO ;
    wire \c0.n29973_THRU_CRY_1_THRU_CO ;
    wire \c0.n29973_THRU_CRY_2_THRU_CO ;
    wire \c0.n29973_THRU_CRY_3_THRU_CO ;
    wire \c0.n29973_THRU_CRY_4_THRU_CO ;
    wire \c0.n29973_THRU_CRY_5_THRU_CO ;
    wire \c0.n29973_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire bfn_24_5_0_;
    wire \c0.n3_adj_4583 ;
    wire \c0.n29974 ;
    wire \c0.n29974_THRU_CRY_0_THRU_CO ;
    wire \c0.n29974_THRU_CRY_1_THRU_CO ;
    wire \c0.n29974_THRU_CRY_2_THRU_CO ;
    wire \c0.n29974_THRU_CRY_3_THRU_CO ;
    wire \c0.n29974_THRU_CRY_4_THRU_CO ;
    wire \c0.n29974_THRU_CRY_5_THRU_CO ;
    wire \c0.n29974_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire bfn_24_6_0_;
    wire \c0.n3_adj_4584 ;
    wire \c0.n29975 ;
    wire \c0.n29975_THRU_CRY_0_THRU_CO ;
    wire \c0.n29975_THRU_CRY_1_THRU_CO ;
    wire \c0.n29975_THRU_CRY_2_THRU_CO ;
    wire \c0.n29975_THRU_CRY_3_THRU_CO ;
    wire \c0.n29975_THRU_CRY_4_THRU_CO ;
    wire \c0.n29975_THRU_CRY_5_THRU_CO ;
    wire \c0.n29975_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire bfn_24_7_0_;
    wire \c0.n3_adj_4585 ;
    wire \c0.n29976 ;
    wire \c0.n29976_THRU_CRY_0_THRU_CO ;
    wire \c0.n29976_THRU_CRY_1_THRU_CO ;
    wire \c0.n29976_THRU_CRY_2_THRU_CO ;
    wire \c0.n29976_THRU_CRY_3_THRU_CO ;
    wire \c0.n29976_THRU_CRY_4_THRU_CO ;
    wire \c0.n29976_THRU_CRY_5_THRU_CO ;
    wire \c0.n29976_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire bfn_24_8_0_;
    wire \c0.n3_adj_4586 ;
    wire \c0.n29977 ;
    wire \c0.n29977_THRU_CRY_0_THRU_CO ;
    wire \c0.n29977_THRU_CRY_1_THRU_CO ;
    wire \c0.n29977_THRU_CRY_2_THRU_CO ;
    wire \c0.n29977_THRU_CRY_3_THRU_CO ;
    wire \c0.n29977_THRU_CRY_4_THRU_CO ;
    wire \c0.n29977_THRU_CRY_5_THRU_CO ;
    wire \c0.n29977_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire bfn_24_9_0_;
    wire \c0.n3_adj_4587 ;
    wire \c0.n29978 ;
    wire \c0.n29978_THRU_CRY_0_THRU_CO ;
    wire \c0.n29978_THRU_CRY_1_THRU_CO ;
    wire \c0.n29978_THRU_CRY_2_THRU_CO ;
    wire \c0.n29978_THRU_CRY_3_THRU_CO ;
    wire \c0.n29978_THRU_CRY_4_THRU_CO ;
    wire \c0.n29978_THRU_CRY_5_THRU_CO ;
    wire \c0.n29978_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire bfn_24_10_0_;
    wire \c0.n3_adj_4588 ;
    wire \c0.n29979 ;
    wire \c0.n29979_THRU_CRY_0_THRU_CO ;
    wire \c0.n29979_THRU_CRY_1_THRU_CO ;
    wire \c0.n29979_THRU_CRY_2_THRU_CO ;
    wire \c0.n29979_THRU_CRY_3_THRU_CO ;
    wire \c0.n29979_THRU_CRY_4_THRU_CO ;
    wire \c0.n29979_THRU_CRY_5_THRU_CO ;
    wire \c0.n29979_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire bfn_24_11_0_;
    wire \c0.n3_adj_4589 ;
    wire \c0.n29980 ;
    wire \c0.n29980_THRU_CRY_0_THRU_CO ;
    wire \c0.n29980_THRU_CRY_1_THRU_CO ;
    wire \c0.n29980_THRU_CRY_2_THRU_CO ;
    wire \c0.n29980_THRU_CRY_3_THRU_CO ;
    wire \c0.n29980_THRU_CRY_4_THRU_CO ;
    wire \c0.n29980_THRU_CRY_5_THRU_CO ;
    wire \c0.n29980_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire bfn_24_12_0_;
    wire \c0.n3_adj_4590 ;
    wire \c0.n29981 ;
    wire \c0.n29981_THRU_CRY_0_THRU_CO ;
    wire \c0.n29981_THRU_CRY_1_THRU_CO ;
    wire \c0.n29981_THRU_CRY_2_THRU_CO ;
    wire \c0.n29981_THRU_CRY_3_THRU_CO ;
    wire \c0.n29981_THRU_CRY_4_THRU_CO ;
    wire \c0.n29981_THRU_CRY_5_THRU_CO ;
    wire \c0.n29981_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire bfn_24_13_0_;
    wire \c0.n3_adj_4591 ;
    wire \c0.n29982 ;
    wire \c0.n29982_THRU_CRY_0_THRU_CO ;
    wire \c0.n29982_THRU_CRY_1_THRU_CO ;
    wire \c0.n29982_THRU_CRY_2_THRU_CO ;
    wire \c0.n29982_THRU_CRY_3_THRU_CO ;
    wire \c0.n29982_THRU_CRY_4_THRU_CO ;
    wire \c0.n29982_THRU_CRY_5_THRU_CO ;
    wire \c0.n29982_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire bfn_24_14_0_;
    wire \c0.n3_adj_4592 ;
    wire \c0.n29983 ;
    wire \c0.n29983_THRU_CRY_0_THRU_CO ;
    wire \c0.n29983_THRU_CRY_1_THRU_CO ;
    wire \c0.n29983_THRU_CRY_2_THRU_CO ;
    wire \c0.n29983_THRU_CRY_3_THRU_CO ;
    wire \c0.n29983_THRU_CRY_4_THRU_CO ;
    wire \c0.n29983_THRU_CRY_5_THRU_CO ;
    wire \c0.n29983_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire bfn_24_15_0_;
    wire \c0.n3_adj_4593 ;
    wire \c0.n29984 ;
    wire \c0.n29984_THRU_CRY_0_THRU_CO ;
    wire \c0.n29984_THRU_CRY_1_THRU_CO ;
    wire \c0.n29984_THRU_CRY_2_THRU_CO ;
    wire \c0.n29984_THRU_CRY_3_THRU_CO ;
    wire \c0.n29984_THRU_CRY_4_THRU_CO ;
    wire \c0.n29984_THRU_CRY_5_THRU_CO ;
    wire \c0.n29984_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire bfn_24_16_0_;
    wire \c0.n3_adj_4594 ;
    wire \c0.n29985 ;
    wire \c0.n29985_THRU_CRY_0_THRU_CO ;
    wire \c0.n29985_THRU_CRY_1_THRU_CO ;
    wire \c0.n29985_THRU_CRY_2_THRU_CO ;
    wire \c0.n29985_THRU_CRY_3_THRU_CO ;
    wire \c0.n29985_THRU_CRY_4_THRU_CO ;
    wire \c0.n29985_THRU_CRY_5_THRU_CO ;
    wire \c0.n29985_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire bfn_24_17_0_;
    wire \c0.n3_adj_4595 ;
    wire \c0.n29986 ;
    wire \c0.n29986_THRU_CRY_0_THRU_CO ;
    wire \c0.n29986_THRU_CRY_1_THRU_CO ;
    wire \c0.n29986_THRU_CRY_2_THRU_CO ;
    wire \c0.n29986_THRU_CRY_3_THRU_CO ;
    wire \c0.n29986_THRU_CRY_4_THRU_CO ;
    wire \c0.n29986_THRU_CRY_5_THRU_CO ;
    wire \c0.n29986_THRU_CRY_6_THRU_CO ;
    wire bfn_24_18_0_;
    wire \c0.n29987 ;
    wire \c0.n29987_THRU_CRY_0_THRU_CO ;
    wire \c0.n29987_THRU_CRY_1_THRU_CO ;
    wire \c0.n29987_THRU_CRY_2_THRU_CO ;
    wire \c0.n29987_THRU_CRY_3_THRU_CO ;
    wire \c0.n29987_THRU_CRY_4_THRU_CO ;
    wire \c0.n29987_THRU_CRY_5_THRU_CO ;
    wire \c0.n29987_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire bfn_24_19_0_;
    wire \c0.n3_adj_4597 ;
    wire \c0.n29988 ;
    wire \c0.n29988_THRU_CRY_0_THRU_CO ;
    wire \c0.n29988_THRU_CRY_1_THRU_CO ;
    wire \c0.n29988_THRU_CRY_2_THRU_CO ;
    wire \c0.n29988_THRU_CRY_3_THRU_CO ;
    wire \c0.n29988_THRU_CRY_4_THRU_CO ;
    wire \c0.n29988_THRU_CRY_5_THRU_CO ;
    wire \c0.n29988_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire bfn_24_20_0_;
    wire \c0.n3_adj_4598 ;
    wire \c0.n29989 ;
    wire \c0.n29989_THRU_CRY_0_THRU_CO ;
    wire \c0.n29989_THRU_CRY_1_THRU_CO ;
    wire \c0.n29989_THRU_CRY_2_THRU_CO ;
    wire \c0.n29989_THRU_CRY_3_THRU_CO ;
    wire \c0.n29989_THRU_CRY_4_THRU_CO ;
    wire \c0.n29989_THRU_CRY_5_THRU_CO ;
    wire \c0.n29989_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire bfn_24_21_0_;
    wire \c0.n3_adj_4599 ;
    wire \c0.n29990 ;
    wire \c0.n29990_THRU_CRY_0_THRU_CO ;
    wire \c0.n29990_THRU_CRY_1_THRU_CO ;
    wire \c0.n29990_THRU_CRY_2_THRU_CO ;
    wire \c0.n29990_THRU_CRY_3_THRU_CO ;
    wire \c0.n29990_THRU_CRY_4_THRU_CO ;
    wire \c0.n29990_THRU_CRY_5_THRU_CO ;
    wire \c0.n29990_THRU_CRY_6_THRU_CO ;
    wire bfn_24_22_0_;
    wire \c0.n29991 ;
    wire \c0.n29991_THRU_CRY_0_THRU_CO ;
    wire \c0.n29991_THRU_CRY_1_THRU_CO ;
    wire \c0.n29991_THRU_CRY_2_THRU_CO ;
    wire \c0.n29991_THRU_CRY_3_THRU_CO ;
    wire \c0.n29991_THRU_CRY_4_THRU_CO ;
    wire \c0.n29991_THRU_CRY_5_THRU_CO ;
    wire \c0.n29991_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire bfn_24_23_0_;
    wire \c0.n3_adj_4601 ;
    wire \c0.n29992 ;
    wire \c0.n29992_THRU_CRY_0_THRU_CO ;
    wire \c0.n29992_THRU_CRY_1_THRU_CO ;
    wire \c0.n29992_THRU_CRY_2_THRU_CO ;
    wire \c0.n29992_THRU_CRY_3_THRU_CO ;
    wire \c0.n29992_THRU_CRY_4_THRU_CO ;
    wire \c0.n29992_THRU_CRY_5_THRU_CO ;
    wire \c0.n29992_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire bfn_24_24_0_;
    wire \c0.n3_adj_4602 ;
    wire \c0.n29993 ;
    wire \c0.n29993_THRU_CRY_0_THRU_CO ;
    wire \c0.n29993_THRU_CRY_1_THRU_CO ;
    wire \c0.n29993_THRU_CRY_2_THRU_CO ;
    wire \c0.n29993_THRU_CRY_3_THRU_CO ;
    wire \c0.n29993_THRU_CRY_4_THRU_CO ;
    wire \c0.n29993_THRU_CRY_5_THRU_CO ;
    wire \c0.n29993_THRU_CRY_6_THRU_CO ;
    wire bfn_24_25_0_;
    wire \c0.n3_adj_4603 ;
    wire \c0.n29994 ;
    wire \c0.n29994_THRU_CRY_0_THRU_CO ;
    wire \c0.n29994_THRU_CRY_1_THRU_CO ;
    wire \c0.n29994_THRU_CRY_2_THRU_CO ;
    wire \c0.n29994_THRU_CRY_3_THRU_CO ;
    wire \c0.n29994_THRU_CRY_4_THRU_CO ;
    wire \c0.n29994_THRU_CRY_5_THRU_CO ;
    wire \c0.n29994_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire bfn_24_26_0_;
    wire \c0.n3_adj_4604 ;
    wire \c0.n29995 ;
    wire \c0.n29995_THRU_CRY_0_THRU_CO ;
    wire \c0.n29995_THRU_CRY_1_THRU_CO ;
    wire \c0.n29995_THRU_CRY_2_THRU_CO ;
    wire \c0.n29995_THRU_CRY_3_THRU_CO ;
    wire \c0.n29995_THRU_CRY_4_THRU_CO ;
    wire \c0.n29995_THRU_CRY_5_THRU_CO ;
    wire \c0.n29995_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire bfn_24_27_0_;
    wire \c0.n3_adj_4605 ;
    wire \c0.n29996 ;
    wire \c0.n29996_THRU_CRY_0_THRU_CO ;
    wire \c0.n29996_THRU_CRY_1_THRU_CO ;
    wire \c0.n29996_THRU_CRY_2_THRU_CO ;
    wire \c0.n29996_THRU_CRY_3_THRU_CO ;
    wire \c0.n29996_THRU_CRY_4_THRU_CO ;
    wire \c0.n29996_THRU_CRY_5_THRU_CO ;
    wire \c0.n29996_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire bfn_24_28_0_;
    wire \c0.n3_adj_4606 ;
    wire \c0.n29997 ;
    wire \c0.n29997_THRU_CRY_0_THRU_CO ;
    wire \c0.n29997_THRU_CRY_1_THRU_CO ;
    wire \c0.n29997_THRU_CRY_2_THRU_CO ;
    wire \c0.n29997_THRU_CRY_3_THRU_CO ;
    wire \c0.n29997_THRU_CRY_4_THRU_CO ;
    wire \c0.n29997_THRU_CRY_5_THRU_CO ;
    wire \c0.n29997_THRU_CRY_6_THRU_CO ;
    wire bfn_24_29_0_;
    wire \c0.n29998 ;
    wire \c0.n29998_THRU_CRY_0_THRU_CO ;
    wire \c0.n29998_THRU_CRY_1_THRU_CO ;
    wire \c0.n29998_THRU_CRY_2_THRU_CO ;
    wire \c0.n29998_THRU_CRY_3_THRU_CO ;
    wire \c0.n29998_THRU_CRY_4_THRU_CO ;
    wire \c0.n29998_THRU_CRY_5_THRU_CO ;
    wire \c0.n29998_THRU_CRY_6_THRU_CO ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire bfn_24_30_0_;
    wire \c0.n3_adj_4608 ;
    wire \c0.n29999 ;
    wire \c0.n29999_THRU_CRY_0_THRU_CO ;
    wire \c0.n29999_THRU_CRY_1_THRU_CO ;
    wire \c0.n29999_THRU_CRY_2_THRU_CO ;
    wire \c0.n29999_THRU_CRY_3_THRU_CO ;
    wire \c0.n29999_THRU_CRY_4_THRU_CO ;
    wire \c0.n29999_THRU_CRY_5_THRU_CO ;
    wire \c0.n29999_THRU_CRY_6_THRU_CO ;
    wire bfn_24_31_0_;
    wire \c0.n3_adj_4609 ;
    wire \c0.n30000 ;
    wire \c0.n30000_THRU_CRY_0_THRU_CO ;
    wire \c0.n30000_THRU_CRY_1_THRU_CO ;
    wire \c0.n30000_THRU_CRY_2_THRU_CO ;
    wire \c0.n30000_THRU_CRY_3_THRU_CO ;
    wire \c0.n30000_THRU_CRY_4_THRU_CO ;
    wire GNDG0;
    wire \c0.n30000_THRU_CRY_5_THRU_CO ;
    wire \c0.n30000_THRU_CRY_6_THRU_CO ;
    wire \c0.n1286 ;
    wire bfn_24_32_0_;
    wire \c0.FRAME_MATCHER_i_31 ;
    wire \c0.n3_adj_4610 ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire \c0.n3_adj_4607 ;
    wire \quad_counter1.n10_adj_4430_cascade_ ;
    wire \quad_counter1.n1847_cascade_ ;
    wire \c0.FRAME_MATCHER_i_0 ;
    wire \c0.n3 ;
    wire \quad_counter1.millisecond_counter_25 ;
    wire bfn_26_8_0_;
    wire \quad_counter1.millisecond_counter_26 ;
    wire \quad_counter1.n1847 ;
    wire \quad_counter1.n30459 ;
    wire \quad_counter1.millisecond_counter_27 ;
    wire \quad_counter1.n30460 ;
    wire \quad_counter1.millisecond_counter_28 ;
    wire \quad_counter1.n30461 ;
    wire \quad_counter1.millisecond_counter_29 ;
    wire \quad_counter1.n30462 ;
    wire \quad_counter1.millisecond_counter_30 ;
    wire \quad_counter1.n30463 ;
    wire \quad_counter1.millisecond_counter_31 ;
    wire \quad_counter1.n36138 ;
    wire \quad_counter1.n30464 ;
    wire bfn_26_9_0_;
    wire \quad_counter1.n30465 ;
    wire \quad_counter1.n30466 ;
    wire \quad_counter1.n30467 ;
    wire \quad_counter1.n30468 ;
    wire \quad_counter1.n30469 ;
    wire \quad_counter1.n30470 ;
    wire \quad_counter1.n30471 ;
    wire \quad_counter1.n28279_cascade_ ;
    wire \quad_counter1.n10_adj_4435_cascade_ ;
    wire \quad_counter1.n7_adj_4436_cascade_ ;
    wire \quad_counter1.n2243_cascade_ ;
    wire \quad_counter1.millisecond_counter_21 ;
    wire \quad_counter1.n2319 ;
    wire bfn_26_11_0_;
    wire \quad_counter1.n2318 ;
    wire \quad_counter1.n30489 ;
    wire \quad_counter1.n2317 ;
    wire \quad_counter1.n30490 ;
    wire \quad_counter1.n2316 ;
    wire \quad_counter1.n30491 ;
    wire \quad_counter1.n2315 ;
    wire \quad_counter1.n30492 ;
    wire \quad_counter1.n2314 ;
    wire \quad_counter1.n30493 ;
    wire \quad_counter1.n36136 ;
    wire \quad_counter1.n2313 ;
    wire \quad_counter1.n30494 ;
    wire \quad_counter1.n30495 ;
    wire \quad_counter1.n30496 ;
    wire \quad_counter1.n2311 ;
    wire bfn_26_12_0_;
    wire \quad_counter1.n2310 ;
    wire \quad_counter1.n30497 ;
    wire \quad_counter1.n2243 ;
    wire \quad_counter1.n30498 ;
    wire \quad_counter1.n2309 ;
    wire \quad_counter1.n2312 ;
    wire \quad_counter1.n8_adj_4438 ;
    wire \c0.n6_adj_4533_cascade_ ;
    wire \c0.data_out_frame_28_2 ;
    wire \c0.n26_adj_4512 ;
    wire \c0.n32271_cascade_ ;
    wire \c0.data_out_frame_28_1 ;
    wire \c0.n26_adj_4506 ;
    wire \c0.data_out_frame_28_4 ;
    wire \c0.n33607 ;
    wire \c0.n33379 ;
    wire \c0.n32271 ;
    wire \c0.n32300_cascade_ ;
    wire \c0.n31280 ;
    wire \c0.n32454 ;
    wire \c0.n32454_cascade_ ;
    wire \c0.n32445 ;
    wire \c0.n32331 ;
    wire \c0.n32377 ;
    wire \c0.n32300 ;
    wire \c0.n32331_cascade_ ;
    wire n35623;
    wire \c0.n4_adj_4630_cascade_ ;
    wire \c0.n4_adj_4630 ;
    wire \c0.data_out_frame_29_5 ;
    wire \c0.data_out_frame_28_5 ;
    wire \c0.n26_adj_4620 ;
    wire \c0.n32476_cascade_ ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire \c0.n44_adj_4639 ;
    wire \c0.n33572 ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire \c0.n3_adj_4596 ;
    wire \c0.n17574_cascade_ ;
    wire \c0.n35251 ;
    wire \c0.n31302 ;
    wire \c0.n32476 ;
    wire \c0.n18901 ;
    wire \c0.n14_adj_4523 ;
    wire \c0.n31463_cascade_ ;
    wire encoder1_position_6;
    wire \c0.n32361 ;
    wire \c0.n32359 ;
    wire \c0.n31466 ;
    wire \c0.n32361_cascade_ ;
    wire \c0.n32333 ;
    wire \c0.n33861 ;
    wire \c0.n21_adj_4551 ;
    wire \c0.n20_adj_4549_cascade_ ;
    wire \c0.n32410 ;
    wire \c0.n32424 ;
    wire \c0.n34466_cascade_ ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire \c0.n2107 ;
    wire \c0.n3_adj_4600 ;
    wire \c0.n18499 ;
    wire \c0.n18898 ;
    wire \quad_counter1.n1913 ;
    wire \quad_counter1.n1946_cascade_ ;
    wire \quad_counter1.n1985 ;
    wire \quad_counter1.n1984 ;
    wire \quad_counter1.n2016_cascade_ ;
    wire \quad_counter1.n1917 ;
    wire \quad_counter1.n28285_cascade_ ;
    wire \quad_counter1.n1918 ;
    wire \quad_counter1.n10_adj_4431 ;
    wire \quad_counter1.n1983 ;
    wire \quad_counter1.n1916 ;
    wire \quad_counter1.n1982 ;
    wire \quad_counter1.n1915 ;
    wire \quad_counter1.millisecond_counter_24 ;
    wire \quad_counter1.n1987 ;
    wire \quad_counter1.n2019_cascade_ ;
    wire \quad_counter1.n28283_cascade_ ;
    wire \quad_counter1.n9 ;
    wire \quad_counter1.n10_adj_4432_cascade_ ;
    wire \quad_counter1.n2045_cascade_ ;
    wire \quad_counter1.n2118_cascade_ ;
    wire \quad_counter1.n1986 ;
    wire \quad_counter1.n1919 ;
    wire \quad_counter1.millisecond_counter_22 ;
    wire \quad_counter1.n2219 ;
    wire bfn_27_11_0_;
    wire \quad_counter1.n2218 ;
    wire \quad_counter1.n30480 ;
    wire \quad_counter1.n2118 ;
    wire \quad_counter1.n2217 ;
    wire \quad_counter1.n30481 ;
    wire \quad_counter1.n2216 ;
    wire \quad_counter1.n30482 ;
    wire \quad_counter1.n2215 ;
    wire \quad_counter1.n30483 ;
    wire \quad_counter1.n2214 ;
    wire \quad_counter1.n30484 ;
    wire \quad_counter1.n2213 ;
    wire \quad_counter1.n30485 ;
    wire \quad_counter1.n2212 ;
    wire \quad_counter1.n30486 ;
    wire \quad_counter1.n30487 ;
    wire \quad_counter1.n2211 ;
    wire bfn_27_12_0_;
    wire \quad_counter1.n30488 ;
    wire \quad_counter1.n2210 ;
    wire \c0.data_out_frame_29_3 ;
    wire \c0.data_out_frame_29_1 ;
    wire \c0.data_out_frame_29__2__N_1749_cascade_ ;
    wire \c0.n31338 ;
    wire \c0.n20 ;
    wire \c0.n21_cascade_ ;
    wire \c0.n19 ;
    wire \c0.n31403 ;
    wire \c0.data_out_frame_29_2 ;
    wire \c0.n32372 ;
    wire \c0.n7_adj_4521_cascade_ ;
    wire \c0.data_out_frame_29__4__N_1639 ;
    wire \c0.n15827 ;
    wire \c0.n32383_cascade_ ;
    wire \c0.data_out_frame_29_0 ;
    wire \c0.data_out_frame_28_0 ;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.n35983 ;
    wire \c0.n4 ;
    wire \c0.n26_cascade_ ;
    wire byte_transmit_counter_3;
    wire \c0.n35819 ;
    wire \c0.n33557 ;
    wire data_out_frame_29__6__N_1518;
    wire \c0.data_out_frame_29_7 ;
    wire \c0.n10_adj_4573_cascade_ ;
    wire \c0.n31236 ;
    wire \c0.n31511 ;
    wire \c0.n33509 ;
    wire \c0.n31372 ;
    wire \c0.n31516 ;
    wire \c0.n31372_cascade_ ;
    wire \c0.n33588 ;
    wire \c0.n32437_cascade_ ;
    wire \c0.n31287 ;
    wire \c0.n32403 ;
    wire \c0.n35212 ;
    wire \c0.n33656 ;
    wire \c0.n35426 ;
    wire data_out_frame_29__7__N_1426;
    wire \c0.n16_cascade_ ;
    wire \c0.data_out_frame_28_7 ;
    wire PIN_9_c;
    wire \c0.n12483 ;
    wire \c0.n31283 ;
    wire \c0.n4_adj_4525 ;
    wire \c0.n15775 ;
    wire \c0.n17576 ;
    wire \c0.n33644_cascade_ ;
    wire \c0.n32273 ;
    wire \c0.n33855 ;
    wire \c0.n31357_cascade_ ;
    wire \c0.n33529 ;
    wire \c0.n17 ;
    wire \c0.n32383 ;
    wire \c0.n33644 ;
    wire \c0.n10_adj_4520 ;
    wire \c0.n14_adj_4562 ;
    wire encoder0_position_5;
    wire \c0.data_out_frame_29__7__N_738 ;
    wire \c0.n15 ;
    wire \c0.n31857 ;
    wire \c0.n35280_cascade_ ;
    wire \c0.n31461 ;
    wire \c0.n32337 ;
    wire \c0.n31461_cascade_ ;
    wire \c0.n33839 ;
    wire \c0.n8_adj_4529 ;
    wire \c0.n31423 ;
    wire \c0.n31387 ;
    wire \c0.n32290 ;
    wire \c0.n33670 ;
    wire \c0.n31446 ;
    wire \c0.n33670_cascade_ ;
    wire \c0.n15744 ;
    wire \c0.n14_adj_4543_cascade_ ;
    wire \c0.n18232 ;
    wire \c0.n32071 ;
    wire \c0.n31878 ;
    wire \c0.n33687 ;
    wire \c0.n19_adj_4550 ;
    wire \c0.n33746 ;
    wire encoder1_position_7;
    wire \c0.n10_adj_4542 ;
    wire bfn_28_9_0_;
    wire \quad_counter1.n2019 ;
    wire \quad_counter1.n2086 ;
    wire \quad_counter1.n30472 ;
    wire \quad_counter1.n30473 ;
    wire \quad_counter1.n30474 ;
    wire \quad_counter1.n2016 ;
    wire \quad_counter1.n2083 ;
    wire \quad_counter1.n30475 ;
    wire \quad_counter1.n30476 ;
    wire \quad_counter1.n30477 ;
    wire \quad_counter1.n30478 ;
    wire \quad_counter1.n30479 ;
    wire CONSTANT_ONE_NET;
    wire \quad_counter1.n2012 ;
    wire bfn_28_10_0_;
    wire \quad_counter1.n1914 ;
    wire \quad_counter1.n1981 ;
    wire \quad_counter1.n1946 ;
    wire \quad_counter1.n2014 ;
    wire \quad_counter1.n2081 ;
    wire \quad_counter1.millisecond_counter_23 ;
    wire \quad_counter1.n2087 ;
    wire \quad_counter1.n2119 ;
    wire \quad_counter1.n2017 ;
    wire \quad_counter1.n2084 ;
    wire \quad_counter1.n2015 ;
    wire \quad_counter1.n2082 ;
    wire \quad_counter1.n2013 ;
    wire \quad_counter1.n2080 ;
    wire \quad_counter1.n2018 ;
    wire \quad_counter1.n2045 ;
    wire \quad_counter1.n2085 ;
    wire \quad_counter1.n2117 ;
    wire \quad_counter1.n2117_cascade_ ;
    wire \quad_counter1.n2114 ;
    wire \quad_counter1.n2116 ;
    wire \quad_counter1.n7_adj_4434 ;
    wire \quad_counter1.n8_adj_4433_cascade_ ;
    wire \quad_counter1.n2115 ;
    wire \quad_counter1.n2113 ;
    wire \quad_counter1.n2112 ;
    wire \quad_counter1.n34427_cascade_ ;
    wire \quad_counter1.n2111 ;
    wire \quad_counter1.n2144 ;
    wire \quad_counter1.n2144_cascade_ ;
    wire \quad_counter1.n36137 ;
    wire \c0.n31463 ;
    wire \c0.n33960 ;
    wire \c0.n32457 ;
    wire \c0.n32412 ;
    wire \c0.n33936 ;
    wire \c0.n32355 ;
    wire \c0.n32437 ;
    wire \c0.n14 ;
    wire \c0.n15711 ;
    wire \c0.n17515 ;
    wire \c0.n33548 ;
    wire \c0.n31468 ;
    wire \c0.n33548_cascade_ ;
    wire \c0.n33635 ;
    wire encoder1_position_0;
    wire \c0.n17536 ;
    wire \c0.n15729 ;
    wire \c0.n33673_cascade_ ;
    wire \c0.n31928 ;
    wire \c0.n15782 ;
    wire \c0.n34929 ;
    wire \c0.n17684 ;
    wire \c0.n32296 ;
    wire \c0.n35280 ;
    wire \c0.n32304 ;
    wire data_out_frame_29__7__N_1240;
    wire \c0.n32275 ;
    wire \c0.n33899 ;
    wire _gnd_net_;

    defparam \pll32MHz_inst.pll32MHz_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll32MHz_inst.pll32MHz_inst .TEST_MODE=1'b0;
    defparam \pll32MHz_inst.pll32MHz_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll32MHz_inst.pll32MHz_inst .PLLOUT_SELECT="SHIFTREG_0deg";
    defparam \pll32MHz_inst.pll32MHz_inst .FILTER_RANGE=3'b001;
    defparam \pll32MHz_inst.pll32MHz_inst .FEEDBACK_PATH="PHASE_AND_DELAY";
    defparam \pll32MHz_inst.pll32MHz_inst .FDA_RELATIVE=4'b0000;
    defparam \pll32MHz_inst.pll32MHz_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll32MHz_inst.pll32MHz_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll32MHz_inst.pll32MHz_inst .DIVR=4'b0000;
    defparam \pll32MHz_inst.pll32MHz_inst .DIVQ=3'b011;
    defparam \pll32MHz_inst.pll32MHz_inst .DIVF=7'b0000001;
    defparam \pll32MHz_inst.pll32MHz_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll32MHz_inst.pll32MHz_inst  (
            .BYPASS(GNDG0),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .LOCK(),
            .PLLOUTCORE(),
            .PLLOUTGLOBAL(PIN_9_c),
            .REFERENCECLK(N__35052),
            .RESETB(N__99330),
            .SCLK(),
            .SDI(),
            .SDO());
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__101572),
            .DIN(N__101571),
            .DOUT(N__101570),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__101572),
            .PADOUT(N__101571),
            .PADIN(N__101570),
            .CLOCKENABLE(),
            .DIN0(CLK_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__101563),
            .DIN(N__101562),
            .DOUT(N__101561),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__101563),
            .PADOUT(N__101562),
            .PADIN(N__101561),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35922),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_12_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_12_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_12_pad_iopad (
            .OE(N__101554),
            .DIN(N__101553),
            .DOUT(N__101552),
            .PACKAGEPIN(PIN_12));
    defparam PIN_12_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_12_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_12_pad_preio (
            .PADOEN(N__101554),
            .PADOUT(N__101553),
            .PADIN(N__101552),
            .CLOCKENABLE(),
            .DIN0(PIN_12_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_13_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_13_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_13_pad_iopad (
            .OE(N__101545),
            .DIN(N__101544),
            .DOUT(N__101543),
            .PACKAGEPIN(PIN_13));
    defparam PIN_13_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_13_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_13_pad_preio (
            .PADOEN(N__101545),
            .PADOUT(N__101544),
            .PADIN(N__101543),
            .CLOCKENABLE(),
            .DIN0(PIN_13_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_1_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_1_pad_iopad (
            .OE(N__101536),
            .DIN(N__101535),
            .DOUT(N__101534),
            .PACKAGEPIN(PIN_1));
    defparam PIN_1_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_1_pad_preio (
            .PADOEN(N__101536),
            .PADOUT(N__101535),
            .PADIN(N__101534),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_22_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_22_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_22_pad_iopad (
            .OE(N__101527),
            .DIN(N__101526),
            .DOUT(N__101525),
            .PACKAGEPIN(PIN_22));
    defparam PIN_22_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_22_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_22_pad_preio (
            .PADOEN(N__101527),
            .PADOUT(N__101526),
            .PADIN(N__101525),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_23_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_23_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_23_pad_iopad (
            .OE(N__101518),
            .DIN(N__101517),
            .DOUT(N__101516),
            .PACKAGEPIN(PIN_23));
    defparam PIN_23_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_23_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_23_pad_preio (
            .PADOEN(N__101518),
            .PADOUT(N__101517),
            .PADIN(N__101516),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_24_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_24_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_24_pad_iopad (
            .OE(N__101509),
            .DIN(N__101508),
            .DOUT(N__101507),
            .PACKAGEPIN(PIN_24));
    defparam PIN_24_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_24_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_24_pad_preio (
            .PADOEN(N__101509),
            .PADOUT(N__101508),
            .PADIN(N__101507),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_2_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_2_pad_iopad (
            .OE(N__101500),
            .DIN(N__101499),
            .DOUT(N__101498),
            .PACKAGEPIN(PIN_2));
    defparam PIN_2_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_2_pad_preio (
            .PADOEN(N__101500),
            .PADOUT(N__101499),
            .PADIN(N__101498),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_3_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_3_pad_iopad (
            .OE(N__101491),
            .DIN(N__101490),
            .DOUT(N__101489),
            .PACKAGEPIN(PIN_3));
    defparam PIN_3_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_3_pad_preio (
            .PADOEN(N__101491),
            .PADOUT(N__101490),
            .PADIN(N__101489),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_7_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_7_pad_iopad (
            .OE(N__101482),
            .DIN(N__101481),
            .DOUT(N__101480),
            .PACKAGEPIN(PIN_7));
    defparam PIN_7_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_7_pad_preio (
            .PADOEN(N__101482),
            .PADOUT(N__101481),
            .PADIN(N__101480),
            .CLOCKENABLE(),
            .DIN0(PIN_7_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_8_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_8_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_8_pad_iopad (
            .OE(N__101473),
            .DIN(N__101472),
            .DOUT(N__101471),
            .PACKAGEPIN(PIN_8));
    defparam PIN_8_pad_preio.PIN_TYPE=6'b000001;
    defparam PIN_8_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_8_pad_preio (
            .PADOEN(N__101473),
            .PADOUT(N__101472),
            .PADIN(N__101471),
            .CLOCKENABLE(),
            .DIN0(PIN_8_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam PIN_9_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam PIN_9_pad_iopad.PULLUP=1'b0;
    IO_PAD PIN_9_pad_iopad (
            .OE(N__101464),
            .DIN(N__101463),
            .DOUT(N__101462),
            .PACKAGEPIN(PIN_9));
    defparam PIN_9_pad_preio.PIN_TYPE=6'b011001;
    defparam PIN_9_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO PIN_9_pad_preio (
            .PADOEN(N__101464),
            .PADOUT(N__101463),
            .PADIN(N__101462),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35013),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__101455),
            .DIN(N__101454),
            .DOUT(N__101453),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__101455),
            .PADOUT(N__101454),
            .PADIN(N__101453),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__101446),
            .DIN(N__101445),
            .DOUT(N__101444),
            .PACKAGEPIN(PIN_4));
    defparam hall1_input_preio.PIN_TYPE=6'b000001;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__101446),
            .PADOUT(N__101445),
            .PADIN(N__101444),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__101437),
            .DIN(N__101436),
            .DOUT(N__101435),
            .PACKAGEPIN(PIN_5));
    defparam hall2_input_preio.PIN_TYPE=6'b000001;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__101437),
            .PADOUT(N__101436),
            .PADIN(N__101435),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__101428),
            .DIN(N__101427),
            .DOUT(N__101426),
            .PACKAGEPIN(PIN_6));
    defparam hall3_input_preio.PIN_TYPE=6'b000001;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__101428),
            .PADOUT(N__101427),
            .PADIN(N__101426),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__101419),
            .DIN(N__101418),
            .DOUT(N__101417),
            .PACKAGEPIN(PIN_11));
    defparam rx_input_preio.PIN_TYPE=6'b000001;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__101419),
            .PADOUT(N__101418),
            .PADIN(N__101417),
            .CLOCKENABLE(),
            .DIN0(rx_i),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__101410),
            .DIN(N__101409),
            .DOUT(N__101408),
            .PACKAGEPIN(PIN_10));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__101410),
            .PADOUT(N__101409),
            .PADIN(N__101408),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35628),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__35025));
    CascadeMux I__25079 (
            .O(N__101391),
            .I(\c0.n33548_cascade_ ));
    InMux I__25078 (
            .O(N__101388),
            .I(N__101384));
    InMux I__25077 (
            .O(N__101387),
            .I(N__101381));
    LocalMux I__25076 (
            .O(N__101384),
            .I(N__101377));
    LocalMux I__25075 (
            .O(N__101381),
            .I(N__101374));
    InMux I__25074 (
            .O(N__101380),
            .I(N__101370));
    Span4Mux_h I__25073 (
            .O(N__101377),
            .I(N__101367));
    Span4Mux_h I__25072 (
            .O(N__101374),
            .I(N__101364));
    InMux I__25071 (
            .O(N__101373),
            .I(N__101361));
    LocalMux I__25070 (
            .O(N__101370),
            .I(N__101358));
    Odrv4 I__25069 (
            .O(N__101367),
            .I(\c0.n33635 ));
    Odrv4 I__25068 (
            .O(N__101364),
            .I(\c0.n33635 ));
    LocalMux I__25067 (
            .O(N__101361),
            .I(\c0.n33635 ));
    Odrv4 I__25066 (
            .O(N__101358),
            .I(\c0.n33635 ));
    CascadeMux I__25065 (
            .O(N__101349),
            .I(N__101344));
    InMux I__25064 (
            .O(N__101348),
            .I(N__101338));
    InMux I__25063 (
            .O(N__101347),
            .I(N__101331));
    InMux I__25062 (
            .O(N__101344),
            .I(N__101328));
    CascadeMux I__25061 (
            .O(N__101343),
            .I(N__101325));
    InMux I__25060 (
            .O(N__101342),
            .I(N__101322));
    CascadeMux I__25059 (
            .O(N__101341),
            .I(N__101318));
    LocalMux I__25058 (
            .O(N__101338),
            .I(N__101315));
    InMux I__25057 (
            .O(N__101337),
            .I(N__101312));
    InMux I__25056 (
            .O(N__101336),
            .I(N__101307));
    InMux I__25055 (
            .O(N__101335),
            .I(N__101307));
    CascadeMux I__25054 (
            .O(N__101334),
            .I(N__101304));
    LocalMux I__25053 (
            .O(N__101331),
            .I(N__101299));
    LocalMux I__25052 (
            .O(N__101328),
            .I(N__101299));
    InMux I__25051 (
            .O(N__101325),
            .I(N__101296));
    LocalMux I__25050 (
            .O(N__101322),
            .I(N__101291));
    InMux I__25049 (
            .O(N__101321),
            .I(N__101286));
    InMux I__25048 (
            .O(N__101318),
            .I(N__101286));
    Span4Mux_v I__25047 (
            .O(N__101315),
            .I(N__101281));
    LocalMux I__25046 (
            .O(N__101312),
            .I(N__101281));
    LocalMux I__25045 (
            .O(N__101307),
            .I(N__101278));
    InMux I__25044 (
            .O(N__101304),
            .I(N__101274));
    Span4Mux_v I__25043 (
            .O(N__101299),
            .I(N__101271));
    LocalMux I__25042 (
            .O(N__101296),
            .I(N__101267));
    InMux I__25041 (
            .O(N__101295),
            .I(N__101262));
    InMux I__25040 (
            .O(N__101294),
            .I(N__101262));
    Span4Mux_v I__25039 (
            .O(N__101291),
            .I(N__101255));
    LocalMux I__25038 (
            .O(N__101286),
            .I(N__101255));
    Span4Mux_h I__25037 (
            .O(N__101281),
            .I(N__101255));
    Span4Mux_v I__25036 (
            .O(N__101278),
            .I(N__101252));
    CascadeMux I__25035 (
            .O(N__101277),
            .I(N__101249));
    LocalMux I__25034 (
            .O(N__101274),
            .I(N__101246));
    Sp12to4 I__25033 (
            .O(N__101271),
            .I(N__101243));
    InMux I__25032 (
            .O(N__101270),
            .I(N__101240));
    Span4Mux_h I__25031 (
            .O(N__101267),
            .I(N__101235));
    LocalMux I__25030 (
            .O(N__101262),
            .I(N__101235));
    Span4Mux_h I__25029 (
            .O(N__101255),
            .I(N__101232));
    Span4Mux_h I__25028 (
            .O(N__101252),
            .I(N__101229));
    InMux I__25027 (
            .O(N__101249),
            .I(N__101226));
    Span12Mux_h I__25026 (
            .O(N__101246),
            .I(N__101221));
    Span12Mux_h I__25025 (
            .O(N__101243),
            .I(N__101221));
    LocalMux I__25024 (
            .O(N__101240),
            .I(N__101214));
    Span4Mux_h I__25023 (
            .O(N__101235),
            .I(N__101214));
    Span4Mux_v I__25022 (
            .O(N__101232),
            .I(N__101214));
    Odrv4 I__25021 (
            .O(N__101229),
            .I(encoder1_position_0));
    LocalMux I__25020 (
            .O(N__101226),
            .I(encoder1_position_0));
    Odrv12 I__25019 (
            .O(N__101221),
            .I(encoder1_position_0));
    Odrv4 I__25018 (
            .O(N__101214),
            .I(encoder1_position_0));
    InMux I__25017 (
            .O(N__101205),
            .I(N__101198));
    InMux I__25016 (
            .O(N__101204),
            .I(N__101191));
    InMux I__25015 (
            .O(N__101203),
            .I(N__101191));
    InMux I__25014 (
            .O(N__101202),
            .I(N__101185));
    InMux I__25013 (
            .O(N__101201),
            .I(N__101182));
    LocalMux I__25012 (
            .O(N__101198),
            .I(N__101179));
    InMux I__25011 (
            .O(N__101197),
            .I(N__101176));
    InMux I__25010 (
            .O(N__101196),
            .I(N__101173));
    LocalMux I__25009 (
            .O(N__101191),
            .I(N__101170));
    InMux I__25008 (
            .O(N__101190),
            .I(N__101165));
    InMux I__25007 (
            .O(N__101189),
            .I(N__101165));
    InMux I__25006 (
            .O(N__101188),
            .I(N__101162));
    LocalMux I__25005 (
            .O(N__101185),
            .I(N__101159));
    LocalMux I__25004 (
            .O(N__101182),
            .I(N__101156));
    Span4Mux_v I__25003 (
            .O(N__101179),
            .I(N__101151));
    LocalMux I__25002 (
            .O(N__101176),
            .I(N__101151));
    LocalMux I__25001 (
            .O(N__101173),
            .I(N__101148));
    Span4Mux_v I__25000 (
            .O(N__101170),
            .I(N__101145));
    LocalMux I__24999 (
            .O(N__101165),
            .I(N__101142));
    LocalMux I__24998 (
            .O(N__101162),
            .I(N__101137));
    Span4Mux_v I__24997 (
            .O(N__101159),
            .I(N__101137));
    Span4Mux_v I__24996 (
            .O(N__101156),
            .I(N__101134));
    Span4Mux_h I__24995 (
            .O(N__101151),
            .I(N__101131));
    Span12Mux_s10_v I__24994 (
            .O(N__101148),
            .I(N__101128));
    Span4Mux_v I__24993 (
            .O(N__101145),
            .I(N__101119));
    Span4Mux_v I__24992 (
            .O(N__101142),
            .I(N__101119));
    Span4Mux_h I__24991 (
            .O(N__101137),
            .I(N__101119));
    Span4Mux_h I__24990 (
            .O(N__101134),
            .I(N__101119));
    Odrv4 I__24989 (
            .O(N__101131),
            .I(\c0.n17536 ));
    Odrv12 I__24988 (
            .O(N__101128),
            .I(\c0.n17536 ));
    Odrv4 I__24987 (
            .O(N__101119),
            .I(\c0.n17536 ));
    InMux I__24986 (
            .O(N__101112),
            .I(N__101107));
    InMux I__24985 (
            .O(N__101111),
            .I(N__101102));
    InMux I__24984 (
            .O(N__101110),
            .I(N__101102));
    LocalMux I__24983 (
            .O(N__101107),
            .I(N__101096));
    LocalMux I__24982 (
            .O(N__101102),
            .I(N__101093));
    InMux I__24981 (
            .O(N__101101),
            .I(N__101090));
    InMux I__24980 (
            .O(N__101100),
            .I(N__101084));
    InMux I__24979 (
            .O(N__101099),
            .I(N__101084));
    Span4Mux_v I__24978 (
            .O(N__101096),
            .I(N__101079));
    Span4Mux_h I__24977 (
            .O(N__101093),
            .I(N__101079));
    LocalMux I__24976 (
            .O(N__101090),
            .I(N__101076));
    InMux I__24975 (
            .O(N__101089),
            .I(N__101073));
    LocalMux I__24974 (
            .O(N__101084),
            .I(N__101070));
    Span4Mux_h I__24973 (
            .O(N__101079),
            .I(N__101067));
    Odrv12 I__24972 (
            .O(N__101076),
            .I(\c0.n15729 ));
    LocalMux I__24971 (
            .O(N__101073),
            .I(\c0.n15729 ));
    Odrv12 I__24970 (
            .O(N__101070),
            .I(\c0.n15729 ));
    Odrv4 I__24969 (
            .O(N__101067),
            .I(\c0.n15729 ));
    CascadeMux I__24968 (
            .O(N__101058),
            .I(\c0.n33673_cascade_ ));
    InMux I__24967 (
            .O(N__101055),
            .I(N__101051));
    InMux I__24966 (
            .O(N__101054),
            .I(N__101047));
    LocalMux I__24965 (
            .O(N__101051),
            .I(N__101042));
    InMux I__24964 (
            .O(N__101050),
            .I(N__101039));
    LocalMux I__24963 (
            .O(N__101047),
            .I(N__101035));
    InMux I__24962 (
            .O(N__101046),
            .I(N__101032));
    InMux I__24961 (
            .O(N__101045),
            .I(N__101029));
    Sp12to4 I__24960 (
            .O(N__101042),
            .I(N__101024));
    LocalMux I__24959 (
            .O(N__101039),
            .I(N__101024));
    InMux I__24958 (
            .O(N__101038),
            .I(N__101021));
    Span4Mux_v I__24957 (
            .O(N__101035),
            .I(N__101018));
    LocalMux I__24956 (
            .O(N__101032),
            .I(N__101011));
    LocalMux I__24955 (
            .O(N__101029),
            .I(N__101011));
    Span12Mux_v I__24954 (
            .O(N__101024),
            .I(N__101011));
    LocalMux I__24953 (
            .O(N__101021),
            .I(N__101006));
    Span4Mux_h I__24952 (
            .O(N__101018),
            .I(N__101006));
    Odrv12 I__24951 (
            .O(N__101011),
            .I(\c0.n31928 ));
    Odrv4 I__24950 (
            .O(N__101006),
            .I(\c0.n31928 ));
    InMux I__24949 (
            .O(N__101001),
            .I(N__100992));
    InMux I__24948 (
            .O(N__101000),
            .I(N__100992));
    InMux I__24947 (
            .O(N__100999),
            .I(N__100992));
    LocalMux I__24946 (
            .O(N__100992),
            .I(N__100987));
    InMux I__24945 (
            .O(N__100991),
            .I(N__100983));
    InMux I__24944 (
            .O(N__100990),
            .I(N__100980));
    Span4Mux_h I__24943 (
            .O(N__100987),
            .I(N__100977));
    InMux I__24942 (
            .O(N__100986),
            .I(N__100974));
    LocalMux I__24941 (
            .O(N__100983),
            .I(\c0.n15782 ));
    LocalMux I__24940 (
            .O(N__100980),
            .I(\c0.n15782 ));
    Odrv4 I__24939 (
            .O(N__100977),
            .I(\c0.n15782 ));
    LocalMux I__24938 (
            .O(N__100974),
            .I(\c0.n15782 ));
    InMux I__24937 (
            .O(N__100965),
            .I(N__100962));
    LocalMux I__24936 (
            .O(N__100962),
            .I(\c0.n34929 ));
    InMux I__24935 (
            .O(N__100959),
            .I(N__100954));
    InMux I__24934 (
            .O(N__100958),
            .I(N__100950));
    InMux I__24933 (
            .O(N__100957),
            .I(N__100947));
    LocalMux I__24932 (
            .O(N__100954),
            .I(N__100944));
    InMux I__24931 (
            .O(N__100953),
            .I(N__100941));
    LocalMux I__24930 (
            .O(N__100950),
            .I(N__100937));
    LocalMux I__24929 (
            .O(N__100947),
            .I(N__100930));
    Span4Mux_v I__24928 (
            .O(N__100944),
            .I(N__100930));
    LocalMux I__24927 (
            .O(N__100941),
            .I(N__100930));
    InMux I__24926 (
            .O(N__100940),
            .I(N__100926));
    Span4Mux_h I__24925 (
            .O(N__100937),
            .I(N__100923));
    Span4Mux_h I__24924 (
            .O(N__100930),
            .I(N__100920));
    InMux I__24923 (
            .O(N__100929),
            .I(N__100917));
    LocalMux I__24922 (
            .O(N__100926),
            .I(N__100914));
    Span4Mux_h I__24921 (
            .O(N__100923),
            .I(N__100911));
    Span4Mux_h I__24920 (
            .O(N__100920),
            .I(N__100908));
    LocalMux I__24919 (
            .O(N__100917),
            .I(N__100905));
    Odrv12 I__24918 (
            .O(N__100914),
            .I(\c0.n17684 ));
    Odrv4 I__24917 (
            .O(N__100911),
            .I(\c0.n17684 ));
    Odrv4 I__24916 (
            .O(N__100908),
            .I(\c0.n17684 ));
    Odrv4 I__24915 (
            .O(N__100905),
            .I(\c0.n17684 ));
    InMux I__24914 (
            .O(N__100896),
            .I(N__100890));
    InMux I__24913 (
            .O(N__100895),
            .I(N__100890));
    LocalMux I__24912 (
            .O(N__100890),
            .I(N__100887));
    Odrv4 I__24911 (
            .O(N__100887),
            .I(\c0.n32296 ));
    InMux I__24910 (
            .O(N__100884),
            .I(N__100881));
    LocalMux I__24909 (
            .O(N__100881),
            .I(N__100875));
    InMux I__24908 (
            .O(N__100880),
            .I(N__100871));
    InMux I__24907 (
            .O(N__100879),
            .I(N__100868));
    InMux I__24906 (
            .O(N__100878),
            .I(N__100863));
    Span4Mux_h I__24905 (
            .O(N__100875),
            .I(N__100860));
    InMux I__24904 (
            .O(N__100874),
            .I(N__100857));
    LocalMux I__24903 (
            .O(N__100871),
            .I(N__100852));
    LocalMux I__24902 (
            .O(N__100868),
            .I(N__100852));
    InMux I__24901 (
            .O(N__100867),
            .I(N__100847));
    InMux I__24900 (
            .O(N__100866),
            .I(N__100847));
    LocalMux I__24899 (
            .O(N__100863),
            .I(\c0.n35280 ));
    Odrv4 I__24898 (
            .O(N__100860),
            .I(\c0.n35280 ));
    LocalMux I__24897 (
            .O(N__100857),
            .I(\c0.n35280 ));
    Odrv4 I__24896 (
            .O(N__100852),
            .I(\c0.n35280 ));
    LocalMux I__24895 (
            .O(N__100847),
            .I(\c0.n35280 ));
    CascadeMux I__24894 (
            .O(N__100836),
            .I(N__100833));
    InMux I__24893 (
            .O(N__100833),
            .I(N__100827));
    InMux I__24892 (
            .O(N__100832),
            .I(N__100827));
    LocalMux I__24891 (
            .O(N__100827),
            .I(N__100821));
    InMux I__24890 (
            .O(N__100826),
            .I(N__100818));
    InMux I__24889 (
            .O(N__100825),
            .I(N__100815));
    InMux I__24888 (
            .O(N__100824),
            .I(N__100812));
    Span4Mux_h I__24887 (
            .O(N__100821),
            .I(N__100807));
    LocalMux I__24886 (
            .O(N__100818),
            .I(N__100807));
    LocalMux I__24885 (
            .O(N__100815),
            .I(N__100801));
    LocalMux I__24884 (
            .O(N__100812),
            .I(N__100801));
    Span4Mux_v I__24883 (
            .O(N__100807),
            .I(N__100798));
    InMux I__24882 (
            .O(N__100806),
            .I(N__100795));
    Span12Mux_s11_h I__24881 (
            .O(N__100801),
            .I(N__100792));
    Span4Mux_h I__24880 (
            .O(N__100798),
            .I(N__100789));
    LocalMux I__24879 (
            .O(N__100795),
            .I(\c0.n32304 ));
    Odrv12 I__24878 (
            .O(N__100792),
            .I(\c0.n32304 ));
    Odrv4 I__24877 (
            .O(N__100789),
            .I(\c0.n32304 ));
    InMux I__24876 (
            .O(N__100782),
            .I(N__100777));
    CascadeMux I__24875 (
            .O(N__100781),
            .I(N__100773));
    CascadeMux I__24874 (
            .O(N__100780),
            .I(N__100769));
    LocalMux I__24873 (
            .O(N__100777),
            .I(N__100766));
    CascadeMux I__24872 (
            .O(N__100776),
            .I(N__100763));
    InMux I__24871 (
            .O(N__100773),
            .I(N__100760));
    InMux I__24870 (
            .O(N__100772),
            .I(N__100757));
    InMux I__24869 (
            .O(N__100769),
            .I(N__100754));
    Span4Mux_v I__24868 (
            .O(N__100766),
            .I(N__100751));
    InMux I__24867 (
            .O(N__100763),
            .I(N__100747));
    LocalMux I__24866 (
            .O(N__100760),
            .I(N__100742));
    LocalMux I__24865 (
            .O(N__100757),
            .I(N__100742));
    LocalMux I__24864 (
            .O(N__100754),
            .I(N__100739));
    Span4Mux_h I__24863 (
            .O(N__100751),
            .I(N__100736));
    CascadeMux I__24862 (
            .O(N__100750),
            .I(N__100733));
    LocalMux I__24861 (
            .O(N__100747),
            .I(N__100730));
    Span4Mux_v I__24860 (
            .O(N__100742),
            .I(N__100727));
    Span4Mux_v I__24859 (
            .O(N__100739),
            .I(N__100723));
    Sp12to4 I__24858 (
            .O(N__100736),
            .I(N__100720));
    InMux I__24857 (
            .O(N__100733),
            .I(N__100717));
    Span4Mux_h I__24856 (
            .O(N__100730),
            .I(N__100714));
    Span4Mux_h I__24855 (
            .O(N__100727),
            .I(N__100711));
    InMux I__24854 (
            .O(N__100726),
            .I(N__100708));
    Sp12to4 I__24853 (
            .O(N__100723),
            .I(N__100701));
    Span12Mux_s8_h I__24852 (
            .O(N__100720),
            .I(N__100701));
    LocalMux I__24851 (
            .O(N__100717),
            .I(N__100701));
    Span4Mux_h I__24850 (
            .O(N__100714),
            .I(N__100696));
    Span4Mux_h I__24849 (
            .O(N__100711),
            .I(N__100696));
    LocalMux I__24848 (
            .O(N__100708),
            .I(data_out_frame_29__7__N_1240));
    Odrv12 I__24847 (
            .O(N__100701),
            .I(data_out_frame_29__7__N_1240));
    Odrv4 I__24846 (
            .O(N__100696),
            .I(data_out_frame_29__7__N_1240));
    InMux I__24845 (
            .O(N__100689),
            .I(N__100686));
    LocalMux I__24844 (
            .O(N__100686),
            .I(N__100679));
    InMux I__24843 (
            .O(N__100685),
            .I(N__100674));
    InMux I__24842 (
            .O(N__100684),
            .I(N__100674));
    InMux I__24841 (
            .O(N__100683),
            .I(N__100671));
    CascadeMux I__24840 (
            .O(N__100682),
            .I(N__100667));
    Span4Mux_v I__24839 (
            .O(N__100679),
            .I(N__100662));
    LocalMux I__24838 (
            .O(N__100674),
            .I(N__100662));
    LocalMux I__24837 (
            .O(N__100671),
            .I(N__100659));
    InMux I__24836 (
            .O(N__100670),
            .I(N__100656));
    InMux I__24835 (
            .O(N__100667),
            .I(N__100653));
    Span4Mux_h I__24834 (
            .O(N__100662),
            .I(N__100650));
    Span4Mux_h I__24833 (
            .O(N__100659),
            .I(N__100647));
    LocalMux I__24832 (
            .O(N__100656),
            .I(N__100642));
    LocalMux I__24831 (
            .O(N__100653),
            .I(N__100642));
    Span4Mux_h I__24830 (
            .O(N__100650),
            .I(N__100639));
    Odrv4 I__24829 (
            .O(N__100647),
            .I(\c0.n32275 ));
    Odrv12 I__24828 (
            .O(N__100642),
            .I(\c0.n32275 ));
    Odrv4 I__24827 (
            .O(N__100639),
            .I(\c0.n32275 ));
    InMux I__24826 (
            .O(N__100632),
            .I(N__100628));
    InMux I__24825 (
            .O(N__100631),
            .I(N__100625));
    LocalMux I__24824 (
            .O(N__100628),
            .I(\c0.n33899 ));
    LocalMux I__24823 (
            .O(N__100625),
            .I(\c0.n33899 ));
    InMux I__24822 (
            .O(N__100620),
            .I(N__100616));
    InMux I__24821 (
            .O(N__100619),
            .I(N__100612));
    LocalMux I__24820 (
            .O(N__100616),
            .I(N__100609));
    InMux I__24819 (
            .O(N__100615),
            .I(N__100606));
    LocalMux I__24818 (
            .O(N__100612),
            .I(\quad_counter1.n2116 ));
    Odrv4 I__24817 (
            .O(N__100609),
            .I(\quad_counter1.n2116 ));
    LocalMux I__24816 (
            .O(N__100606),
            .I(\quad_counter1.n2116 ));
    InMux I__24815 (
            .O(N__100599),
            .I(N__100596));
    LocalMux I__24814 (
            .O(N__100596),
            .I(\quad_counter1.n7_adj_4434 ));
    CascadeMux I__24813 (
            .O(N__100593),
            .I(\quad_counter1.n8_adj_4433_cascade_ ));
    InMux I__24812 (
            .O(N__100590),
            .I(N__100586));
    InMux I__24811 (
            .O(N__100589),
            .I(N__100582));
    LocalMux I__24810 (
            .O(N__100586),
            .I(N__100579));
    InMux I__24809 (
            .O(N__100585),
            .I(N__100576));
    LocalMux I__24808 (
            .O(N__100582),
            .I(\quad_counter1.n2115 ));
    Odrv4 I__24807 (
            .O(N__100579),
            .I(\quad_counter1.n2115 ));
    LocalMux I__24806 (
            .O(N__100576),
            .I(\quad_counter1.n2115 ));
    InMux I__24805 (
            .O(N__100569),
            .I(N__100564));
    InMux I__24804 (
            .O(N__100568),
            .I(N__100561));
    InMux I__24803 (
            .O(N__100567),
            .I(N__100558));
    LocalMux I__24802 (
            .O(N__100564),
            .I(\quad_counter1.n2113 ));
    LocalMux I__24801 (
            .O(N__100561),
            .I(\quad_counter1.n2113 ));
    LocalMux I__24800 (
            .O(N__100558),
            .I(\quad_counter1.n2113 ));
    InMux I__24799 (
            .O(N__100551),
            .I(N__100546));
    InMux I__24798 (
            .O(N__100550),
            .I(N__100543));
    InMux I__24797 (
            .O(N__100549),
            .I(N__100540));
    LocalMux I__24796 (
            .O(N__100546),
            .I(\quad_counter1.n2112 ));
    LocalMux I__24795 (
            .O(N__100543),
            .I(\quad_counter1.n2112 ));
    LocalMux I__24794 (
            .O(N__100540),
            .I(\quad_counter1.n2112 ));
    CascadeMux I__24793 (
            .O(N__100533),
            .I(\quad_counter1.n34427_cascade_ ));
    InMux I__24792 (
            .O(N__100530),
            .I(N__100526));
    InMux I__24791 (
            .O(N__100529),
            .I(N__100523));
    LocalMux I__24790 (
            .O(N__100526),
            .I(N__100520));
    LocalMux I__24789 (
            .O(N__100523),
            .I(N__100514));
    Span4Mux_h I__24788 (
            .O(N__100520),
            .I(N__100514));
    InMux I__24787 (
            .O(N__100519),
            .I(N__100511));
    Odrv4 I__24786 (
            .O(N__100514),
            .I(\quad_counter1.n2111 ));
    LocalMux I__24785 (
            .O(N__100511),
            .I(\quad_counter1.n2111 ));
    CascadeMux I__24784 (
            .O(N__100506),
            .I(N__100500));
    CascadeMux I__24783 (
            .O(N__100505),
            .I(N__100497));
    CascadeMux I__24782 (
            .O(N__100504),
            .I(N__100494));
    CascadeMux I__24781 (
            .O(N__100503),
            .I(N__100491));
    InMux I__24780 (
            .O(N__100500),
            .I(N__100488));
    InMux I__24779 (
            .O(N__100497),
            .I(N__100485));
    InMux I__24778 (
            .O(N__100494),
            .I(N__100480));
    InMux I__24777 (
            .O(N__100491),
            .I(N__100480));
    LocalMux I__24776 (
            .O(N__100488),
            .I(\quad_counter1.n2144 ));
    LocalMux I__24775 (
            .O(N__100485),
            .I(\quad_counter1.n2144 ));
    LocalMux I__24774 (
            .O(N__100480),
            .I(\quad_counter1.n2144 ));
    CascadeMux I__24773 (
            .O(N__100473),
            .I(\quad_counter1.n2144_cascade_ ));
    CascadeMux I__24772 (
            .O(N__100470),
            .I(N__100462));
    CascadeMux I__24771 (
            .O(N__100469),
            .I(N__100459));
    CascadeMux I__24770 (
            .O(N__100468),
            .I(N__100456));
    CascadeMux I__24769 (
            .O(N__100467),
            .I(N__100453));
    CascadeMux I__24768 (
            .O(N__100466),
            .I(N__100450));
    CascadeMux I__24767 (
            .O(N__100465),
            .I(N__100447));
    InMux I__24766 (
            .O(N__100462),
            .I(N__100442));
    InMux I__24765 (
            .O(N__100459),
            .I(N__100442));
    InMux I__24764 (
            .O(N__100456),
            .I(N__100433));
    InMux I__24763 (
            .O(N__100453),
            .I(N__100433));
    InMux I__24762 (
            .O(N__100450),
            .I(N__100433));
    InMux I__24761 (
            .O(N__100447),
            .I(N__100433));
    LocalMux I__24760 (
            .O(N__100442),
            .I(\quad_counter1.n36137 ));
    LocalMux I__24759 (
            .O(N__100433),
            .I(\quad_counter1.n36137 ));
    CascadeMux I__24758 (
            .O(N__100428),
            .I(N__100422));
    CascadeMux I__24757 (
            .O(N__100427),
            .I(N__100419));
    InMux I__24756 (
            .O(N__100426),
            .I(N__100416));
    InMux I__24755 (
            .O(N__100425),
            .I(N__100411));
    InMux I__24754 (
            .O(N__100422),
            .I(N__100406));
    InMux I__24753 (
            .O(N__100419),
            .I(N__100406));
    LocalMux I__24752 (
            .O(N__100416),
            .I(N__100403));
    InMux I__24751 (
            .O(N__100415),
            .I(N__100400));
    InMux I__24750 (
            .O(N__100414),
            .I(N__100397));
    LocalMux I__24749 (
            .O(N__100411),
            .I(N__100392));
    LocalMux I__24748 (
            .O(N__100406),
            .I(N__100392));
    Span4Mux_v I__24747 (
            .O(N__100403),
            .I(N__100389));
    LocalMux I__24746 (
            .O(N__100400),
            .I(\c0.n31463 ));
    LocalMux I__24745 (
            .O(N__100397),
            .I(\c0.n31463 ));
    Odrv4 I__24744 (
            .O(N__100392),
            .I(\c0.n31463 ));
    Odrv4 I__24743 (
            .O(N__100389),
            .I(\c0.n31463 ));
    InMux I__24742 (
            .O(N__100380),
            .I(N__100376));
    InMux I__24741 (
            .O(N__100379),
            .I(N__100373));
    LocalMux I__24740 (
            .O(N__100376),
            .I(N__100370));
    LocalMux I__24739 (
            .O(N__100373),
            .I(N__100367));
    Span4Mux_v I__24738 (
            .O(N__100370),
            .I(N__100364));
    Odrv4 I__24737 (
            .O(N__100367),
            .I(\c0.n33960 ));
    Odrv4 I__24736 (
            .O(N__100364),
            .I(\c0.n33960 ));
    CascadeMux I__24735 (
            .O(N__100359),
            .I(N__100354));
    InMux I__24734 (
            .O(N__100358),
            .I(N__100351));
    CascadeMux I__24733 (
            .O(N__100357),
            .I(N__100348));
    InMux I__24732 (
            .O(N__100354),
            .I(N__100345));
    LocalMux I__24731 (
            .O(N__100351),
            .I(N__100342));
    InMux I__24730 (
            .O(N__100348),
            .I(N__100339));
    LocalMux I__24729 (
            .O(N__100345),
            .I(N__100336));
    Span4Mux_h I__24728 (
            .O(N__100342),
            .I(N__100331));
    LocalMux I__24727 (
            .O(N__100339),
            .I(N__100331));
    Odrv4 I__24726 (
            .O(N__100336),
            .I(\c0.n32457 ));
    Odrv4 I__24725 (
            .O(N__100331),
            .I(\c0.n32457 ));
    CascadeMux I__24724 (
            .O(N__100326),
            .I(N__100323));
    InMux I__24723 (
            .O(N__100323),
            .I(N__100320));
    LocalMux I__24722 (
            .O(N__100320),
            .I(N__100316));
    InMux I__24721 (
            .O(N__100319),
            .I(N__100313));
    Odrv4 I__24720 (
            .O(N__100316),
            .I(\c0.n32412 ));
    LocalMux I__24719 (
            .O(N__100313),
            .I(\c0.n32412 ));
    InMux I__24718 (
            .O(N__100308),
            .I(N__100305));
    LocalMux I__24717 (
            .O(N__100305),
            .I(N__100301));
    InMux I__24716 (
            .O(N__100304),
            .I(N__100298));
    Span4Mux_v I__24715 (
            .O(N__100301),
            .I(N__100295));
    LocalMux I__24714 (
            .O(N__100298),
            .I(\c0.n33936 ));
    Odrv4 I__24713 (
            .O(N__100295),
            .I(\c0.n33936 ));
    CascadeMux I__24712 (
            .O(N__100290),
            .I(N__100287));
    InMux I__24711 (
            .O(N__100287),
            .I(N__100284));
    LocalMux I__24710 (
            .O(N__100284),
            .I(\c0.n32355 ));
    InMux I__24709 (
            .O(N__100281),
            .I(N__100277));
    InMux I__24708 (
            .O(N__100280),
            .I(N__100274));
    LocalMux I__24707 (
            .O(N__100277),
            .I(\c0.n32437 ));
    LocalMux I__24706 (
            .O(N__100274),
            .I(\c0.n32437 ));
    InMux I__24705 (
            .O(N__100269),
            .I(N__100263));
    InMux I__24704 (
            .O(N__100268),
            .I(N__100263));
    LocalMux I__24703 (
            .O(N__100263),
            .I(N__100260));
    Odrv4 I__24702 (
            .O(N__100260),
            .I(\c0.n14 ));
    CascadeMux I__24701 (
            .O(N__100257),
            .I(N__100250));
    InMux I__24700 (
            .O(N__100256),
            .I(N__100247));
    CascadeMux I__24699 (
            .O(N__100255),
            .I(N__100243));
    InMux I__24698 (
            .O(N__100254),
            .I(N__100240));
    InMux I__24697 (
            .O(N__100253),
            .I(N__100237));
    InMux I__24696 (
            .O(N__100250),
            .I(N__100234));
    LocalMux I__24695 (
            .O(N__100247),
            .I(N__100231));
    InMux I__24694 (
            .O(N__100246),
            .I(N__100228));
    InMux I__24693 (
            .O(N__100243),
            .I(N__100225));
    LocalMux I__24692 (
            .O(N__100240),
            .I(N__100222));
    LocalMux I__24691 (
            .O(N__100237),
            .I(N__100219));
    LocalMux I__24690 (
            .O(N__100234),
            .I(N__100216));
    Span4Mux_h I__24689 (
            .O(N__100231),
            .I(N__100213));
    LocalMux I__24688 (
            .O(N__100228),
            .I(N__100210));
    LocalMux I__24687 (
            .O(N__100225),
            .I(N__100207));
    Span4Mux_v I__24686 (
            .O(N__100222),
            .I(N__100203));
    Span4Mux_h I__24685 (
            .O(N__100219),
            .I(N__100198));
    Span4Mux_v I__24684 (
            .O(N__100216),
            .I(N__100198));
    Span4Mux_h I__24683 (
            .O(N__100213),
            .I(N__100195));
    Span4Mux_h I__24682 (
            .O(N__100210),
            .I(N__100190));
    Span4Mux_v I__24681 (
            .O(N__100207),
            .I(N__100190));
    InMux I__24680 (
            .O(N__100206),
            .I(N__100187));
    Span4Mux_h I__24679 (
            .O(N__100203),
            .I(N__100182));
    Span4Mux_v I__24678 (
            .O(N__100198),
            .I(N__100182));
    Span4Mux_v I__24677 (
            .O(N__100195),
            .I(N__100179));
    Span4Mux_h I__24676 (
            .O(N__100190),
            .I(N__100176));
    LocalMux I__24675 (
            .O(N__100187),
            .I(\c0.n15711 ));
    Odrv4 I__24674 (
            .O(N__100182),
            .I(\c0.n15711 ));
    Odrv4 I__24673 (
            .O(N__100179),
            .I(\c0.n15711 ));
    Odrv4 I__24672 (
            .O(N__100176),
            .I(\c0.n15711 ));
    InMux I__24671 (
            .O(N__100167),
            .I(N__100162));
    InMux I__24670 (
            .O(N__100166),
            .I(N__100156));
    InMux I__24669 (
            .O(N__100165),
            .I(N__100153));
    LocalMux I__24668 (
            .O(N__100162),
            .I(N__100150));
    InMux I__24667 (
            .O(N__100161),
            .I(N__100143));
    InMux I__24666 (
            .O(N__100160),
            .I(N__100143));
    InMux I__24665 (
            .O(N__100159),
            .I(N__100143));
    LocalMux I__24664 (
            .O(N__100156),
            .I(N__100140));
    LocalMux I__24663 (
            .O(N__100153),
            .I(N__100137));
    Span4Mux_h I__24662 (
            .O(N__100150),
            .I(N__100134));
    LocalMux I__24661 (
            .O(N__100143),
            .I(N__100131));
    Span4Mux_h I__24660 (
            .O(N__100140),
            .I(N__100128));
    Span4Mux_v I__24659 (
            .O(N__100137),
            .I(N__100123));
    Span4Mux_h I__24658 (
            .O(N__100134),
            .I(N__100123));
    Odrv12 I__24657 (
            .O(N__100131),
            .I(\c0.n17515 ));
    Odrv4 I__24656 (
            .O(N__100128),
            .I(\c0.n17515 ));
    Odrv4 I__24655 (
            .O(N__100123),
            .I(\c0.n17515 ));
    InMux I__24654 (
            .O(N__100116),
            .I(N__100113));
    LocalMux I__24653 (
            .O(N__100113),
            .I(N__100110));
    Span4Mux_h I__24652 (
            .O(N__100110),
            .I(N__100107));
    Odrv4 I__24651 (
            .O(N__100107),
            .I(\c0.n33548 ));
    InMux I__24650 (
            .O(N__100104),
            .I(N__100094));
    InMux I__24649 (
            .O(N__100103),
            .I(N__100094));
    InMux I__24648 (
            .O(N__100102),
            .I(N__100091));
    InMux I__24647 (
            .O(N__100101),
            .I(N__100088));
    InMux I__24646 (
            .O(N__100100),
            .I(N__100083));
    InMux I__24645 (
            .O(N__100099),
            .I(N__100083));
    LocalMux I__24644 (
            .O(N__100094),
            .I(N__100079));
    LocalMux I__24643 (
            .O(N__100091),
            .I(N__100071));
    LocalMux I__24642 (
            .O(N__100088),
            .I(N__100071));
    LocalMux I__24641 (
            .O(N__100083),
            .I(N__100071));
    CascadeMux I__24640 (
            .O(N__100082),
            .I(N__100067));
    Span4Mux_h I__24639 (
            .O(N__100079),
            .I(N__100064));
    InMux I__24638 (
            .O(N__100078),
            .I(N__100061));
    Span4Mux_v I__24637 (
            .O(N__100071),
            .I(N__100058));
    InMux I__24636 (
            .O(N__100070),
            .I(N__100055));
    InMux I__24635 (
            .O(N__100067),
            .I(N__100052));
    Odrv4 I__24634 (
            .O(N__100064),
            .I(\c0.n31468 ));
    LocalMux I__24633 (
            .O(N__100061),
            .I(\c0.n31468 ));
    Odrv4 I__24632 (
            .O(N__100058),
            .I(\c0.n31468 ));
    LocalMux I__24631 (
            .O(N__100055),
            .I(\c0.n31468 ));
    LocalMux I__24630 (
            .O(N__100052),
            .I(\c0.n31468 ));
    InMux I__24629 (
            .O(N__100041),
            .I(bfn_28_10_0_));
    InMux I__24628 (
            .O(N__100038),
            .I(N__100035));
    LocalMux I__24627 (
            .O(N__100035),
            .I(N__100031));
    CascadeMux I__24626 (
            .O(N__100034),
            .I(N__100028));
    Span4Mux_h I__24625 (
            .O(N__100031),
            .I(N__100024));
    InMux I__24624 (
            .O(N__100028),
            .I(N__100021));
    InMux I__24623 (
            .O(N__100027),
            .I(N__100018));
    Odrv4 I__24622 (
            .O(N__100024),
            .I(\quad_counter1.n1914 ));
    LocalMux I__24621 (
            .O(N__100021),
            .I(\quad_counter1.n1914 ));
    LocalMux I__24620 (
            .O(N__100018),
            .I(\quad_counter1.n1914 ));
    CascadeMux I__24619 (
            .O(N__100011),
            .I(N__100008));
    InMux I__24618 (
            .O(N__100008),
            .I(N__100005));
    LocalMux I__24617 (
            .O(N__100005),
            .I(N__100002));
    Span4Mux_h I__24616 (
            .O(N__100002),
            .I(N__99999));
    Odrv4 I__24615 (
            .O(N__99999),
            .I(\quad_counter1.n1981 ));
    CascadeMux I__24614 (
            .O(N__99996),
            .I(N__99991));
    CascadeMux I__24613 (
            .O(N__99995),
            .I(N__99987));
    CascadeMux I__24612 (
            .O(N__99994),
            .I(N__99983));
    InMux I__24611 (
            .O(N__99991),
            .I(N__99978));
    InMux I__24610 (
            .O(N__99990),
            .I(N__99975));
    InMux I__24609 (
            .O(N__99987),
            .I(N__99970));
    InMux I__24608 (
            .O(N__99986),
            .I(N__99970));
    InMux I__24607 (
            .O(N__99983),
            .I(N__99963));
    InMux I__24606 (
            .O(N__99982),
            .I(N__99963));
    InMux I__24605 (
            .O(N__99981),
            .I(N__99963));
    LocalMux I__24604 (
            .O(N__99978),
            .I(\quad_counter1.n1946 ));
    LocalMux I__24603 (
            .O(N__99975),
            .I(\quad_counter1.n1946 ));
    LocalMux I__24602 (
            .O(N__99970),
            .I(\quad_counter1.n1946 ));
    LocalMux I__24601 (
            .O(N__99963),
            .I(\quad_counter1.n1946 ));
    InMux I__24600 (
            .O(N__99954),
            .I(N__99949));
    InMux I__24599 (
            .O(N__99953),
            .I(N__99946));
    InMux I__24598 (
            .O(N__99952),
            .I(N__99943));
    LocalMux I__24597 (
            .O(N__99949),
            .I(\quad_counter1.n2014 ));
    LocalMux I__24596 (
            .O(N__99946),
            .I(\quad_counter1.n2014 ));
    LocalMux I__24595 (
            .O(N__99943),
            .I(\quad_counter1.n2014 ));
    InMux I__24594 (
            .O(N__99936),
            .I(N__99933));
    LocalMux I__24593 (
            .O(N__99933),
            .I(\quad_counter1.n2081 ));
    InMux I__24592 (
            .O(N__99930),
            .I(N__99926));
    InMux I__24591 (
            .O(N__99929),
            .I(N__99923));
    LocalMux I__24590 (
            .O(N__99926),
            .I(N__99917));
    LocalMux I__24589 (
            .O(N__99923),
            .I(N__99917));
    InMux I__24588 (
            .O(N__99922),
            .I(N__99913));
    Span4Mux_h I__24587 (
            .O(N__99917),
            .I(N__99910));
    InMux I__24586 (
            .O(N__99916),
            .I(N__99907));
    LocalMux I__24585 (
            .O(N__99913),
            .I(N__99904));
    Span4Mux_h I__24584 (
            .O(N__99910),
            .I(N__99901));
    LocalMux I__24583 (
            .O(N__99907),
            .I(\quad_counter1.millisecond_counter_23 ));
    Odrv12 I__24582 (
            .O(N__99904),
            .I(\quad_counter1.millisecond_counter_23 ));
    Odrv4 I__24581 (
            .O(N__99901),
            .I(\quad_counter1.millisecond_counter_23 ));
    InMux I__24580 (
            .O(N__99894),
            .I(N__99891));
    LocalMux I__24579 (
            .O(N__99891),
            .I(\quad_counter1.n2087 ));
    InMux I__24578 (
            .O(N__99888),
            .I(N__99883));
    InMux I__24577 (
            .O(N__99887),
            .I(N__99880));
    InMux I__24576 (
            .O(N__99886),
            .I(N__99877));
    LocalMux I__24575 (
            .O(N__99883),
            .I(\quad_counter1.n2119 ));
    LocalMux I__24574 (
            .O(N__99880),
            .I(\quad_counter1.n2119 ));
    LocalMux I__24573 (
            .O(N__99877),
            .I(\quad_counter1.n2119 ));
    CascadeMux I__24572 (
            .O(N__99870),
            .I(N__99865));
    InMux I__24571 (
            .O(N__99869),
            .I(N__99862));
    InMux I__24570 (
            .O(N__99868),
            .I(N__99859));
    InMux I__24569 (
            .O(N__99865),
            .I(N__99856));
    LocalMux I__24568 (
            .O(N__99862),
            .I(N__99853));
    LocalMux I__24567 (
            .O(N__99859),
            .I(\quad_counter1.n2017 ));
    LocalMux I__24566 (
            .O(N__99856),
            .I(\quad_counter1.n2017 ));
    Odrv4 I__24565 (
            .O(N__99853),
            .I(\quad_counter1.n2017 ));
    InMux I__24564 (
            .O(N__99846),
            .I(N__99843));
    LocalMux I__24563 (
            .O(N__99843),
            .I(\quad_counter1.n2084 ));
    CascadeMux I__24562 (
            .O(N__99840),
            .I(N__99836));
    CascadeMux I__24561 (
            .O(N__99839),
            .I(N__99833));
    InMux I__24560 (
            .O(N__99836),
            .I(N__99829));
    InMux I__24559 (
            .O(N__99833),
            .I(N__99826));
    InMux I__24558 (
            .O(N__99832),
            .I(N__99823));
    LocalMux I__24557 (
            .O(N__99829),
            .I(\quad_counter1.n2015 ));
    LocalMux I__24556 (
            .O(N__99826),
            .I(\quad_counter1.n2015 ));
    LocalMux I__24555 (
            .O(N__99823),
            .I(\quad_counter1.n2015 ));
    InMux I__24554 (
            .O(N__99816),
            .I(N__99813));
    LocalMux I__24553 (
            .O(N__99813),
            .I(\quad_counter1.n2082 ));
    InMux I__24552 (
            .O(N__99810),
            .I(N__99805));
    InMux I__24551 (
            .O(N__99809),
            .I(N__99802));
    InMux I__24550 (
            .O(N__99808),
            .I(N__99799));
    LocalMux I__24549 (
            .O(N__99805),
            .I(\quad_counter1.n2013 ));
    LocalMux I__24548 (
            .O(N__99802),
            .I(\quad_counter1.n2013 ));
    LocalMux I__24547 (
            .O(N__99799),
            .I(\quad_counter1.n2013 ));
    CascadeMux I__24546 (
            .O(N__99792),
            .I(N__99789));
    InMux I__24545 (
            .O(N__99789),
            .I(N__99786));
    LocalMux I__24544 (
            .O(N__99786),
            .I(N__99783));
    Odrv4 I__24543 (
            .O(N__99783),
            .I(\quad_counter1.n2080 ));
    InMux I__24542 (
            .O(N__99780),
            .I(N__99775));
    InMux I__24541 (
            .O(N__99779),
            .I(N__99772));
    InMux I__24540 (
            .O(N__99778),
            .I(N__99769));
    LocalMux I__24539 (
            .O(N__99775),
            .I(\quad_counter1.n2018 ));
    LocalMux I__24538 (
            .O(N__99772),
            .I(\quad_counter1.n2018 ));
    LocalMux I__24537 (
            .O(N__99769),
            .I(\quad_counter1.n2018 ));
    CascadeMux I__24536 (
            .O(N__99762),
            .I(N__99754));
    CascadeMux I__24535 (
            .O(N__99761),
            .I(N__99751));
    CascadeMux I__24534 (
            .O(N__99760),
            .I(N__99748));
    InMux I__24533 (
            .O(N__99759),
            .I(N__99741));
    InMux I__24532 (
            .O(N__99758),
            .I(N__99741));
    InMux I__24531 (
            .O(N__99757),
            .I(N__99738));
    InMux I__24530 (
            .O(N__99754),
            .I(N__99727));
    InMux I__24529 (
            .O(N__99751),
            .I(N__99727));
    InMux I__24528 (
            .O(N__99748),
            .I(N__99727));
    InMux I__24527 (
            .O(N__99747),
            .I(N__99727));
    InMux I__24526 (
            .O(N__99746),
            .I(N__99727));
    LocalMux I__24525 (
            .O(N__99741),
            .I(\quad_counter1.n2045 ));
    LocalMux I__24524 (
            .O(N__99738),
            .I(\quad_counter1.n2045 ));
    LocalMux I__24523 (
            .O(N__99727),
            .I(\quad_counter1.n2045 ));
    InMux I__24522 (
            .O(N__99720),
            .I(N__99717));
    LocalMux I__24521 (
            .O(N__99717),
            .I(N__99714));
    Odrv4 I__24520 (
            .O(N__99714),
            .I(\quad_counter1.n2085 ));
    InMux I__24519 (
            .O(N__99711),
            .I(N__99707));
    InMux I__24518 (
            .O(N__99710),
            .I(N__99704));
    LocalMux I__24517 (
            .O(N__99707),
            .I(\quad_counter1.n2117 ));
    LocalMux I__24516 (
            .O(N__99704),
            .I(\quad_counter1.n2117 ));
    CascadeMux I__24515 (
            .O(N__99699),
            .I(\quad_counter1.n2117_cascade_ ));
    InMux I__24514 (
            .O(N__99696),
            .I(N__99692));
    InMux I__24513 (
            .O(N__99695),
            .I(N__99689));
    LocalMux I__24512 (
            .O(N__99692),
            .I(N__99683));
    LocalMux I__24511 (
            .O(N__99689),
            .I(N__99683));
    InMux I__24510 (
            .O(N__99688),
            .I(N__99680));
    Odrv4 I__24509 (
            .O(N__99683),
            .I(\quad_counter1.n2114 ));
    LocalMux I__24508 (
            .O(N__99680),
            .I(\quad_counter1.n2114 ));
    InMux I__24507 (
            .O(N__99675),
            .I(bfn_28_9_0_));
    CascadeMux I__24506 (
            .O(N__99672),
            .I(N__99668));
    CascadeMux I__24505 (
            .O(N__99671),
            .I(N__99665));
    InMux I__24504 (
            .O(N__99668),
            .I(N__99662));
    InMux I__24503 (
            .O(N__99665),
            .I(N__99659));
    LocalMux I__24502 (
            .O(N__99662),
            .I(\quad_counter1.n2019 ));
    LocalMux I__24501 (
            .O(N__99659),
            .I(\quad_counter1.n2019 ));
    InMux I__24500 (
            .O(N__99654),
            .I(N__99651));
    LocalMux I__24499 (
            .O(N__99651),
            .I(\quad_counter1.n2086 ));
    InMux I__24498 (
            .O(N__99648),
            .I(\quad_counter1.n30472 ));
    InMux I__24497 (
            .O(N__99645),
            .I(\quad_counter1.n30473 ));
    InMux I__24496 (
            .O(N__99642),
            .I(\quad_counter1.n30474 ));
    CascadeMux I__24495 (
            .O(N__99639),
            .I(N__99635));
    InMux I__24494 (
            .O(N__99638),
            .I(N__99632));
    InMux I__24493 (
            .O(N__99635),
            .I(N__99629));
    LocalMux I__24492 (
            .O(N__99632),
            .I(\quad_counter1.n2016 ));
    LocalMux I__24491 (
            .O(N__99629),
            .I(\quad_counter1.n2016 ));
    InMux I__24490 (
            .O(N__99624),
            .I(N__99621));
    LocalMux I__24489 (
            .O(N__99621),
            .I(\quad_counter1.n2083 ));
    InMux I__24488 (
            .O(N__99618),
            .I(\quad_counter1.n30475 ));
    InMux I__24487 (
            .O(N__99615),
            .I(\quad_counter1.n30476 ));
    InMux I__24486 (
            .O(N__99612),
            .I(\quad_counter1.n30477 ));
    InMux I__24485 (
            .O(N__99609),
            .I(\quad_counter1.n30478 ));
    CascadeMux I__24484 (
            .O(N__99606),
            .I(N__99597));
    CascadeMux I__24483 (
            .O(N__99605),
            .I(N__99593));
    CascadeMux I__24482 (
            .O(N__99604),
            .I(N__99589));
    CascadeMux I__24481 (
            .O(N__99603),
            .I(N__99577));
    CascadeMux I__24480 (
            .O(N__99602),
            .I(N__99573));
    CascadeMux I__24479 (
            .O(N__99601),
            .I(N__99569));
    InMux I__24478 (
            .O(N__99600),
            .I(N__99543));
    InMux I__24477 (
            .O(N__99597),
            .I(N__99543));
    InMux I__24476 (
            .O(N__99596),
            .I(N__99543));
    InMux I__24475 (
            .O(N__99593),
            .I(N__99543));
    InMux I__24474 (
            .O(N__99592),
            .I(N__99543));
    InMux I__24473 (
            .O(N__99589),
            .I(N__99543));
    InMux I__24472 (
            .O(N__99588),
            .I(N__99543));
    InMux I__24471 (
            .O(N__99587),
            .I(N__99536));
    InMux I__24470 (
            .O(N__99586),
            .I(N__99536));
    InMux I__24469 (
            .O(N__99585),
            .I(N__99536));
    InMux I__24468 (
            .O(N__99584),
            .I(N__99527));
    InMux I__24467 (
            .O(N__99583),
            .I(N__99527));
    InMux I__24466 (
            .O(N__99582),
            .I(N__99527));
    InMux I__24465 (
            .O(N__99581),
            .I(N__99527));
    InMux I__24464 (
            .O(N__99580),
            .I(N__99512));
    InMux I__24463 (
            .O(N__99577),
            .I(N__99512));
    InMux I__24462 (
            .O(N__99576),
            .I(N__99512));
    InMux I__24461 (
            .O(N__99573),
            .I(N__99512));
    InMux I__24460 (
            .O(N__99572),
            .I(N__99512));
    InMux I__24459 (
            .O(N__99569),
            .I(N__99512));
    InMux I__24458 (
            .O(N__99568),
            .I(N__99512));
    CascadeMux I__24457 (
            .O(N__99567),
            .I(N__99505));
    CascadeMux I__24456 (
            .O(N__99566),
            .I(N__99501));
    CascadeMux I__24455 (
            .O(N__99565),
            .I(N__99497));
    CascadeMux I__24454 (
            .O(N__99564),
            .I(N__99485));
    CascadeMux I__24453 (
            .O(N__99563),
            .I(N__99481));
    CascadeMux I__24452 (
            .O(N__99562),
            .I(N__99477));
    InMux I__24451 (
            .O(N__99561),
            .I(N__99458));
    InMux I__24450 (
            .O(N__99560),
            .I(N__99458));
    InMux I__24449 (
            .O(N__99559),
            .I(N__99458));
    InMux I__24448 (
            .O(N__99558),
            .I(N__99458));
    LocalMux I__24447 (
            .O(N__99543),
            .I(N__99449));
    LocalMux I__24446 (
            .O(N__99536),
            .I(N__99449));
    LocalMux I__24445 (
            .O(N__99527),
            .I(N__99449));
    LocalMux I__24444 (
            .O(N__99512),
            .I(N__99449));
    InMux I__24443 (
            .O(N__99511),
            .I(N__99442));
    InMux I__24442 (
            .O(N__99510),
            .I(N__99442));
    InMux I__24441 (
            .O(N__99509),
            .I(N__99442));
    InMux I__24440 (
            .O(N__99508),
            .I(N__99427));
    InMux I__24439 (
            .O(N__99505),
            .I(N__99427));
    InMux I__24438 (
            .O(N__99504),
            .I(N__99427));
    InMux I__24437 (
            .O(N__99501),
            .I(N__99427));
    InMux I__24436 (
            .O(N__99500),
            .I(N__99427));
    InMux I__24435 (
            .O(N__99497),
            .I(N__99427));
    InMux I__24434 (
            .O(N__99496),
            .I(N__99427));
    InMux I__24433 (
            .O(N__99495),
            .I(N__99420));
    InMux I__24432 (
            .O(N__99494),
            .I(N__99420));
    InMux I__24431 (
            .O(N__99493),
            .I(N__99420));
    InMux I__24430 (
            .O(N__99492),
            .I(N__99411));
    InMux I__24429 (
            .O(N__99491),
            .I(N__99411));
    InMux I__24428 (
            .O(N__99490),
            .I(N__99411));
    InMux I__24427 (
            .O(N__99489),
            .I(N__99411));
    InMux I__24426 (
            .O(N__99488),
            .I(N__99396));
    InMux I__24425 (
            .O(N__99485),
            .I(N__99396));
    InMux I__24424 (
            .O(N__99484),
            .I(N__99396));
    InMux I__24423 (
            .O(N__99481),
            .I(N__99396));
    InMux I__24422 (
            .O(N__99480),
            .I(N__99396));
    InMux I__24421 (
            .O(N__99477),
            .I(N__99396));
    InMux I__24420 (
            .O(N__99476),
            .I(N__99396));
    CascadeMux I__24419 (
            .O(N__99475),
            .I(N__99392));
    CascadeMux I__24418 (
            .O(N__99474),
            .I(N__99388));
    CascadeMux I__24417 (
            .O(N__99473),
            .I(N__99384));
    CascadeMux I__24416 (
            .O(N__99472),
            .I(N__99379));
    CascadeMux I__24415 (
            .O(N__99471),
            .I(N__99375));
    CascadeMux I__24414 (
            .O(N__99470),
            .I(N__99371));
    CascadeMux I__24413 (
            .O(N__99469),
            .I(N__99359));
    CascadeMux I__24412 (
            .O(N__99468),
            .I(N__99355));
    CascadeMux I__24411 (
            .O(N__99467),
            .I(N__99351));
    LocalMux I__24410 (
            .O(N__99458),
            .I(N__99327));
    Span4Mux_v I__24409 (
            .O(N__99449),
            .I(N__99314));
    LocalMux I__24408 (
            .O(N__99442),
            .I(N__99314));
    LocalMux I__24407 (
            .O(N__99427),
            .I(N__99314));
    LocalMux I__24406 (
            .O(N__99420),
            .I(N__99314));
    LocalMux I__24405 (
            .O(N__99411),
            .I(N__99314));
    LocalMux I__24404 (
            .O(N__99396),
            .I(N__99314));
    InMux I__24403 (
            .O(N__99395),
            .I(N__99299));
    InMux I__24402 (
            .O(N__99392),
            .I(N__99299));
    InMux I__24401 (
            .O(N__99391),
            .I(N__99299));
    InMux I__24400 (
            .O(N__99388),
            .I(N__99299));
    InMux I__24399 (
            .O(N__99387),
            .I(N__99299));
    InMux I__24398 (
            .O(N__99384),
            .I(N__99299));
    InMux I__24397 (
            .O(N__99383),
            .I(N__99299));
    InMux I__24396 (
            .O(N__99382),
            .I(N__99284));
    InMux I__24395 (
            .O(N__99379),
            .I(N__99284));
    InMux I__24394 (
            .O(N__99378),
            .I(N__99284));
    InMux I__24393 (
            .O(N__99375),
            .I(N__99284));
    InMux I__24392 (
            .O(N__99374),
            .I(N__99284));
    InMux I__24391 (
            .O(N__99371),
            .I(N__99284));
    InMux I__24390 (
            .O(N__99370),
            .I(N__99284));
    InMux I__24389 (
            .O(N__99369),
            .I(N__99277));
    InMux I__24388 (
            .O(N__99368),
            .I(N__99277));
    InMux I__24387 (
            .O(N__99367),
            .I(N__99277));
    InMux I__24386 (
            .O(N__99366),
            .I(N__99268));
    InMux I__24385 (
            .O(N__99365),
            .I(N__99268));
    InMux I__24384 (
            .O(N__99364),
            .I(N__99268));
    InMux I__24383 (
            .O(N__99363),
            .I(N__99268));
    InMux I__24382 (
            .O(N__99362),
            .I(N__99253));
    InMux I__24381 (
            .O(N__99359),
            .I(N__99253));
    InMux I__24380 (
            .O(N__99358),
            .I(N__99253));
    InMux I__24379 (
            .O(N__99355),
            .I(N__99253));
    InMux I__24378 (
            .O(N__99354),
            .I(N__99253));
    InMux I__24377 (
            .O(N__99351),
            .I(N__99253));
    InMux I__24376 (
            .O(N__99350),
            .I(N__99253));
    CascadeMux I__24375 (
            .O(N__99349),
            .I(N__99249));
    CascadeMux I__24374 (
            .O(N__99348),
            .I(N__99245));
    CascadeMux I__24373 (
            .O(N__99347),
            .I(N__99241));
    CascadeMux I__24372 (
            .O(N__99346),
            .I(N__99236));
    CascadeMux I__24371 (
            .O(N__99345),
            .I(N__99232));
    CascadeMux I__24370 (
            .O(N__99344),
            .I(N__99228));
    CascadeMux I__24369 (
            .O(N__99343),
            .I(N__99216));
    CascadeMux I__24368 (
            .O(N__99342),
            .I(N__99212));
    CascadeMux I__24367 (
            .O(N__99341),
            .I(N__99208));
    CascadeMux I__24366 (
            .O(N__99340),
            .I(N__99197));
    CascadeMux I__24365 (
            .O(N__99339),
            .I(N__99193));
    CascadeMux I__24364 (
            .O(N__99338),
            .I(N__99189));
    CascadeMux I__24363 (
            .O(N__99337),
            .I(N__99184));
    CascadeMux I__24362 (
            .O(N__99336),
            .I(N__99180));
    CascadeMux I__24361 (
            .O(N__99335),
            .I(N__99176));
    CascadeMux I__24360 (
            .O(N__99334),
            .I(N__99171));
    CascadeMux I__24359 (
            .O(N__99333),
            .I(N__99167));
    CascadeMux I__24358 (
            .O(N__99332),
            .I(N__99163));
    CascadeMux I__24357 (
            .O(N__99331),
            .I(N__99158));
    IoInMux I__24356 (
            .O(N__99330),
            .I(N__99155));
    Span4Mux_v I__24355 (
            .O(N__99327),
            .I(N__99131));
    Span4Mux_v I__24354 (
            .O(N__99314),
            .I(N__99131));
    LocalMux I__24353 (
            .O(N__99299),
            .I(N__99131));
    LocalMux I__24352 (
            .O(N__99284),
            .I(N__99131));
    LocalMux I__24351 (
            .O(N__99277),
            .I(N__99131));
    LocalMux I__24350 (
            .O(N__99268),
            .I(N__99131));
    LocalMux I__24349 (
            .O(N__99253),
            .I(N__99131));
    InMux I__24348 (
            .O(N__99252),
            .I(N__99116));
    InMux I__24347 (
            .O(N__99249),
            .I(N__99116));
    InMux I__24346 (
            .O(N__99248),
            .I(N__99116));
    InMux I__24345 (
            .O(N__99245),
            .I(N__99116));
    InMux I__24344 (
            .O(N__99244),
            .I(N__99116));
    InMux I__24343 (
            .O(N__99241),
            .I(N__99116));
    InMux I__24342 (
            .O(N__99240),
            .I(N__99116));
    InMux I__24341 (
            .O(N__99239),
            .I(N__99101));
    InMux I__24340 (
            .O(N__99236),
            .I(N__99101));
    InMux I__24339 (
            .O(N__99235),
            .I(N__99101));
    InMux I__24338 (
            .O(N__99232),
            .I(N__99101));
    InMux I__24337 (
            .O(N__99231),
            .I(N__99101));
    InMux I__24336 (
            .O(N__99228),
            .I(N__99101));
    InMux I__24335 (
            .O(N__99227),
            .I(N__99101));
    InMux I__24334 (
            .O(N__99226),
            .I(N__99094));
    InMux I__24333 (
            .O(N__99225),
            .I(N__99094));
    InMux I__24332 (
            .O(N__99224),
            .I(N__99094));
    InMux I__24331 (
            .O(N__99223),
            .I(N__99085));
    InMux I__24330 (
            .O(N__99222),
            .I(N__99085));
    InMux I__24329 (
            .O(N__99221),
            .I(N__99085));
    InMux I__24328 (
            .O(N__99220),
            .I(N__99085));
    InMux I__24327 (
            .O(N__99219),
            .I(N__99070));
    InMux I__24326 (
            .O(N__99216),
            .I(N__99070));
    InMux I__24325 (
            .O(N__99215),
            .I(N__99070));
    InMux I__24324 (
            .O(N__99212),
            .I(N__99070));
    InMux I__24323 (
            .O(N__99211),
            .I(N__99070));
    InMux I__24322 (
            .O(N__99208),
            .I(N__99070));
    InMux I__24321 (
            .O(N__99207),
            .I(N__99070));
    CascadeMux I__24320 (
            .O(N__99206),
            .I(N__99059));
    CascadeMux I__24319 (
            .O(N__99205),
            .I(N__99055));
    CascadeMux I__24318 (
            .O(N__99204),
            .I(N__99051));
    CascadeMux I__24317 (
            .O(N__99203),
            .I(N__99039));
    CascadeMux I__24316 (
            .O(N__99202),
            .I(N__99035));
    CascadeMux I__24315 (
            .O(N__99201),
            .I(N__99031));
    InMux I__24314 (
            .O(N__99200),
            .I(N__99012));
    InMux I__24313 (
            .O(N__99197),
            .I(N__99012));
    InMux I__24312 (
            .O(N__99196),
            .I(N__99012));
    InMux I__24311 (
            .O(N__99193),
            .I(N__99012));
    InMux I__24310 (
            .O(N__99192),
            .I(N__99012));
    InMux I__24309 (
            .O(N__99189),
            .I(N__99012));
    InMux I__24308 (
            .O(N__99188),
            .I(N__99012));
    InMux I__24307 (
            .O(N__99187),
            .I(N__98997));
    InMux I__24306 (
            .O(N__99184),
            .I(N__98997));
    InMux I__24305 (
            .O(N__99183),
            .I(N__98997));
    InMux I__24304 (
            .O(N__99180),
            .I(N__98997));
    InMux I__24303 (
            .O(N__99179),
            .I(N__98997));
    InMux I__24302 (
            .O(N__99176),
            .I(N__98997));
    InMux I__24301 (
            .O(N__99175),
            .I(N__98997));
    InMux I__24300 (
            .O(N__99174),
            .I(N__98982));
    InMux I__24299 (
            .O(N__99171),
            .I(N__98982));
    InMux I__24298 (
            .O(N__99170),
            .I(N__98982));
    InMux I__24297 (
            .O(N__99167),
            .I(N__98982));
    InMux I__24296 (
            .O(N__99166),
            .I(N__98982));
    InMux I__24295 (
            .O(N__99163),
            .I(N__98982));
    InMux I__24294 (
            .O(N__99162),
            .I(N__98982));
    InMux I__24293 (
            .O(N__99161),
            .I(N__98967));
    InMux I__24292 (
            .O(N__99158),
            .I(N__98967));
    LocalMux I__24291 (
            .O(N__99155),
            .I(N__98962));
    CascadeMux I__24290 (
            .O(N__99154),
            .I(N__98958));
    CascadeMux I__24289 (
            .O(N__99153),
            .I(N__98954));
    CascadeMux I__24288 (
            .O(N__99152),
            .I(N__98950));
    InMux I__24287 (
            .O(N__99151),
            .I(N__98944));
    InMux I__24286 (
            .O(N__99150),
            .I(N__98944));
    InMux I__24285 (
            .O(N__99149),
            .I(N__98941));
    CascadeMux I__24284 (
            .O(N__99148),
            .I(N__98934));
    CascadeMux I__24283 (
            .O(N__99147),
            .I(N__98930));
    CascadeMux I__24282 (
            .O(N__99146),
            .I(N__98926));
    Span4Mux_v I__24281 (
            .O(N__99131),
            .I(N__98912));
    LocalMux I__24280 (
            .O(N__99116),
            .I(N__98912));
    LocalMux I__24279 (
            .O(N__99101),
            .I(N__98912));
    LocalMux I__24278 (
            .O(N__99094),
            .I(N__98912));
    LocalMux I__24277 (
            .O(N__99085),
            .I(N__98912));
    LocalMux I__24276 (
            .O(N__99070),
            .I(N__98912));
    InMux I__24275 (
            .O(N__99069),
            .I(N__98903));
    InMux I__24274 (
            .O(N__99068),
            .I(N__98903));
    InMux I__24273 (
            .O(N__99067),
            .I(N__98903));
    InMux I__24272 (
            .O(N__99066),
            .I(N__98903));
    InMux I__24271 (
            .O(N__99065),
            .I(N__98896));
    InMux I__24270 (
            .O(N__99064),
            .I(N__98896));
    InMux I__24269 (
            .O(N__99063),
            .I(N__98896));
    InMux I__24268 (
            .O(N__99062),
            .I(N__98881));
    InMux I__24267 (
            .O(N__99059),
            .I(N__98881));
    InMux I__24266 (
            .O(N__99058),
            .I(N__98881));
    InMux I__24265 (
            .O(N__99055),
            .I(N__98881));
    InMux I__24264 (
            .O(N__99054),
            .I(N__98881));
    InMux I__24263 (
            .O(N__99051),
            .I(N__98881));
    InMux I__24262 (
            .O(N__99050),
            .I(N__98881));
    InMux I__24261 (
            .O(N__99049),
            .I(N__98874));
    InMux I__24260 (
            .O(N__99048),
            .I(N__98874));
    InMux I__24259 (
            .O(N__99047),
            .I(N__98874));
    InMux I__24258 (
            .O(N__99046),
            .I(N__98865));
    InMux I__24257 (
            .O(N__99045),
            .I(N__98865));
    InMux I__24256 (
            .O(N__99044),
            .I(N__98865));
    InMux I__24255 (
            .O(N__99043),
            .I(N__98865));
    InMux I__24254 (
            .O(N__99042),
            .I(N__98850));
    InMux I__24253 (
            .O(N__99039),
            .I(N__98850));
    InMux I__24252 (
            .O(N__99038),
            .I(N__98850));
    InMux I__24251 (
            .O(N__99035),
            .I(N__98850));
    InMux I__24250 (
            .O(N__99034),
            .I(N__98850));
    InMux I__24249 (
            .O(N__99031),
            .I(N__98850));
    InMux I__24248 (
            .O(N__99030),
            .I(N__98850));
    CascadeMux I__24247 (
            .O(N__99029),
            .I(N__98846));
    CascadeMux I__24246 (
            .O(N__99028),
            .I(N__98842));
    CascadeMux I__24245 (
            .O(N__99027),
            .I(N__98838));
    LocalMux I__24244 (
            .O(N__99012),
            .I(N__98830));
    LocalMux I__24243 (
            .O(N__98997),
            .I(N__98830));
    LocalMux I__24242 (
            .O(N__98982),
            .I(N__98830));
    InMux I__24241 (
            .O(N__98981),
            .I(N__98821));
    InMux I__24240 (
            .O(N__98980),
            .I(N__98821));
    InMux I__24239 (
            .O(N__98979),
            .I(N__98821));
    InMux I__24238 (
            .O(N__98978),
            .I(N__98821));
    CascadeMux I__24237 (
            .O(N__98977),
            .I(N__98817));
    CascadeMux I__24236 (
            .O(N__98976),
            .I(N__98813));
    CascadeMux I__24235 (
            .O(N__98975),
            .I(N__98809));
    CascadeMux I__24234 (
            .O(N__98974),
            .I(N__98797));
    CascadeMux I__24233 (
            .O(N__98973),
            .I(N__98793));
    CascadeMux I__24232 (
            .O(N__98972),
            .I(N__98789));
    LocalMux I__24231 (
            .O(N__98967),
            .I(N__98785));
    InMux I__24230 (
            .O(N__98966),
            .I(N__98782));
    InMux I__24229 (
            .O(N__98965),
            .I(N__98774));
    Span4Mux_s2_v I__24228 (
            .O(N__98962),
            .I(N__98771));
    InMux I__24227 (
            .O(N__98961),
            .I(N__98756));
    InMux I__24226 (
            .O(N__98958),
            .I(N__98756));
    InMux I__24225 (
            .O(N__98957),
            .I(N__98756));
    InMux I__24224 (
            .O(N__98954),
            .I(N__98756));
    InMux I__24223 (
            .O(N__98953),
            .I(N__98756));
    InMux I__24222 (
            .O(N__98950),
            .I(N__98756));
    InMux I__24221 (
            .O(N__98949),
            .I(N__98756));
    LocalMux I__24220 (
            .O(N__98944),
            .I(N__98743));
    LocalMux I__24219 (
            .O(N__98941),
            .I(N__98743));
    InMux I__24218 (
            .O(N__98940),
            .I(N__98736));
    InMux I__24217 (
            .O(N__98939),
            .I(N__98736));
    InMux I__24216 (
            .O(N__98938),
            .I(N__98736));
    InMux I__24215 (
            .O(N__98937),
            .I(N__98721));
    InMux I__24214 (
            .O(N__98934),
            .I(N__98721));
    InMux I__24213 (
            .O(N__98933),
            .I(N__98721));
    InMux I__24212 (
            .O(N__98930),
            .I(N__98721));
    InMux I__24211 (
            .O(N__98929),
            .I(N__98721));
    InMux I__24210 (
            .O(N__98926),
            .I(N__98721));
    InMux I__24209 (
            .O(N__98925),
            .I(N__98721));
    Span4Mux_v I__24208 (
            .O(N__98912),
            .I(N__98716));
    LocalMux I__24207 (
            .O(N__98903),
            .I(N__98716));
    LocalMux I__24206 (
            .O(N__98896),
            .I(N__98705));
    LocalMux I__24205 (
            .O(N__98881),
            .I(N__98705));
    LocalMux I__24204 (
            .O(N__98874),
            .I(N__98705));
    LocalMux I__24203 (
            .O(N__98865),
            .I(N__98705));
    LocalMux I__24202 (
            .O(N__98850),
            .I(N__98705));
    InMux I__24201 (
            .O(N__98849),
            .I(N__98690));
    InMux I__24200 (
            .O(N__98846),
            .I(N__98690));
    InMux I__24199 (
            .O(N__98845),
            .I(N__98690));
    InMux I__24198 (
            .O(N__98842),
            .I(N__98690));
    InMux I__24197 (
            .O(N__98841),
            .I(N__98690));
    InMux I__24196 (
            .O(N__98838),
            .I(N__98690));
    InMux I__24195 (
            .O(N__98837),
            .I(N__98690));
    Span4Mux_s3_v I__24194 (
            .O(N__98830),
            .I(N__98685));
    LocalMux I__24193 (
            .O(N__98821),
            .I(N__98685));
    InMux I__24192 (
            .O(N__98820),
            .I(N__98670));
    InMux I__24191 (
            .O(N__98817),
            .I(N__98670));
    InMux I__24190 (
            .O(N__98816),
            .I(N__98670));
    InMux I__24189 (
            .O(N__98813),
            .I(N__98670));
    InMux I__24188 (
            .O(N__98812),
            .I(N__98670));
    InMux I__24187 (
            .O(N__98809),
            .I(N__98670));
    InMux I__24186 (
            .O(N__98808),
            .I(N__98670));
    InMux I__24185 (
            .O(N__98807),
            .I(N__98663));
    InMux I__24184 (
            .O(N__98806),
            .I(N__98663));
    InMux I__24183 (
            .O(N__98805),
            .I(N__98663));
    InMux I__24182 (
            .O(N__98804),
            .I(N__98654));
    InMux I__24181 (
            .O(N__98803),
            .I(N__98654));
    InMux I__24180 (
            .O(N__98802),
            .I(N__98654));
    InMux I__24179 (
            .O(N__98801),
            .I(N__98654));
    InMux I__24178 (
            .O(N__98800),
            .I(N__98639));
    InMux I__24177 (
            .O(N__98797),
            .I(N__98639));
    InMux I__24176 (
            .O(N__98796),
            .I(N__98639));
    InMux I__24175 (
            .O(N__98793),
            .I(N__98639));
    InMux I__24174 (
            .O(N__98792),
            .I(N__98639));
    InMux I__24173 (
            .O(N__98789),
            .I(N__98639));
    InMux I__24172 (
            .O(N__98788),
            .I(N__98639));
    Span4Mux_v I__24171 (
            .O(N__98785),
            .I(N__98636));
    LocalMux I__24170 (
            .O(N__98782),
            .I(N__98633));
    CascadeMux I__24169 (
            .O(N__98781),
            .I(N__98629));
    CascadeMux I__24168 (
            .O(N__98780),
            .I(N__98625));
    CascadeMux I__24167 (
            .O(N__98779),
            .I(N__98621));
    InMux I__24166 (
            .O(N__98778),
            .I(N__98617));
    InMux I__24165 (
            .O(N__98777),
            .I(N__98614));
    LocalMux I__24164 (
            .O(N__98774),
            .I(N__98611));
    Span4Mux_h I__24163 (
            .O(N__98771),
            .I(N__98606));
    LocalMux I__24162 (
            .O(N__98756),
            .I(N__98606));
    InMux I__24161 (
            .O(N__98755),
            .I(N__98599));
    InMux I__24160 (
            .O(N__98754),
            .I(N__98599));
    InMux I__24159 (
            .O(N__98753),
            .I(N__98599));
    InMux I__24158 (
            .O(N__98752),
            .I(N__98590));
    InMux I__24157 (
            .O(N__98751),
            .I(N__98590));
    InMux I__24156 (
            .O(N__98750),
            .I(N__98590));
    InMux I__24155 (
            .O(N__98749),
            .I(N__98590));
    CascadeMux I__24154 (
            .O(N__98748),
            .I(N__98586));
    Span12Mux_s7_v I__24153 (
            .O(N__98743),
            .I(N__98583));
    LocalMux I__24152 (
            .O(N__98736),
            .I(N__98578));
    LocalMux I__24151 (
            .O(N__98721),
            .I(N__98578));
    Span4Mux_v I__24150 (
            .O(N__98716),
            .I(N__98561));
    Span4Mux_v I__24149 (
            .O(N__98705),
            .I(N__98561));
    LocalMux I__24148 (
            .O(N__98690),
            .I(N__98561));
    Span4Mux_v I__24147 (
            .O(N__98685),
            .I(N__98561));
    LocalMux I__24146 (
            .O(N__98670),
            .I(N__98561));
    LocalMux I__24145 (
            .O(N__98663),
            .I(N__98561));
    LocalMux I__24144 (
            .O(N__98654),
            .I(N__98561));
    LocalMux I__24143 (
            .O(N__98639),
            .I(N__98561));
    Span4Mux_h I__24142 (
            .O(N__98636),
            .I(N__98556));
    Span4Mux_v I__24141 (
            .O(N__98633),
            .I(N__98556));
    InMux I__24140 (
            .O(N__98632),
            .I(N__98541));
    InMux I__24139 (
            .O(N__98629),
            .I(N__98541));
    InMux I__24138 (
            .O(N__98628),
            .I(N__98541));
    InMux I__24137 (
            .O(N__98625),
            .I(N__98541));
    InMux I__24136 (
            .O(N__98624),
            .I(N__98541));
    InMux I__24135 (
            .O(N__98621),
            .I(N__98541));
    InMux I__24134 (
            .O(N__98620),
            .I(N__98541));
    LocalMux I__24133 (
            .O(N__98617),
            .I(N__98538));
    LocalMux I__24132 (
            .O(N__98614),
            .I(N__98535));
    Span4Mux_h I__24131 (
            .O(N__98611),
            .I(N__98532));
    Span4Mux_v I__24130 (
            .O(N__98606),
            .I(N__98525));
    LocalMux I__24129 (
            .O(N__98599),
            .I(N__98525));
    LocalMux I__24128 (
            .O(N__98590),
            .I(N__98525));
    InMux I__24127 (
            .O(N__98589),
            .I(N__98522));
    InMux I__24126 (
            .O(N__98586),
            .I(N__98519));
    Span12Mux_h I__24125 (
            .O(N__98583),
            .I(N__98515));
    Span4Mux_v I__24124 (
            .O(N__98578),
            .I(N__98510));
    Span4Mux_v I__24123 (
            .O(N__98561),
            .I(N__98510));
    Sp12to4 I__24122 (
            .O(N__98556),
            .I(N__98505));
    LocalMux I__24121 (
            .O(N__98541),
            .I(N__98505));
    Span4Mux_v I__24120 (
            .O(N__98538),
            .I(N__98500));
    Span4Mux_v I__24119 (
            .O(N__98535),
            .I(N__98500));
    Span4Mux_h I__24118 (
            .O(N__98532),
            .I(N__98491));
    Span4Mux_h I__24117 (
            .O(N__98525),
            .I(N__98491));
    LocalMux I__24116 (
            .O(N__98522),
            .I(N__98491));
    LocalMux I__24115 (
            .O(N__98519),
            .I(N__98491));
    InMux I__24114 (
            .O(N__98518),
            .I(N__98488));
    Odrv12 I__24113 (
            .O(N__98515),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__24112 (
            .O(N__98510),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__24111 (
            .O(N__98505),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__24110 (
            .O(N__98500),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__24109 (
            .O(N__98491),
            .I(CONSTANT_ONE_NET));
    LocalMux I__24108 (
            .O(N__98488),
            .I(CONSTANT_ONE_NET));
    InMux I__24107 (
            .O(N__98475),
            .I(N__98472));
    LocalMux I__24106 (
            .O(N__98472),
            .I(N__98469));
    Span4Mux_h I__24105 (
            .O(N__98469),
            .I(N__98465));
    InMux I__24104 (
            .O(N__98468),
            .I(N__98462));
    Odrv4 I__24103 (
            .O(N__98465),
            .I(\quad_counter1.n2012 ));
    LocalMux I__24102 (
            .O(N__98462),
            .I(\quad_counter1.n2012 ));
    CascadeMux I__24101 (
            .O(N__98457),
            .I(N__98454));
    InMux I__24100 (
            .O(N__98454),
            .I(N__98451));
    LocalMux I__24099 (
            .O(N__98451),
            .I(N__98442));
    InMux I__24098 (
            .O(N__98450),
            .I(N__98437));
    InMux I__24097 (
            .O(N__98449),
            .I(N__98437));
    InMux I__24096 (
            .O(N__98448),
            .I(N__98434));
    InMux I__24095 (
            .O(N__98447),
            .I(N__98431));
    InMux I__24094 (
            .O(N__98446),
            .I(N__98426));
    InMux I__24093 (
            .O(N__98445),
            .I(N__98426));
    Span4Mux_h I__24092 (
            .O(N__98442),
            .I(N__98419));
    LocalMux I__24091 (
            .O(N__98437),
            .I(N__98419));
    LocalMux I__24090 (
            .O(N__98434),
            .I(N__98419));
    LocalMux I__24089 (
            .O(N__98431),
            .I(\c0.n31857 ));
    LocalMux I__24088 (
            .O(N__98426),
            .I(\c0.n31857 ));
    Odrv4 I__24087 (
            .O(N__98419),
            .I(\c0.n31857 ));
    CascadeMux I__24086 (
            .O(N__98412),
            .I(\c0.n35280_cascade_ ));
    InMux I__24085 (
            .O(N__98409),
            .I(N__98406));
    LocalMux I__24084 (
            .O(N__98406),
            .I(N__98403));
    Span4Mux_h I__24083 (
            .O(N__98403),
            .I(N__98400));
    Odrv4 I__24082 (
            .O(N__98400),
            .I(\c0.n31461 ));
    CascadeMux I__24081 (
            .O(N__98397),
            .I(N__98394));
    InMux I__24080 (
            .O(N__98394),
            .I(N__98391));
    LocalMux I__24079 (
            .O(N__98391),
            .I(N__98387));
    InMux I__24078 (
            .O(N__98390),
            .I(N__98384));
    Span4Mux_h I__24077 (
            .O(N__98387),
            .I(N__98381));
    LocalMux I__24076 (
            .O(N__98384),
            .I(N__98378));
    Odrv4 I__24075 (
            .O(N__98381),
            .I(\c0.n32337 ));
    Odrv12 I__24074 (
            .O(N__98378),
            .I(\c0.n32337 ));
    CascadeMux I__24073 (
            .O(N__98373),
            .I(\c0.n31461_cascade_ ));
    InMux I__24072 (
            .O(N__98370),
            .I(N__98366));
    InMux I__24071 (
            .O(N__98369),
            .I(N__98363));
    LocalMux I__24070 (
            .O(N__98366),
            .I(\c0.n33839 ));
    LocalMux I__24069 (
            .O(N__98363),
            .I(\c0.n33839 ));
    InMux I__24068 (
            .O(N__98358),
            .I(N__98355));
    LocalMux I__24067 (
            .O(N__98355),
            .I(\c0.n8_adj_4529 ));
    InMux I__24066 (
            .O(N__98352),
            .I(N__98346));
    InMux I__24065 (
            .O(N__98351),
            .I(N__98346));
    LocalMux I__24064 (
            .O(N__98346),
            .I(N__98339));
    InMux I__24063 (
            .O(N__98345),
            .I(N__98336));
    InMux I__24062 (
            .O(N__98344),
            .I(N__98330));
    InMux I__24061 (
            .O(N__98343),
            .I(N__98330));
    InMux I__24060 (
            .O(N__98342),
            .I(N__98327));
    Span4Mux_h I__24059 (
            .O(N__98339),
            .I(N__98322));
    LocalMux I__24058 (
            .O(N__98336),
            .I(N__98322));
    InMux I__24057 (
            .O(N__98335),
            .I(N__98319));
    LocalMux I__24056 (
            .O(N__98330),
            .I(N__98314));
    LocalMux I__24055 (
            .O(N__98327),
            .I(N__98314));
    Span4Mux_h I__24054 (
            .O(N__98322),
            .I(N__98311));
    LocalMux I__24053 (
            .O(N__98319),
            .I(N__98308));
    Span12Mux_h I__24052 (
            .O(N__98314),
            .I(N__98305));
    Odrv4 I__24051 (
            .O(N__98311),
            .I(\c0.n31423 ));
    Odrv4 I__24050 (
            .O(N__98308),
            .I(\c0.n31423 ));
    Odrv12 I__24049 (
            .O(N__98305),
            .I(\c0.n31423 ));
    InMux I__24048 (
            .O(N__98298),
            .I(N__98295));
    LocalMux I__24047 (
            .O(N__98295),
            .I(N__98292));
    Span4Mux_h I__24046 (
            .O(N__98292),
            .I(N__98288));
    InMux I__24045 (
            .O(N__98291),
            .I(N__98285));
    Odrv4 I__24044 (
            .O(N__98288),
            .I(\c0.n31387 ));
    LocalMux I__24043 (
            .O(N__98285),
            .I(\c0.n31387 ));
    CascadeMux I__24042 (
            .O(N__98280),
            .I(N__98277));
    InMux I__24041 (
            .O(N__98277),
            .I(N__98268));
    InMux I__24040 (
            .O(N__98276),
            .I(N__98268));
    InMux I__24039 (
            .O(N__98275),
            .I(N__98265));
    CascadeMux I__24038 (
            .O(N__98274),
            .I(N__98262));
    InMux I__24037 (
            .O(N__98273),
            .I(N__98258));
    LocalMux I__24036 (
            .O(N__98268),
            .I(N__98253));
    LocalMux I__24035 (
            .O(N__98265),
            .I(N__98253));
    InMux I__24034 (
            .O(N__98262),
            .I(N__98248));
    InMux I__24033 (
            .O(N__98261),
            .I(N__98248));
    LocalMux I__24032 (
            .O(N__98258),
            .I(N__98244));
    Span4Mux_v I__24031 (
            .O(N__98253),
            .I(N__98238));
    LocalMux I__24030 (
            .O(N__98248),
            .I(N__98238));
    InMux I__24029 (
            .O(N__98247),
            .I(N__98235));
    Span4Mux_h I__24028 (
            .O(N__98244),
            .I(N__98232));
    InMux I__24027 (
            .O(N__98243),
            .I(N__98229));
    Span4Mux_h I__24026 (
            .O(N__98238),
            .I(N__98222));
    LocalMux I__24025 (
            .O(N__98235),
            .I(N__98222));
    Span4Mux_h I__24024 (
            .O(N__98232),
            .I(N__98222));
    LocalMux I__24023 (
            .O(N__98229),
            .I(\c0.n32290 ));
    Odrv4 I__24022 (
            .O(N__98222),
            .I(\c0.n32290 ));
    CascadeMux I__24021 (
            .O(N__98217),
            .I(N__98214));
    InMux I__24020 (
            .O(N__98214),
            .I(N__98211));
    LocalMux I__24019 (
            .O(N__98211),
            .I(N__98208));
    Odrv12 I__24018 (
            .O(N__98208),
            .I(\c0.n33670 ));
    InMux I__24017 (
            .O(N__98205),
            .I(N__98202));
    LocalMux I__24016 (
            .O(N__98202),
            .I(N__98199));
    Span4Mux_h I__24015 (
            .O(N__98199),
            .I(N__98196));
    Span4Mux_v I__24014 (
            .O(N__98196),
            .I(N__98193));
    Odrv4 I__24013 (
            .O(N__98193),
            .I(\c0.n31446 ));
    CascadeMux I__24012 (
            .O(N__98190),
            .I(\c0.n33670_cascade_ ));
    InMux I__24011 (
            .O(N__98187),
            .I(N__98184));
    LocalMux I__24010 (
            .O(N__98184),
            .I(N__98180));
    InMux I__24009 (
            .O(N__98183),
            .I(N__98177));
    Odrv4 I__24008 (
            .O(N__98180),
            .I(\c0.n15744 ));
    LocalMux I__24007 (
            .O(N__98177),
            .I(\c0.n15744 ));
    CascadeMux I__24006 (
            .O(N__98172),
            .I(\c0.n14_adj_4543_cascade_ ));
    InMux I__24005 (
            .O(N__98169),
            .I(N__98165));
    InMux I__24004 (
            .O(N__98168),
            .I(N__98162));
    LocalMux I__24003 (
            .O(N__98165),
            .I(N__98159));
    LocalMux I__24002 (
            .O(N__98162),
            .I(N__98155));
    Span4Mux_h I__24001 (
            .O(N__98159),
            .I(N__98152));
    CascadeMux I__24000 (
            .O(N__98158),
            .I(N__98149));
    Span4Mux_h I__23999 (
            .O(N__98155),
            .I(N__98144));
    Span4Mux_v I__23998 (
            .O(N__98152),
            .I(N__98144));
    InMux I__23997 (
            .O(N__98149),
            .I(N__98141));
    Odrv4 I__23996 (
            .O(N__98144),
            .I(\c0.n18232 ));
    LocalMux I__23995 (
            .O(N__98141),
            .I(\c0.n18232 ));
    InMux I__23994 (
            .O(N__98136),
            .I(N__98133));
    LocalMux I__23993 (
            .O(N__98133),
            .I(N__98129));
    InMux I__23992 (
            .O(N__98132),
            .I(N__98126));
    Odrv12 I__23991 (
            .O(N__98129),
            .I(\c0.n32071 ));
    LocalMux I__23990 (
            .O(N__98126),
            .I(\c0.n32071 ));
    InMux I__23989 (
            .O(N__98121),
            .I(N__98112));
    InMux I__23988 (
            .O(N__98120),
            .I(N__98112));
    InMux I__23987 (
            .O(N__98119),
            .I(N__98105));
    InMux I__23986 (
            .O(N__98118),
            .I(N__98105));
    InMux I__23985 (
            .O(N__98117),
            .I(N__98102));
    LocalMux I__23984 (
            .O(N__98112),
            .I(N__98099));
    InMux I__23983 (
            .O(N__98111),
            .I(N__98096));
    InMux I__23982 (
            .O(N__98110),
            .I(N__98093));
    LocalMux I__23981 (
            .O(N__98105),
            .I(N__98088));
    LocalMux I__23980 (
            .O(N__98102),
            .I(N__98088));
    Span4Mux_v I__23979 (
            .O(N__98099),
            .I(N__98084));
    LocalMux I__23978 (
            .O(N__98096),
            .I(N__98081));
    LocalMux I__23977 (
            .O(N__98093),
            .I(N__98076));
    Span4Mux_h I__23976 (
            .O(N__98088),
            .I(N__98076));
    InMux I__23975 (
            .O(N__98087),
            .I(N__98073));
    Odrv4 I__23974 (
            .O(N__98084),
            .I(\c0.n31878 ));
    Odrv12 I__23973 (
            .O(N__98081),
            .I(\c0.n31878 ));
    Odrv4 I__23972 (
            .O(N__98076),
            .I(\c0.n31878 ));
    LocalMux I__23971 (
            .O(N__98073),
            .I(\c0.n31878 ));
    InMux I__23970 (
            .O(N__98064),
            .I(N__98061));
    LocalMux I__23969 (
            .O(N__98061),
            .I(N__98058));
    Span4Mux_v I__23968 (
            .O(N__98058),
            .I(N__98055));
    Span4Mux_h I__23967 (
            .O(N__98055),
            .I(N__98052));
    Odrv4 I__23966 (
            .O(N__98052),
            .I(\c0.n33687 ));
    InMux I__23965 (
            .O(N__98049),
            .I(N__98046));
    LocalMux I__23964 (
            .O(N__98046),
            .I(\c0.n19_adj_4550 ));
    CascadeMux I__23963 (
            .O(N__98043),
            .I(N__98039));
    InMux I__23962 (
            .O(N__98042),
            .I(N__98035));
    InMux I__23961 (
            .O(N__98039),
            .I(N__98030));
    CascadeMux I__23960 (
            .O(N__98038),
            .I(N__98027));
    LocalMux I__23959 (
            .O(N__98035),
            .I(N__98023));
    InMux I__23958 (
            .O(N__98034),
            .I(N__98020));
    InMux I__23957 (
            .O(N__98033),
            .I(N__98017));
    LocalMux I__23956 (
            .O(N__98030),
            .I(N__98014));
    InMux I__23955 (
            .O(N__98027),
            .I(N__98009));
    InMux I__23954 (
            .O(N__98026),
            .I(N__98009));
    Span4Mux_h I__23953 (
            .O(N__98023),
            .I(N__98006));
    LocalMux I__23952 (
            .O(N__98020),
            .I(N__98003));
    LocalMux I__23951 (
            .O(N__98017),
            .I(N__98000));
    Span4Mux_v I__23950 (
            .O(N__98014),
            .I(N__97995));
    LocalMux I__23949 (
            .O(N__98009),
            .I(N__97995));
    Span4Mux_h I__23948 (
            .O(N__98006),
            .I(N__97992));
    Span4Mux_v I__23947 (
            .O(N__98003),
            .I(N__97987));
    Span4Mux_v I__23946 (
            .O(N__98000),
            .I(N__97987));
    Odrv4 I__23945 (
            .O(N__97995),
            .I(\c0.n33746 ));
    Odrv4 I__23944 (
            .O(N__97992),
            .I(\c0.n33746 ));
    Odrv4 I__23943 (
            .O(N__97987),
            .I(\c0.n33746 ));
    InMux I__23942 (
            .O(N__97980),
            .I(N__97977));
    LocalMux I__23941 (
            .O(N__97977),
            .I(N__97971));
    InMux I__23940 (
            .O(N__97976),
            .I(N__97968));
    InMux I__23939 (
            .O(N__97975),
            .I(N__97963));
    InMux I__23938 (
            .O(N__97974),
            .I(N__97963));
    Span4Mux_v I__23937 (
            .O(N__97971),
            .I(N__97958));
    LocalMux I__23936 (
            .O(N__97968),
            .I(N__97955));
    LocalMux I__23935 (
            .O(N__97963),
            .I(N__97952));
    CascadeMux I__23934 (
            .O(N__97962),
            .I(N__97948));
    CascadeMux I__23933 (
            .O(N__97961),
            .I(N__97945));
    Span4Mux_v I__23932 (
            .O(N__97958),
            .I(N__97942));
    Span4Mux_v I__23931 (
            .O(N__97955),
            .I(N__97937));
    Span4Mux_h I__23930 (
            .O(N__97952),
            .I(N__97937));
    InMux I__23929 (
            .O(N__97951),
            .I(N__97932));
    InMux I__23928 (
            .O(N__97948),
            .I(N__97932));
    InMux I__23927 (
            .O(N__97945),
            .I(N__97929));
    Sp12to4 I__23926 (
            .O(N__97942),
            .I(N__97926));
    Span4Mux_h I__23925 (
            .O(N__97937),
            .I(N__97923));
    LocalMux I__23924 (
            .O(N__97932),
            .I(encoder1_position_7));
    LocalMux I__23923 (
            .O(N__97929),
            .I(encoder1_position_7));
    Odrv12 I__23922 (
            .O(N__97926),
            .I(encoder1_position_7));
    Odrv4 I__23921 (
            .O(N__97923),
            .I(encoder1_position_7));
    InMux I__23920 (
            .O(N__97914),
            .I(N__97911));
    LocalMux I__23919 (
            .O(N__97911),
            .I(\c0.n10_adj_4542 ));
    InMux I__23918 (
            .O(N__97908),
            .I(N__97905));
    LocalMux I__23917 (
            .O(N__97905),
            .I(N__97902));
    Span4Mux_v I__23916 (
            .O(N__97902),
            .I(N__97897));
    InMux I__23915 (
            .O(N__97901),
            .I(N__97892));
    InMux I__23914 (
            .O(N__97900),
            .I(N__97892));
    Span4Mux_h I__23913 (
            .O(N__97897),
            .I(N__97887));
    LocalMux I__23912 (
            .O(N__97892),
            .I(N__97887));
    Span4Mux_v I__23911 (
            .O(N__97887),
            .I(N__97884));
    Odrv4 I__23910 (
            .O(N__97884),
            .I(\c0.n35426 ));
    InMux I__23909 (
            .O(N__97881),
            .I(N__97877));
    CascadeMux I__23908 (
            .O(N__97880),
            .I(N__97871));
    LocalMux I__23907 (
            .O(N__97877),
            .I(N__97868));
    InMux I__23906 (
            .O(N__97876),
            .I(N__97865));
    InMux I__23905 (
            .O(N__97875),
            .I(N__97858));
    InMux I__23904 (
            .O(N__97874),
            .I(N__97858));
    InMux I__23903 (
            .O(N__97871),
            .I(N__97858));
    Span4Mux_v I__23902 (
            .O(N__97868),
            .I(N__97853));
    LocalMux I__23901 (
            .O(N__97865),
            .I(N__97853));
    LocalMux I__23900 (
            .O(N__97858),
            .I(N__97850));
    Span4Mux_v I__23899 (
            .O(N__97853),
            .I(N__97845));
    Span4Mux_v I__23898 (
            .O(N__97850),
            .I(N__97845));
    Span4Mux_v I__23897 (
            .O(N__97845),
            .I(N__97840));
    InMux I__23896 (
            .O(N__97844),
            .I(N__97835));
    InMux I__23895 (
            .O(N__97843),
            .I(N__97835));
    Span4Mux_h I__23894 (
            .O(N__97840),
            .I(N__97832));
    LocalMux I__23893 (
            .O(N__97835),
            .I(data_out_frame_29__7__N_1426));
    Odrv4 I__23892 (
            .O(N__97832),
            .I(data_out_frame_29__7__N_1426));
    CascadeMux I__23891 (
            .O(N__97827),
            .I(\c0.n16_cascade_ ));
    InMux I__23890 (
            .O(N__97824),
            .I(N__97821));
    LocalMux I__23889 (
            .O(N__97821),
            .I(N__97818));
    Span4Mux_h I__23888 (
            .O(N__97818),
            .I(N__97815));
    Span4Mux_h I__23887 (
            .O(N__97815),
            .I(N__97812));
    Odrv4 I__23886 (
            .O(N__97812),
            .I(\c0.data_out_frame_28_7 ));
    InMux I__23885 (
            .O(N__97809),
            .I(N__97806));
    LocalMux I__23884 (
            .O(N__97806),
            .I(N__97798));
    ClkMux I__23883 (
            .O(N__97805),
            .I(N__97002));
    ClkMux I__23882 (
            .O(N__97804),
            .I(N__97002));
    ClkMux I__23881 (
            .O(N__97803),
            .I(N__97002));
    ClkMux I__23880 (
            .O(N__97802),
            .I(N__97002));
    ClkMux I__23879 (
            .O(N__97801),
            .I(N__97002));
    Glb2LocalMux I__23878 (
            .O(N__97798),
            .I(N__97002));
    ClkMux I__23877 (
            .O(N__97797),
            .I(N__97002));
    ClkMux I__23876 (
            .O(N__97796),
            .I(N__97002));
    ClkMux I__23875 (
            .O(N__97795),
            .I(N__97002));
    ClkMux I__23874 (
            .O(N__97794),
            .I(N__97002));
    ClkMux I__23873 (
            .O(N__97793),
            .I(N__97002));
    ClkMux I__23872 (
            .O(N__97792),
            .I(N__97002));
    ClkMux I__23871 (
            .O(N__97791),
            .I(N__97002));
    ClkMux I__23870 (
            .O(N__97790),
            .I(N__97002));
    ClkMux I__23869 (
            .O(N__97789),
            .I(N__97002));
    ClkMux I__23868 (
            .O(N__97788),
            .I(N__97002));
    ClkMux I__23867 (
            .O(N__97787),
            .I(N__97002));
    ClkMux I__23866 (
            .O(N__97786),
            .I(N__97002));
    ClkMux I__23865 (
            .O(N__97785),
            .I(N__97002));
    ClkMux I__23864 (
            .O(N__97784),
            .I(N__97002));
    ClkMux I__23863 (
            .O(N__97783),
            .I(N__97002));
    ClkMux I__23862 (
            .O(N__97782),
            .I(N__97002));
    ClkMux I__23861 (
            .O(N__97781),
            .I(N__97002));
    ClkMux I__23860 (
            .O(N__97780),
            .I(N__97002));
    ClkMux I__23859 (
            .O(N__97779),
            .I(N__97002));
    ClkMux I__23858 (
            .O(N__97778),
            .I(N__97002));
    ClkMux I__23857 (
            .O(N__97777),
            .I(N__97002));
    ClkMux I__23856 (
            .O(N__97776),
            .I(N__97002));
    ClkMux I__23855 (
            .O(N__97775),
            .I(N__97002));
    ClkMux I__23854 (
            .O(N__97774),
            .I(N__97002));
    ClkMux I__23853 (
            .O(N__97773),
            .I(N__97002));
    ClkMux I__23852 (
            .O(N__97772),
            .I(N__97002));
    ClkMux I__23851 (
            .O(N__97771),
            .I(N__97002));
    ClkMux I__23850 (
            .O(N__97770),
            .I(N__97002));
    ClkMux I__23849 (
            .O(N__97769),
            .I(N__97002));
    ClkMux I__23848 (
            .O(N__97768),
            .I(N__97002));
    ClkMux I__23847 (
            .O(N__97767),
            .I(N__97002));
    ClkMux I__23846 (
            .O(N__97766),
            .I(N__97002));
    ClkMux I__23845 (
            .O(N__97765),
            .I(N__97002));
    ClkMux I__23844 (
            .O(N__97764),
            .I(N__97002));
    ClkMux I__23843 (
            .O(N__97763),
            .I(N__97002));
    ClkMux I__23842 (
            .O(N__97762),
            .I(N__97002));
    ClkMux I__23841 (
            .O(N__97761),
            .I(N__97002));
    ClkMux I__23840 (
            .O(N__97760),
            .I(N__97002));
    ClkMux I__23839 (
            .O(N__97759),
            .I(N__97002));
    ClkMux I__23838 (
            .O(N__97758),
            .I(N__97002));
    ClkMux I__23837 (
            .O(N__97757),
            .I(N__97002));
    ClkMux I__23836 (
            .O(N__97756),
            .I(N__97002));
    ClkMux I__23835 (
            .O(N__97755),
            .I(N__97002));
    ClkMux I__23834 (
            .O(N__97754),
            .I(N__97002));
    ClkMux I__23833 (
            .O(N__97753),
            .I(N__97002));
    ClkMux I__23832 (
            .O(N__97752),
            .I(N__97002));
    ClkMux I__23831 (
            .O(N__97751),
            .I(N__97002));
    ClkMux I__23830 (
            .O(N__97750),
            .I(N__97002));
    ClkMux I__23829 (
            .O(N__97749),
            .I(N__97002));
    ClkMux I__23828 (
            .O(N__97748),
            .I(N__97002));
    ClkMux I__23827 (
            .O(N__97747),
            .I(N__97002));
    ClkMux I__23826 (
            .O(N__97746),
            .I(N__97002));
    ClkMux I__23825 (
            .O(N__97745),
            .I(N__97002));
    ClkMux I__23824 (
            .O(N__97744),
            .I(N__97002));
    ClkMux I__23823 (
            .O(N__97743),
            .I(N__97002));
    ClkMux I__23822 (
            .O(N__97742),
            .I(N__97002));
    ClkMux I__23821 (
            .O(N__97741),
            .I(N__97002));
    ClkMux I__23820 (
            .O(N__97740),
            .I(N__97002));
    ClkMux I__23819 (
            .O(N__97739),
            .I(N__97002));
    ClkMux I__23818 (
            .O(N__97738),
            .I(N__97002));
    ClkMux I__23817 (
            .O(N__97737),
            .I(N__97002));
    ClkMux I__23816 (
            .O(N__97736),
            .I(N__97002));
    ClkMux I__23815 (
            .O(N__97735),
            .I(N__97002));
    ClkMux I__23814 (
            .O(N__97734),
            .I(N__97002));
    ClkMux I__23813 (
            .O(N__97733),
            .I(N__97002));
    ClkMux I__23812 (
            .O(N__97732),
            .I(N__97002));
    ClkMux I__23811 (
            .O(N__97731),
            .I(N__97002));
    ClkMux I__23810 (
            .O(N__97730),
            .I(N__97002));
    ClkMux I__23809 (
            .O(N__97729),
            .I(N__97002));
    ClkMux I__23808 (
            .O(N__97728),
            .I(N__97002));
    ClkMux I__23807 (
            .O(N__97727),
            .I(N__97002));
    ClkMux I__23806 (
            .O(N__97726),
            .I(N__97002));
    ClkMux I__23805 (
            .O(N__97725),
            .I(N__97002));
    ClkMux I__23804 (
            .O(N__97724),
            .I(N__97002));
    ClkMux I__23803 (
            .O(N__97723),
            .I(N__97002));
    ClkMux I__23802 (
            .O(N__97722),
            .I(N__97002));
    ClkMux I__23801 (
            .O(N__97721),
            .I(N__97002));
    ClkMux I__23800 (
            .O(N__97720),
            .I(N__97002));
    ClkMux I__23799 (
            .O(N__97719),
            .I(N__97002));
    ClkMux I__23798 (
            .O(N__97718),
            .I(N__97002));
    ClkMux I__23797 (
            .O(N__97717),
            .I(N__97002));
    ClkMux I__23796 (
            .O(N__97716),
            .I(N__97002));
    ClkMux I__23795 (
            .O(N__97715),
            .I(N__97002));
    ClkMux I__23794 (
            .O(N__97714),
            .I(N__97002));
    ClkMux I__23793 (
            .O(N__97713),
            .I(N__97002));
    ClkMux I__23792 (
            .O(N__97712),
            .I(N__97002));
    ClkMux I__23791 (
            .O(N__97711),
            .I(N__97002));
    ClkMux I__23790 (
            .O(N__97710),
            .I(N__97002));
    ClkMux I__23789 (
            .O(N__97709),
            .I(N__97002));
    ClkMux I__23788 (
            .O(N__97708),
            .I(N__97002));
    ClkMux I__23787 (
            .O(N__97707),
            .I(N__97002));
    ClkMux I__23786 (
            .O(N__97706),
            .I(N__97002));
    ClkMux I__23785 (
            .O(N__97705),
            .I(N__97002));
    ClkMux I__23784 (
            .O(N__97704),
            .I(N__97002));
    ClkMux I__23783 (
            .O(N__97703),
            .I(N__97002));
    ClkMux I__23782 (
            .O(N__97702),
            .I(N__97002));
    ClkMux I__23781 (
            .O(N__97701),
            .I(N__97002));
    ClkMux I__23780 (
            .O(N__97700),
            .I(N__97002));
    ClkMux I__23779 (
            .O(N__97699),
            .I(N__97002));
    ClkMux I__23778 (
            .O(N__97698),
            .I(N__97002));
    ClkMux I__23777 (
            .O(N__97697),
            .I(N__97002));
    ClkMux I__23776 (
            .O(N__97696),
            .I(N__97002));
    ClkMux I__23775 (
            .O(N__97695),
            .I(N__97002));
    ClkMux I__23774 (
            .O(N__97694),
            .I(N__97002));
    ClkMux I__23773 (
            .O(N__97693),
            .I(N__97002));
    ClkMux I__23772 (
            .O(N__97692),
            .I(N__97002));
    ClkMux I__23771 (
            .O(N__97691),
            .I(N__97002));
    ClkMux I__23770 (
            .O(N__97690),
            .I(N__97002));
    ClkMux I__23769 (
            .O(N__97689),
            .I(N__97002));
    ClkMux I__23768 (
            .O(N__97688),
            .I(N__97002));
    ClkMux I__23767 (
            .O(N__97687),
            .I(N__97002));
    ClkMux I__23766 (
            .O(N__97686),
            .I(N__97002));
    ClkMux I__23765 (
            .O(N__97685),
            .I(N__97002));
    ClkMux I__23764 (
            .O(N__97684),
            .I(N__97002));
    ClkMux I__23763 (
            .O(N__97683),
            .I(N__97002));
    ClkMux I__23762 (
            .O(N__97682),
            .I(N__97002));
    ClkMux I__23761 (
            .O(N__97681),
            .I(N__97002));
    ClkMux I__23760 (
            .O(N__97680),
            .I(N__97002));
    ClkMux I__23759 (
            .O(N__97679),
            .I(N__97002));
    ClkMux I__23758 (
            .O(N__97678),
            .I(N__97002));
    ClkMux I__23757 (
            .O(N__97677),
            .I(N__97002));
    ClkMux I__23756 (
            .O(N__97676),
            .I(N__97002));
    ClkMux I__23755 (
            .O(N__97675),
            .I(N__97002));
    ClkMux I__23754 (
            .O(N__97674),
            .I(N__97002));
    ClkMux I__23753 (
            .O(N__97673),
            .I(N__97002));
    ClkMux I__23752 (
            .O(N__97672),
            .I(N__97002));
    ClkMux I__23751 (
            .O(N__97671),
            .I(N__97002));
    ClkMux I__23750 (
            .O(N__97670),
            .I(N__97002));
    ClkMux I__23749 (
            .O(N__97669),
            .I(N__97002));
    ClkMux I__23748 (
            .O(N__97668),
            .I(N__97002));
    ClkMux I__23747 (
            .O(N__97667),
            .I(N__97002));
    ClkMux I__23746 (
            .O(N__97666),
            .I(N__97002));
    ClkMux I__23745 (
            .O(N__97665),
            .I(N__97002));
    ClkMux I__23744 (
            .O(N__97664),
            .I(N__97002));
    ClkMux I__23743 (
            .O(N__97663),
            .I(N__97002));
    ClkMux I__23742 (
            .O(N__97662),
            .I(N__97002));
    ClkMux I__23741 (
            .O(N__97661),
            .I(N__97002));
    ClkMux I__23740 (
            .O(N__97660),
            .I(N__97002));
    ClkMux I__23739 (
            .O(N__97659),
            .I(N__97002));
    ClkMux I__23738 (
            .O(N__97658),
            .I(N__97002));
    ClkMux I__23737 (
            .O(N__97657),
            .I(N__97002));
    ClkMux I__23736 (
            .O(N__97656),
            .I(N__97002));
    ClkMux I__23735 (
            .O(N__97655),
            .I(N__97002));
    ClkMux I__23734 (
            .O(N__97654),
            .I(N__97002));
    ClkMux I__23733 (
            .O(N__97653),
            .I(N__97002));
    ClkMux I__23732 (
            .O(N__97652),
            .I(N__97002));
    ClkMux I__23731 (
            .O(N__97651),
            .I(N__97002));
    ClkMux I__23730 (
            .O(N__97650),
            .I(N__97002));
    ClkMux I__23729 (
            .O(N__97649),
            .I(N__97002));
    ClkMux I__23728 (
            .O(N__97648),
            .I(N__97002));
    ClkMux I__23727 (
            .O(N__97647),
            .I(N__97002));
    ClkMux I__23726 (
            .O(N__97646),
            .I(N__97002));
    ClkMux I__23725 (
            .O(N__97645),
            .I(N__97002));
    ClkMux I__23724 (
            .O(N__97644),
            .I(N__97002));
    ClkMux I__23723 (
            .O(N__97643),
            .I(N__97002));
    ClkMux I__23722 (
            .O(N__97642),
            .I(N__97002));
    ClkMux I__23721 (
            .O(N__97641),
            .I(N__97002));
    ClkMux I__23720 (
            .O(N__97640),
            .I(N__97002));
    ClkMux I__23719 (
            .O(N__97639),
            .I(N__97002));
    ClkMux I__23718 (
            .O(N__97638),
            .I(N__97002));
    ClkMux I__23717 (
            .O(N__97637),
            .I(N__97002));
    ClkMux I__23716 (
            .O(N__97636),
            .I(N__97002));
    ClkMux I__23715 (
            .O(N__97635),
            .I(N__97002));
    ClkMux I__23714 (
            .O(N__97634),
            .I(N__97002));
    ClkMux I__23713 (
            .O(N__97633),
            .I(N__97002));
    ClkMux I__23712 (
            .O(N__97632),
            .I(N__97002));
    ClkMux I__23711 (
            .O(N__97631),
            .I(N__97002));
    ClkMux I__23710 (
            .O(N__97630),
            .I(N__97002));
    ClkMux I__23709 (
            .O(N__97629),
            .I(N__97002));
    ClkMux I__23708 (
            .O(N__97628),
            .I(N__97002));
    ClkMux I__23707 (
            .O(N__97627),
            .I(N__97002));
    ClkMux I__23706 (
            .O(N__97626),
            .I(N__97002));
    ClkMux I__23705 (
            .O(N__97625),
            .I(N__97002));
    ClkMux I__23704 (
            .O(N__97624),
            .I(N__97002));
    ClkMux I__23703 (
            .O(N__97623),
            .I(N__97002));
    ClkMux I__23702 (
            .O(N__97622),
            .I(N__97002));
    ClkMux I__23701 (
            .O(N__97621),
            .I(N__97002));
    ClkMux I__23700 (
            .O(N__97620),
            .I(N__97002));
    ClkMux I__23699 (
            .O(N__97619),
            .I(N__97002));
    ClkMux I__23698 (
            .O(N__97618),
            .I(N__97002));
    ClkMux I__23697 (
            .O(N__97617),
            .I(N__97002));
    ClkMux I__23696 (
            .O(N__97616),
            .I(N__97002));
    ClkMux I__23695 (
            .O(N__97615),
            .I(N__97002));
    ClkMux I__23694 (
            .O(N__97614),
            .I(N__97002));
    ClkMux I__23693 (
            .O(N__97613),
            .I(N__97002));
    ClkMux I__23692 (
            .O(N__97612),
            .I(N__97002));
    ClkMux I__23691 (
            .O(N__97611),
            .I(N__97002));
    ClkMux I__23690 (
            .O(N__97610),
            .I(N__97002));
    ClkMux I__23689 (
            .O(N__97609),
            .I(N__97002));
    ClkMux I__23688 (
            .O(N__97608),
            .I(N__97002));
    ClkMux I__23687 (
            .O(N__97607),
            .I(N__97002));
    ClkMux I__23686 (
            .O(N__97606),
            .I(N__97002));
    ClkMux I__23685 (
            .O(N__97605),
            .I(N__97002));
    ClkMux I__23684 (
            .O(N__97604),
            .I(N__97002));
    ClkMux I__23683 (
            .O(N__97603),
            .I(N__97002));
    ClkMux I__23682 (
            .O(N__97602),
            .I(N__97002));
    ClkMux I__23681 (
            .O(N__97601),
            .I(N__97002));
    ClkMux I__23680 (
            .O(N__97600),
            .I(N__97002));
    ClkMux I__23679 (
            .O(N__97599),
            .I(N__97002));
    ClkMux I__23678 (
            .O(N__97598),
            .I(N__97002));
    ClkMux I__23677 (
            .O(N__97597),
            .I(N__97002));
    ClkMux I__23676 (
            .O(N__97596),
            .I(N__97002));
    ClkMux I__23675 (
            .O(N__97595),
            .I(N__97002));
    ClkMux I__23674 (
            .O(N__97594),
            .I(N__97002));
    ClkMux I__23673 (
            .O(N__97593),
            .I(N__97002));
    ClkMux I__23672 (
            .O(N__97592),
            .I(N__97002));
    ClkMux I__23671 (
            .O(N__97591),
            .I(N__97002));
    ClkMux I__23670 (
            .O(N__97590),
            .I(N__97002));
    ClkMux I__23669 (
            .O(N__97589),
            .I(N__97002));
    ClkMux I__23668 (
            .O(N__97588),
            .I(N__97002));
    ClkMux I__23667 (
            .O(N__97587),
            .I(N__97002));
    ClkMux I__23666 (
            .O(N__97586),
            .I(N__97002));
    ClkMux I__23665 (
            .O(N__97585),
            .I(N__97002));
    ClkMux I__23664 (
            .O(N__97584),
            .I(N__97002));
    ClkMux I__23663 (
            .O(N__97583),
            .I(N__97002));
    ClkMux I__23662 (
            .O(N__97582),
            .I(N__97002));
    ClkMux I__23661 (
            .O(N__97581),
            .I(N__97002));
    ClkMux I__23660 (
            .O(N__97580),
            .I(N__97002));
    ClkMux I__23659 (
            .O(N__97579),
            .I(N__97002));
    ClkMux I__23658 (
            .O(N__97578),
            .I(N__97002));
    ClkMux I__23657 (
            .O(N__97577),
            .I(N__97002));
    ClkMux I__23656 (
            .O(N__97576),
            .I(N__97002));
    ClkMux I__23655 (
            .O(N__97575),
            .I(N__97002));
    ClkMux I__23654 (
            .O(N__97574),
            .I(N__97002));
    ClkMux I__23653 (
            .O(N__97573),
            .I(N__97002));
    ClkMux I__23652 (
            .O(N__97572),
            .I(N__97002));
    ClkMux I__23651 (
            .O(N__97571),
            .I(N__97002));
    ClkMux I__23650 (
            .O(N__97570),
            .I(N__97002));
    ClkMux I__23649 (
            .O(N__97569),
            .I(N__97002));
    ClkMux I__23648 (
            .O(N__97568),
            .I(N__97002));
    ClkMux I__23647 (
            .O(N__97567),
            .I(N__97002));
    ClkMux I__23646 (
            .O(N__97566),
            .I(N__97002));
    ClkMux I__23645 (
            .O(N__97565),
            .I(N__97002));
    ClkMux I__23644 (
            .O(N__97564),
            .I(N__97002));
    ClkMux I__23643 (
            .O(N__97563),
            .I(N__97002));
    ClkMux I__23642 (
            .O(N__97562),
            .I(N__97002));
    ClkMux I__23641 (
            .O(N__97561),
            .I(N__97002));
    ClkMux I__23640 (
            .O(N__97560),
            .I(N__97002));
    ClkMux I__23639 (
            .O(N__97559),
            .I(N__97002));
    ClkMux I__23638 (
            .O(N__97558),
            .I(N__97002));
    ClkMux I__23637 (
            .O(N__97557),
            .I(N__97002));
    ClkMux I__23636 (
            .O(N__97556),
            .I(N__97002));
    ClkMux I__23635 (
            .O(N__97555),
            .I(N__97002));
    ClkMux I__23634 (
            .O(N__97554),
            .I(N__97002));
    ClkMux I__23633 (
            .O(N__97553),
            .I(N__97002));
    ClkMux I__23632 (
            .O(N__97552),
            .I(N__97002));
    ClkMux I__23631 (
            .O(N__97551),
            .I(N__97002));
    ClkMux I__23630 (
            .O(N__97550),
            .I(N__97002));
    ClkMux I__23629 (
            .O(N__97549),
            .I(N__97002));
    ClkMux I__23628 (
            .O(N__97548),
            .I(N__97002));
    ClkMux I__23627 (
            .O(N__97547),
            .I(N__97002));
    ClkMux I__23626 (
            .O(N__97546),
            .I(N__97002));
    ClkMux I__23625 (
            .O(N__97545),
            .I(N__97002));
    ClkMux I__23624 (
            .O(N__97544),
            .I(N__97002));
    ClkMux I__23623 (
            .O(N__97543),
            .I(N__97002));
    ClkMux I__23622 (
            .O(N__97542),
            .I(N__97002));
    ClkMux I__23621 (
            .O(N__97541),
            .I(N__97002));
    ClkMux I__23620 (
            .O(N__97540),
            .I(N__97002));
    ClkMux I__23619 (
            .O(N__97539),
            .I(N__97002));
    ClkMux I__23618 (
            .O(N__97538),
            .I(N__97002));
    ClkMux I__23617 (
            .O(N__97537),
            .I(N__97002));
    GlobalMux I__23616 (
            .O(N__97002),
            .I(PIN_9_c));
    CEMux I__23615 (
            .O(N__96999),
            .I(N__96992));
    CEMux I__23614 (
            .O(N__96998),
            .I(N__96989));
    CEMux I__23613 (
            .O(N__96997),
            .I(N__96985));
    CEMux I__23612 (
            .O(N__96996),
            .I(N__96982));
    CEMux I__23611 (
            .O(N__96995),
            .I(N__96979));
    LocalMux I__23610 (
            .O(N__96992),
            .I(N__96976));
    LocalMux I__23609 (
            .O(N__96989),
            .I(N__96973));
    CEMux I__23608 (
            .O(N__96988),
            .I(N__96970));
    LocalMux I__23607 (
            .O(N__96985),
            .I(N__96966));
    LocalMux I__23606 (
            .O(N__96982),
            .I(N__96961));
    LocalMux I__23605 (
            .O(N__96979),
            .I(N__96961));
    Span4Mux_v I__23604 (
            .O(N__96976),
            .I(N__96958));
    Span4Mux_v I__23603 (
            .O(N__96973),
            .I(N__96953));
    LocalMux I__23602 (
            .O(N__96970),
            .I(N__96953));
    CEMux I__23601 (
            .O(N__96969),
            .I(N__96950));
    Span4Mux_v I__23600 (
            .O(N__96966),
            .I(N__96945));
    Span4Mux_v I__23599 (
            .O(N__96961),
            .I(N__96936));
    Span4Mux_h I__23598 (
            .O(N__96958),
            .I(N__96936));
    Span4Mux_h I__23597 (
            .O(N__96953),
            .I(N__96936));
    LocalMux I__23596 (
            .O(N__96950),
            .I(N__96936));
    SRMux I__23595 (
            .O(N__96949),
            .I(N__96933));
    CEMux I__23594 (
            .O(N__96948),
            .I(N__96930));
    Span4Mux_v I__23593 (
            .O(N__96945),
            .I(N__96924));
    Span4Mux_h I__23592 (
            .O(N__96936),
            .I(N__96924));
    LocalMux I__23591 (
            .O(N__96933),
            .I(N__96921));
    LocalMux I__23590 (
            .O(N__96930),
            .I(N__96918));
    CEMux I__23589 (
            .O(N__96929),
            .I(N__96915));
    Span4Mux_h I__23588 (
            .O(N__96924),
            .I(N__96911));
    Span4Mux_h I__23587 (
            .O(N__96921),
            .I(N__96908));
    Span4Mux_h I__23586 (
            .O(N__96918),
            .I(N__96905));
    LocalMux I__23585 (
            .O(N__96915),
            .I(N__96902));
    SRMux I__23584 (
            .O(N__96914),
            .I(N__96899));
    Span4Mux_h I__23583 (
            .O(N__96911),
            .I(N__96894));
    Span4Mux_h I__23582 (
            .O(N__96908),
            .I(N__96894));
    Sp12to4 I__23581 (
            .O(N__96905),
            .I(N__96887));
    Span12Mux_v I__23580 (
            .O(N__96902),
            .I(N__96887));
    LocalMux I__23579 (
            .O(N__96899),
            .I(N__96887));
    Odrv4 I__23578 (
            .O(N__96894),
            .I(\c0.n12483 ));
    Odrv12 I__23577 (
            .O(N__96887),
            .I(\c0.n12483 ));
    InMux I__23576 (
            .O(N__96882),
            .I(N__96878));
    InMux I__23575 (
            .O(N__96881),
            .I(N__96875));
    LocalMux I__23574 (
            .O(N__96878),
            .I(\c0.n31283 ));
    LocalMux I__23573 (
            .O(N__96875),
            .I(\c0.n31283 ));
    InMux I__23572 (
            .O(N__96870),
            .I(N__96867));
    LocalMux I__23571 (
            .O(N__96867),
            .I(\c0.n4_adj_4525 ));
    CascadeMux I__23570 (
            .O(N__96864),
            .I(N__96860));
    InMux I__23569 (
            .O(N__96863),
            .I(N__96857));
    InMux I__23568 (
            .O(N__96860),
            .I(N__96854));
    LocalMux I__23567 (
            .O(N__96857),
            .I(N__96851));
    LocalMux I__23566 (
            .O(N__96854),
            .I(N__96848));
    Span4Mux_v I__23565 (
            .O(N__96851),
            .I(N__96843));
    Span4Mux_h I__23564 (
            .O(N__96848),
            .I(N__96843));
    Span4Mux_h I__23563 (
            .O(N__96843),
            .I(N__96840));
    Odrv4 I__23562 (
            .O(N__96840),
            .I(\c0.n15775 ));
    InMux I__23561 (
            .O(N__96837),
            .I(N__96834));
    LocalMux I__23560 (
            .O(N__96834),
            .I(N__96830));
    InMux I__23559 (
            .O(N__96833),
            .I(N__96827));
    Odrv4 I__23558 (
            .O(N__96830),
            .I(\c0.n17576 ));
    LocalMux I__23557 (
            .O(N__96827),
            .I(\c0.n17576 ));
    CascadeMux I__23556 (
            .O(N__96822),
            .I(\c0.n33644_cascade_ ));
    InMux I__23555 (
            .O(N__96819),
            .I(N__96815));
    InMux I__23554 (
            .O(N__96818),
            .I(N__96812));
    LocalMux I__23553 (
            .O(N__96815),
            .I(N__96806));
    LocalMux I__23552 (
            .O(N__96812),
            .I(N__96803));
    InMux I__23551 (
            .O(N__96811),
            .I(N__96800));
    InMux I__23550 (
            .O(N__96810),
            .I(N__96797));
    InMux I__23549 (
            .O(N__96809),
            .I(N__96794));
    Odrv12 I__23548 (
            .O(N__96806),
            .I(\c0.n32273 ));
    Odrv4 I__23547 (
            .O(N__96803),
            .I(\c0.n32273 ));
    LocalMux I__23546 (
            .O(N__96800),
            .I(\c0.n32273 ));
    LocalMux I__23545 (
            .O(N__96797),
            .I(\c0.n32273 ));
    LocalMux I__23544 (
            .O(N__96794),
            .I(\c0.n32273 ));
    InMux I__23543 (
            .O(N__96783),
            .I(N__96780));
    LocalMux I__23542 (
            .O(N__96780),
            .I(N__96777));
    Span4Mux_h I__23541 (
            .O(N__96777),
            .I(N__96773));
    InMux I__23540 (
            .O(N__96776),
            .I(N__96770));
    Odrv4 I__23539 (
            .O(N__96773),
            .I(\c0.n33855 ));
    LocalMux I__23538 (
            .O(N__96770),
            .I(\c0.n33855 ));
    CascadeMux I__23537 (
            .O(N__96765),
            .I(\c0.n31357_cascade_ ));
    InMux I__23536 (
            .O(N__96762),
            .I(N__96759));
    LocalMux I__23535 (
            .O(N__96759),
            .I(N__96755));
    InMux I__23534 (
            .O(N__96758),
            .I(N__96752));
    Span12Mux_v I__23533 (
            .O(N__96755),
            .I(N__96749));
    LocalMux I__23532 (
            .O(N__96752),
            .I(N__96746));
    Odrv12 I__23531 (
            .O(N__96749),
            .I(\c0.n33529 ));
    Odrv12 I__23530 (
            .O(N__96746),
            .I(\c0.n33529 ));
    InMux I__23529 (
            .O(N__96741),
            .I(N__96738));
    LocalMux I__23528 (
            .O(N__96738),
            .I(\c0.n17 ));
    InMux I__23527 (
            .O(N__96735),
            .I(N__96730));
    InMux I__23526 (
            .O(N__96734),
            .I(N__96726));
    CascadeMux I__23525 (
            .O(N__96733),
            .I(N__96722));
    LocalMux I__23524 (
            .O(N__96730),
            .I(N__96719));
    InMux I__23523 (
            .O(N__96729),
            .I(N__96716));
    LocalMux I__23522 (
            .O(N__96726),
            .I(N__96713));
    InMux I__23521 (
            .O(N__96725),
            .I(N__96708));
    InMux I__23520 (
            .O(N__96722),
            .I(N__96708));
    Odrv4 I__23519 (
            .O(N__96719),
            .I(\c0.n32383 ));
    LocalMux I__23518 (
            .O(N__96716),
            .I(\c0.n32383 ));
    Odrv4 I__23517 (
            .O(N__96713),
            .I(\c0.n32383 ));
    LocalMux I__23516 (
            .O(N__96708),
            .I(\c0.n32383 ));
    CascadeMux I__23515 (
            .O(N__96699),
            .I(N__96695));
    InMux I__23514 (
            .O(N__96698),
            .I(N__96692));
    InMux I__23513 (
            .O(N__96695),
            .I(N__96689));
    LocalMux I__23512 (
            .O(N__96692),
            .I(N__96683));
    LocalMux I__23511 (
            .O(N__96689),
            .I(N__96683));
    InMux I__23510 (
            .O(N__96688),
            .I(N__96680));
    Odrv12 I__23509 (
            .O(N__96683),
            .I(\c0.n33644 ));
    LocalMux I__23508 (
            .O(N__96680),
            .I(\c0.n33644 ));
    CascadeMux I__23507 (
            .O(N__96675),
            .I(N__96671));
    CascadeMux I__23506 (
            .O(N__96674),
            .I(N__96668));
    InMux I__23505 (
            .O(N__96671),
            .I(N__96663));
    InMux I__23504 (
            .O(N__96668),
            .I(N__96663));
    LocalMux I__23503 (
            .O(N__96663),
            .I(N__96660));
    Odrv12 I__23502 (
            .O(N__96660),
            .I(\c0.n10_adj_4520 ));
    InMux I__23501 (
            .O(N__96657),
            .I(N__96654));
    LocalMux I__23500 (
            .O(N__96654),
            .I(N__96651));
    Span4Mux_h I__23499 (
            .O(N__96651),
            .I(N__96648));
    Span4Mux_h I__23498 (
            .O(N__96648),
            .I(N__96645));
    Odrv4 I__23497 (
            .O(N__96645),
            .I(\c0.n14_adj_4562 ));
    CascadeMux I__23496 (
            .O(N__96642),
            .I(N__96639));
    InMux I__23495 (
            .O(N__96639),
            .I(N__96635));
    CascadeMux I__23494 (
            .O(N__96638),
            .I(N__96631));
    LocalMux I__23493 (
            .O(N__96635),
            .I(N__96627));
    InMux I__23492 (
            .O(N__96634),
            .I(N__96623));
    InMux I__23491 (
            .O(N__96631),
            .I(N__96620));
    CascadeMux I__23490 (
            .O(N__96630),
            .I(N__96617));
    Span4Mux_h I__23489 (
            .O(N__96627),
            .I(N__96614));
    InMux I__23488 (
            .O(N__96626),
            .I(N__96611));
    LocalMux I__23487 (
            .O(N__96623),
            .I(N__96608));
    LocalMux I__23486 (
            .O(N__96620),
            .I(N__96605));
    InMux I__23485 (
            .O(N__96617),
            .I(N__96602));
    Span4Mux_v I__23484 (
            .O(N__96614),
            .I(N__96596));
    LocalMux I__23483 (
            .O(N__96611),
            .I(N__96596));
    Span4Mux_h I__23482 (
            .O(N__96608),
            .I(N__96593));
    Span4Mux_v I__23481 (
            .O(N__96605),
            .I(N__96588));
    LocalMux I__23480 (
            .O(N__96602),
            .I(N__96588));
    InMux I__23479 (
            .O(N__96601),
            .I(N__96585));
    Span4Mux_h I__23478 (
            .O(N__96596),
            .I(N__96582));
    Span4Mux_h I__23477 (
            .O(N__96593),
            .I(N__96577));
    Span4Mux_h I__23476 (
            .O(N__96588),
            .I(N__96577));
    LocalMux I__23475 (
            .O(N__96585),
            .I(encoder0_position_5));
    Odrv4 I__23474 (
            .O(N__96582),
            .I(encoder0_position_5));
    Odrv4 I__23473 (
            .O(N__96577),
            .I(encoder0_position_5));
    CascadeMux I__23472 (
            .O(N__96570),
            .I(N__96567));
    InMux I__23471 (
            .O(N__96567),
            .I(N__96564));
    LocalMux I__23470 (
            .O(N__96564),
            .I(N__96561));
    Odrv12 I__23469 (
            .O(N__96561),
            .I(\c0.data_out_frame_29__7__N_738 ));
    InMux I__23468 (
            .O(N__96558),
            .I(N__96555));
    LocalMux I__23467 (
            .O(N__96555),
            .I(N__96552));
    Span4Mux_v I__23466 (
            .O(N__96552),
            .I(N__96549));
    Span4Mux_h I__23465 (
            .O(N__96549),
            .I(N__96546));
    Odrv4 I__23464 (
            .O(N__96546),
            .I(\c0.n15 ));
    InMux I__23463 (
            .O(N__96543),
            .I(N__96540));
    LocalMux I__23462 (
            .O(N__96540),
            .I(N__96537));
    Odrv12 I__23461 (
            .O(N__96537),
            .I(\c0.data_out_frame_29_7 ));
    CascadeMux I__23460 (
            .O(N__96534),
            .I(\c0.n10_adj_4573_cascade_ ));
    CascadeMux I__23459 (
            .O(N__96531),
            .I(N__96527));
    InMux I__23458 (
            .O(N__96530),
            .I(N__96522));
    InMux I__23457 (
            .O(N__96527),
            .I(N__96522));
    LocalMux I__23456 (
            .O(N__96522),
            .I(N__96519));
    Odrv4 I__23455 (
            .O(N__96519),
            .I(\c0.n31236 ));
    CascadeMux I__23454 (
            .O(N__96516),
            .I(N__96513));
    InMux I__23453 (
            .O(N__96513),
            .I(N__96507));
    InMux I__23452 (
            .O(N__96512),
            .I(N__96502));
    InMux I__23451 (
            .O(N__96511),
            .I(N__96502));
    InMux I__23450 (
            .O(N__96510),
            .I(N__96499));
    LocalMux I__23449 (
            .O(N__96507),
            .I(N__96496));
    LocalMux I__23448 (
            .O(N__96502),
            .I(N__96493));
    LocalMux I__23447 (
            .O(N__96499),
            .I(N__96488));
    Span4Mux_v I__23446 (
            .O(N__96496),
            .I(N__96485));
    Span4Mux_v I__23445 (
            .O(N__96493),
            .I(N__96482));
    InMux I__23444 (
            .O(N__96492),
            .I(N__96479));
    InMux I__23443 (
            .O(N__96491),
            .I(N__96476));
    Span4Mux_h I__23442 (
            .O(N__96488),
            .I(N__96473));
    Span4Mux_h I__23441 (
            .O(N__96485),
            .I(N__96466));
    Span4Mux_h I__23440 (
            .O(N__96482),
            .I(N__96466));
    LocalMux I__23439 (
            .O(N__96479),
            .I(N__96466));
    LocalMux I__23438 (
            .O(N__96476),
            .I(\c0.n31511 ));
    Odrv4 I__23437 (
            .O(N__96473),
            .I(\c0.n31511 ));
    Odrv4 I__23436 (
            .O(N__96466),
            .I(\c0.n31511 ));
    InMux I__23435 (
            .O(N__96459),
            .I(N__96455));
    InMux I__23434 (
            .O(N__96458),
            .I(N__96452));
    LocalMux I__23433 (
            .O(N__96455),
            .I(N__96448));
    LocalMux I__23432 (
            .O(N__96452),
            .I(N__96445));
    InMux I__23431 (
            .O(N__96451),
            .I(N__96442));
    Span4Mux_h I__23430 (
            .O(N__96448),
            .I(N__96437));
    Span4Mux_v I__23429 (
            .O(N__96445),
            .I(N__96437));
    LocalMux I__23428 (
            .O(N__96442),
            .I(N__96434));
    Span4Mux_v I__23427 (
            .O(N__96437),
            .I(N__96431));
    Odrv4 I__23426 (
            .O(N__96434),
            .I(\c0.n33509 ));
    Odrv4 I__23425 (
            .O(N__96431),
            .I(\c0.n33509 ));
    InMux I__23424 (
            .O(N__96426),
            .I(N__96423));
    LocalMux I__23423 (
            .O(N__96423),
            .I(\c0.n31372 ));
    InMux I__23422 (
            .O(N__96420),
            .I(N__96411));
    InMux I__23421 (
            .O(N__96419),
            .I(N__96411));
    InMux I__23420 (
            .O(N__96418),
            .I(N__96408));
    InMux I__23419 (
            .O(N__96417),
            .I(N__96405));
    InMux I__23418 (
            .O(N__96416),
            .I(N__96402));
    LocalMux I__23417 (
            .O(N__96411),
            .I(N__96397));
    LocalMux I__23416 (
            .O(N__96408),
            .I(N__96397));
    LocalMux I__23415 (
            .O(N__96405),
            .I(\c0.n31516 ));
    LocalMux I__23414 (
            .O(N__96402),
            .I(\c0.n31516 ));
    Odrv4 I__23413 (
            .O(N__96397),
            .I(\c0.n31516 ));
    CascadeMux I__23412 (
            .O(N__96390),
            .I(\c0.n31372_cascade_ ));
    InMux I__23411 (
            .O(N__96387),
            .I(N__96378));
    InMux I__23410 (
            .O(N__96386),
            .I(N__96378));
    InMux I__23409 (
            .O(N__96385),
            .I(N__96378));
    LocalMux I__23408 (
            .O(N__96378),
            .I(\c0.n33588 ));
    CascadeMux I__23407 (
            .O(N__96375),
            .I(\c0.n32437_cascade_ ));
    InMux I__23406 (
            .O(N__96372),
            .I(N__96368));
    InMux I__23405 (
            .O(N__96371),
            .I(N__96365));
    LocalMux I__23404 (
            .O(N__96368),
            .I(N__96362));
    LocalMux I__23403 (
            .O(N__96365),
            .I(\c0.n31287 ));
    Odrv4 I__23402 (
            .O(N__96362),
            .I(\c0.n31287 ));
    InMux I__23401 (
            .O(N__96357),
            .I(N__96351));
    InMux I__23400 (
            .O(N__96356),
            .I(N__96351));
    LocalMux I__23399 (
            .O(N__96351),
            .I(N__96346));
    InMux I__23398 (
            .O(N__96350),
            .I(N__96343));
    InMux I__23397 (
            .O(N__96349),
            .I(N__96340));
    Odrv4 I__23396 (
            .O(N__96346),
            .I(\c0.n32403 ));
    LocalMux I__23395 (
            .O(N__96343),
            .I(\c0.n32403 ));
    LocalMux I__23394 (
            .O(N__96340),
            .I(\c0.n32403 ));
    InMux I__23393 (
            .O(N__96333),
            .I(N__96329));
    InMux I__23392 (
            .O(N__96332),
            .I(N__96325));
    LocalMux I__23391 (
            .O(N__96329),
            .I(N__96322));
    InMux I__23390 (
            .O(N__96328),
            .I(N__96319));
    LocalMux I__23389 (
            .O(N__96325),
            .I(\c0.n35212 ));
    Odrv4 I__23388 (
            .O(N__96322),
            .I(\c0.n35212 ));
    LocalMux I__23387 (
            .O(N__96319),
            .I(\c0.n35212 ));
    CascadeMux I__23386 (
            .O(N__96312),
            .I(N__96309));
    InMux I__23385 (
            .O(N__96309),
            .I(N__96306));
    LocalMux I__23384 (
            .O(N__96306),
            .I(N__96303));
    Odrv4 I__23383 (
            .O(N__96303),
            .I(\c0.n33656 ));
    InMux I__23382 (
            .O(N__96300),
            .I(N__96293));
    InMux I__23381 (
            .O(N__96299),
            .I(N__96288));
    InMux I__23380 (
            .O(N__96298),
            .I(N__96288));
    InMux I__23379 (
            .O(N__96297),
            .I(N__96285));
    InMux I__23378 (
            .O(N__96296),
            .I(N__96282));
    LocalMux I__23377 (
            .O(N__96293),
            .I(N__96279));
    LocalMux I__23376 (
            .O(N__96288),
            .I(N__96274));
    LocalMux I__23375 (
            .O(N__96285),
            .I(N__96274));
    LocalMux I__23374 (
            .O(N__96282),
            .I(N__96271));
    Span4Mux_h I__23373 (
            .O(N__96279),
            .I(N__96265));
    Span4Mux_v I__23372 (
            .O(N__96274),
            .I(N__96265));
    Span4Mux_h I__23371 (
            .O(N__96271),
            .I(N__96262));
    InMux I__23370 (
            .O(N__96270),
            .I(N__96259));
    Span4Mux_h I__23369 (
            .O(N__96265),
            .I(N__96256));
    Odrv4 I__23368 (
            .O(N__96262),
            .I(\c0.n32372 ));
    LocalMux I__23367 (
            .O(N__96259),
            .I(\c0.n32372 ));
    Odrv4 I__23366 (
            .O(N__96256),
            .I(\c0.n32372 ));
    CascadeMux I__23365 (
            .O(N__96249),
            .I(\c0.n7_adj_4521_cascade_ ));
    InMux I__23364 (
            .O(N__96246),
            .I(N__96243));
    LocalMux I__23363 (
            .O(N__96243),
            .I(N__96236));
    InMux I__23362 (
            .O(N__96242),
            .I(N__96227));
    InMux I__23361 (
            .O(N__96241),
            .I(N__96227));
    InMux I__23360 (
            .O(N__96240),
            .I(N__96227));
    InMux I__23359 (
            .O(N__96239),
            .I(N__96227));
    Odrv4 I__23358 (
            .O(N__96236),
            .I(\c0.data_out_frame_29__4__N_1639 ));
    LocalMux I__23357 (
            .O(N__96227),
            .I(\c0.data_out_frame_29__4__N_1639 ));
    InMux I__23356 (
            .O(N__96222),
            .I(N__96219));
    LocalMux I__23355 (
            .O(N__96219),
            .I(N__96214));
    InMux I__23354 (
            .O(N__96218),
            .I(N__96209));
    InMux I__23353 (
            .O(N__96217),
            .I(N__96209));
    Span4Mux_v I__23352 (
            .O(N__96214),
            .I(N__96204));
    LocalMux I__23351 (
            .O(N__96209),
            .I(N__96204));
    Span4Mux_h I__23350 (
            .O(N__96204),
            .I(N__96201));
    Odrv4 I__23349 (
            .O(N__96201),
            .I(\c0.n15827 ));
    CascadeMux I__23348 (
            .O(N__96198),
            .I(\c0.n32383_cascade_ ));
    InMux I__23347 (
            .O(N__96195),
            .I(N__96192));
    LocalMux I__23346 (
            .O(N__96192),
            .I(\c0.data_out_frame_29_0 ));
    InMux I__23345 (
            .O(N__96189),
            .I(N__96186));
    LocalMux I__23344 (
            .O(N__96186),
            .I(\c0.data_out_frame_28_0 ));
    InMux I__23343 (
            .O(N__96183),
            .I(N__96171));
    InMux I__23342 (
            .O(N__96182),
            .I(N__96164));
    InMux I__23341 (
            .O(N__96181),
            .I(N__96161));
    InMux I__23340 (
            .O(N__96180),
            .I(N__96156));
    InMux I__23339 (
            .O(N__96179),
            .I(N__96152));
    CascadeMux I__23338 (
            .O(N__96178),
            .I(N__96149));
    InMux I__23337 (
            .O(N__96177),
            .I(N__96146));
    CascadeMux I__23336 (
            .O(N__96176),
            .I(N__96142));
    CascadeMux I__23335 (
            .O(N__96175),
            .I(N__96139));
    CascadeMux I__23334 (
            .O(N__96174),
            .I(N__96136));
    LocalMux I__23333 (
            .O(N__96171),
            .I(N__96132));
    InMux I__23332 (
            .O(N__96170),
            .I(N__96127));
    InMux I__23331 (
            .O(N__96169),
            .I(N__96127));
    InMux I__23330 (
            .O(N__96168),
            .I(N__96124));
    CascadeMux I__23329 (
            .O(N__96167),
            .I(N__96115));
    LocalMux I__23328 (
            .O(N__96164),
            .I(N__96104));
    LocalMux I__23327 (
            .O(N__96161),
            .I(N__96101));
    InMux I__23326 (
            .O(N__96160),
            .I(N__96096));
    InMux I__23325 (
            .O(N__96159),
            .I(N__96096));
    LocalMux I__23324 (
            .O(N__96156),
            .I(N__96093));
    InMux I__23323 (
            .O(N__96155),
            .I(N__96090));
    LocalMux I__23322 (
            .O(N__96152),
            .I(N__96087));
    InMux I__23321 (
            .O(N__96149),
            .I(N__96084));
    LocalMux I__23320 (
            .O(N__96146),
            .I(N__96081));
    InMux I__23319 (
            .O(N__96145),
            .I(N__96078));
    InMux I__23318 (
            .O(N__96142),
            .I(N__96075));
    InMux I__23317 (
            .O(N__96139),
            .I(N__96072));
    InMux I__23316 (
            .O(N__96136),
            .I(N__96069));
    InMux I__23315 (
            .O(N__96135),
            .I(N__96064));
    Span4Mux_v I__23314 (
            .O(N__96132),
            .I(N__96059));
    LocalMux I__23313 (
            .O(N__96127),
            .I(N__96059));
    LocalMux I__23312 (
            .O(N__96124),
            .I(N__96056));
    CascadeMux I__23311 (
            .O(N__96123),
            .I(N__96052));
    InMux I__23310 (
            .O(N__96122),
            .I(N__96049));
    InMux I__23309 (
            .O(N__96121),
            .I(N__96044));
    InMux I__23308 (
            .O(N__96120),
            .I(N__96044));
    InMux I__23307 (
            .O(N__96119),
            .I(N__96039));
    InMux I__23306 (
            .O(N__96118),
            .I(N__96039));
    InMux I__23305 (
            .O(N__96115),
            .I(N__96036));
    InMux I__23304 (
            .O(N__96114),
            .I(N__96033));
    InMux I__23303 (
            .O(N__96113),
            .I(N__96030));
    InMux I__23302 (
            .O(N__96112),
            .I(N__96027));
    InMux I__23301 (
            .O(N__96111),
            .I(N__96022));
    InMux I__23300 (
            .O(N__96110),
            .I(N__96022));
    CascadeMux I__23299 (
            .O(N__96109),
            .I(N__96017));
    InMux I__23298 (
            .O(N__96108),
            .I(N__96011));
    InMux I__23297 (
            .O(N__96107),
            .I(N__96008));
    Span4Mux_v I__23296 (
            .O(N__96104),
            .I(N__95999));
    Span4Mux_h I__23295 (
            .O(N__96101),
            .I(N__95999));
    LocalMux I__23294 (
            .O(N__96096),
            .I(N__95999));
    Span4Mux_v I__23293 (
            .O(N__96093),
            .I(N__95999));
    LocalMux I__23292 (
            .O(N__96090),
            .I(N__95990));
    Span4Mux_h I__23291 (
            .O(N__96087),
            .I(N__95990));
    LocalMux I__23290 (
            .O(N__96084),
            .I(N__95990));
    Span4Mux_v I__23289 (
            .O(N__96081),
            .I(N__95990));
    LocalMux I__23288 (
            .O(N__96078),
            .I(N__95986));
    LocalMux I__23287 (
            .O(N__96075),
            .I(N__95979));
    LocalMux I__23286 (
            .O(N__96072),
            .I(N__95979));
    LocalMux I__23285 (
            .O(N__96069),
            .I(N__95979));
    InMux I__23284 (
            .O(N__96068),
            .I(N__95976));
    InMux I__23283 (
            .O(N__96067),
            .I(N__95973));
    LocalMux I__23282 (
            .O(N__96064),
            .I(N__95970));
    Span4Mux_v I__23281 (
            .O(N__96059),
            .I(N__95967));
    Span4Mux_v I__23280 (
            .O(N__96056),
            .I(N__95963));
    InMux I__23279 (
            .O(N__96055),
            .I(N__95958));
    InMux I__23278 (
            .O(N__96052),
            .I(N__95958));
    LocalMux I__23277 (
            .O(N__96049),
            .I(N__95951));
    LocalMux I__23276 (
            .O(N__96044),
            .I(N__95951));
    LocalMux I__23275 (
            .O(N__96039),
            .I(N__95951));
    LocalMux I__23274 (
            .O(N__96036),
            .I(N__95940));
    LocalMux I__23273 (
            .O(N__96033),
            .I(N__95940));
    LocalMux I__23272 (
            .O(N__96030),
            .I(N__95940));
    LocalMux I__23271 (
            .O(N__96027),
            .I(N__95940));
    LocalMux I__23270 (
            .O(N__96022),
            .I(N__95940));
    InMux I__23269 (
            .O(N__96021),
            .I(N__95935));
    InMux I__23268 (
            .O(N__96020),
            .I(N__95935));
    InMux I__23267 (
            .O(N__96017),
            .I(N__95930));
    InMux I__23266 (
            .O(N__96016),
            .I(N__95930));
    InMux I__23265 (
            .O(N__96015),
            .I(N__95927));
    InMux I__23264 (
            .O(N__96014),
            .I(N__95924));
    LocalMux I__23263 (
            .O(N__96011),
            .I(N__95919));
    LocalMux I__23262 (
            .O(N__96008),
            .I(N__95919));
    Span4Mux_h I__23261 (
            .O(N__95999),
            .I(N__95914));
    Span4Mux_v I__23260 (
            .O(N__95990),
            .I(N__95914));
    InMux I__23259 (
            .O(N__95989),
            .I(N__95909));
    Span4Mux_v I__23258 (
            .O(N__95986),
            .I(N__95904));
    Span4Mux_v I__23257 (
            .O(N__95979),
            .I(N__95904));
    LocalMux I__23256 (
            .O(N__95976),
            .I(N__95899));
    LocalMux I__23255 (
            .O(N__95973),
            .I(N__95899));
    Span4Mux_v I__23254 (
            .O(N__95970),
            .I(N__95896));
    Span4Mux_h I__23253 (
            .O(N__95967),
            .I(N__95893));
    InMux I__23252 (
            .O(N__95966),
            .I(N__95890));
    Span4Mux_h I__23251 (
            .O(N__95963),
            .I(N__95883));
    LocalMux I__23250 (
            .O(N__95958),
            .I(N__95883));
    Span4Mux_v I__23249 (
            .O(N__95951),
            .I(N__95883));
    Span4Mux_v I__23248 (
            .O(N__95940),
            .I(N__95880));
    LocalMux I__23247 (
            .O(N__95935),
            .I(N__95867));
    LocalMux I__23246 (
            .O(N__95930),
            .I(N__95867));
    LocalMux I__23245 (
            .O(N__95927),
            .I(N__95867));
    LocalMux I__23244 (
            .O(N__95924),
            .I(N__95867));
    Span4Mux_v I__23243 (
            .O(N__95919),
            .I(N__95867));
    Span4Mux_h I__23242 (
            .O(N__95914),
            .I(N__95867));
    InMux I__23241 (
            .O(N__95913),
            .I(N__95864));
    InMux I__23240 (
            .O(N__95912),
            .I(N__95861));
    LocalMux I__23239 (
            .O(N__95909),
            .I(N__95856));
    Span4Mux_h I__23238 (
            .O(N__95904),
            .I(N__95856));
    Span4Mux_v I__23237 (
            .O(N__95899),
            .I(N__95845));
    Span4Mux_v I__23236 (
            .O(N__95896),
            .I(N__95845));
    Span4Mux_h I__23235 (
            .O(N__95893),
            .I(N__95845));
    LocalMux I__23234 (
            .O(N__95890),
            .I(N__95845));
    Span4Mux_v I__23233 (
            .O(N__95883),
            .I(N__95845));
    Span4Mux_h I__23232 (
            .O(N__95880),
            .I(N__95840));
    Span4Mux_v I__23231 (
            .O(N__95867),
            .I(N__95840));
    LocalMux I__23230 (
            .O(N__95864),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__23229 (
            .O(N__95861),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__23228 (
            .O(N__95856),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__23227 (
            .O(N__95845),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__23226 (
            .O(N__95840),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__23225 (
            .O(N__95829),
            .I(N__95826));
    LocalMux I__23224 (
            .O(N__95826),
            .I(N__95823));
    Span4Mux_v I__23223 (
            .O(N__95823),
            .I(N__95820));
    Span4Mux_h I__23222 (
            .O(N__95820),
            .I(N__95817));
    Odrv4 I__23221 (
            .O(N__95817),
            .I(\c0.n35983 ));
    InMux I__23220 (
            .O(N__95814),
            .I(N__95811));
    LocalMux I__23219 (
            .O(N__95811),
            .I(N__95808));
    Span4Mux_h I__23218 (
            .O(N__95808),
            .I(N__95805));
    Span4Mux_h I__23217 (
            .O(N__95805),
            .I(N__95802));
    Odrv4 I__23216 (
            .O(N__95802),
            .I(\c0.n4 ));
    CascadeMux I__23215 (
            .O(N__95799),
            .I(\c0.n26_cascade_ ));
    InMux I__23214 (
            .O(N__95796),
            .I(N__95792));
    InMux I__23213 (
            .O(N__95795),
            .I(N__95786));
    LocalMux I__23212 (
            .O(N__95792),
            .I(N__95783));
    InMux I__23211 (
            .O(N__95791),
            .I(N__95780));
    InMux I__23210 (
            .O(N__95790),
            .I(N__95777));
    CascadeMux I__23209 (
            .O(N__95789),
            .I(N__95773));
    LocalMux I__23208 (
            .O(N__95786),
            .I(N__95769));
    Span4Mux_h I__23207 (
            .O(N__95783),
            .I(N__95766));
    LocalMux I__23206 (
            .O(N__95780),
            .I(N__95763));
    LocalMux I__23205 (
            .O(N__95777),
            .I(N__95759));
    InMux I__23204 (
            .O(N__95776),
            .I(N__95756));
    InMux I__23203 (
            .O(N__95773),
            .I(N__95753));
    InMux I__23202 (
            .O(N__95772),
            .I(N__95750));
    Span4Mux_v I__23201 (
            .O(N__95769),
            .I(N__95747));
    Span4Mux_h I__23200 (
            .O(N__95766),
            .I(N__95742));
    Span4Mux_v I__23199 (
            .O(N__95763),
            .I(N__95742));
    InMux I__23198 (
            .O(N__95762),
            .I(N__95738));
    Span4Mux_v I__23197 (
            .O(N__95759),
            .I(N__95735));
    LocalMux I__23196 (
            .O(N__95756),
            .I(N__95729));
    LocalMux I__23195 (
            .O(N__95753),
            .I(N__95720));
    LocalMux I__23194 (
            .O(N__95750),
            .I(N__95720));
    Span4Mux_v I__23193 (
            .O(N__95747),
            .I(N__95720));
    Span4Mux_h I__23192 (
            .O(N__95742),
            .I(N__95720));
    InMux I__23191 (
            .O(N__95741),
            .I(N__95717));
    LocalMux I__23190 (
            .O(N__95738),
            .I(N__95714));
    Span4Mux_h I__23189 (
            .O(N__95735),
            .I(N__95711));
    InMux I__23188 (
            .O(N__95734),
            .I(N__95708));
    InMux I__23187 (
            .O(N__95733),
            .I(N__95705));
    InMux I__23186 (
            .O(N__95732),
            .I(N__95702));
    Span12Mux_v I__23185 (
            .O(N__95729),
            .I(N__95699));
    Span4Mux_v I__23184 (
            .O(N__95720),
            .I(N__95694));
    LocalMux I__23183 (
            .O(N__95717),
            .I(N__95694));
    Span4Mux_v I__23182 (
            .O(N__95714),
            .I(N__95689));
    Span4Mux_h I__23181 (
            .O(N__95711),
            .I(N__95689));
    LocalMux I__23180 (
            .O(N__95708),
            .I(byte_transmit_counter_3));
    LocalMux I__23179 (
            .O(N__95705),
            .I(byte_transmit_counter_3));
    LocalMux I__23178 (
            .O(N__95702),
            .I(byte_transmit_counter_3));
    Odrv12 I__23177 (
            .O(N__95699),
            .I(byte_transmit_counter_3));
    Odrv4 I__23176 (
            .O(N__95694),
            .I(byte_transmit_counter_3));
    Odrv4 I__23175 (
            .O(N__95689),
            .I(byte_transmit_counter_3));
    InMux I__23174 (
            .O(N__95676),
            .I(N__95673));
    LocalMux I__23173 (
            .O(N__95673),
            .I(N__95670));
    Odrv12 I__23172 (
            .O(N__95670),
            .I(\c0.n35819 ));
    InMux I__23171 (
            .O(N__95667),
            .I(N__95663));
    InMux I__23170 (
            .O(N__95666),
            .I(N__95660));
    LocalMux I__23169 (
            .O(N__95663),
            .I(N__95657));
    LocalMux I__23168 (
            .O(N__95660),
            .I(\c0.n33557 ));
    Odrv4 I__23167 (
            .O(N__95657),
            .I(\c0.n33557 ));
    CascadeMux I__23166 (
            .O(N__95652),
            .I(N__95649));
    InMux I__23165 (
            .O(N__95649),
            .I(N__95646));
    LocalMux I__23164 (
            .O(N__95646),
            .I(N__95643));
    Span4Mux_v I__23163 (
            .O(N__95643),
            .I(N__95639));
    InMux I__23162 (
            .O(N__95642),
            .I(N__95636));
    Span4Mux_h I__23161 (
            .O(N__95639),
            .I(N__95633));
    LocalMux I__23160 (
            .O(N__95636),
            .I(N__95630));
    Odrv4 I__23159 (
            .O(N__95633),
            .I(data_out_frame_29__6__N_1518));
    Odrv4 I__23158 (
            .O(N__95630),
            .I(data_out_frame_29__6__N_1518));
    InMux I__23157 (
            .O(N__95625),
            .I(\quad_counter1.n30488 ));
    InMux I__23156 (
            .O(N__95622),
            .I(N__95617));
    InMux I__23155 (
            .O(N__95621),
            .I(N__95614));
    InMux I__23154 (
            .O(N__95620),
            .I(N__95611));
    LocalMux I__23153 (
            .O(N__95617),
            .I(N__95608));
    LocalMux I__23152 (
            .O(N__95614),
            .I(\quad_counter1.n2210 ));
    LocalMux I__23151 (
            .O(N__95611),
            .I(\quad_counter1.n2210 ));
    Odrv4 I__23150 (
            .O(N__95608),
            .I(\quad_counter1.n2210 ));
    InMux I__23149 (
            .O(N__95601),
            .I(N__95598));
    LocalMux I__23148 (
            .O(N__95598),
            .I(N__95595));
    Span4Mux_h I__23147 (
            .O(N__95595),
            .I(N__95592));
    Odrv4 I__23146 (
            .O(N__95592),
            .I(\c0.data_out_frame_29_3 ));
    InMux I__23145 (
            .O(N__95589),
            .I(N__95586));
    LocalMux I__23144 (
            .O(N__95586),
            .I(\c0.data_out_frame_29_1 ));
    CascadeMux I__23143 (
            .O(N__95583),
            .I(\c0.data_out_frame_29__2__N_1749_cascade_ ));
    InMux I__23142 (
            .O(N__95580),
            .I(N__95577));
    LocalMux I__23141 (
            .O(N__95577),
            .I(N__95573));
    InMux I__23140 (
            .O(N__95576),
            .I(N__95570));
    Odrv4 I__23139 (
            .O(N__95573),
            .I(\c0.n31338 ));
    LocalMux I__23138 (
            .O(N__95570),
            .I(\c0.n31338 ));
    InMux I__23137 (
            .O(N__95565),
            .I(N__95562));
    LocalMux I__23136 (
            .O(N__95562),
            .I(N__95559));
    Span4Mux_v I__23135 (
            .O(N__95559),
            .I(N__95556));
    Odrv4 I__23134 (
            .O(N__95556),
            .I(\c0.n20 ));
    CascadeMux I__23133 (
            .O(N__95553),
            .I(\c0.n21_cascade_ ));
    InMux I__23132 (
            .O(N__95550),
            .I(N__95547));
    LocalMux I__23131 (
            .O(N__95547),
            .I(\c0.n19 ));
    InMux I__23130 (
            .O(N__95544),
            .I(N__95538));
    InMux I__23129 (
            .O(N__95543),
            .I(N__95538));
    LocalMux I__23128 (
            .O(N__95538),
            .I(\c0.n31403 ));
    InMux I__23127 (
            .O(N__95535),
            .I(N__95532));
    LocalMux I__23126 (
            .O(N__95532),
            .I(\c0.data_out_frame_29_2 ));
    InMux I__23125 (
            .O(N__95529),
            .I(N__95524));
    InMux I__23124 (
            .O(N__95528),
            .I(N__95521));
    InMux I__23123 (
            .O(N__95527),
            .I(N__95518));
    LocalMux I__23122 (
            .O(N__95524),
            .I(\quad_counter1.n2219 ));
    LocalMux I__23121 (
            .O(N__95521),
            .I(\quad_counter1.n2219 ));
    LocalMux I__23120 (
            .O(N__95518),
            .I(\quad_counter1.n2219 ));
    InMux I__23119 (
            .O(N__95511),
            .I(bfn_27_11_0_));
    InMux I__23118 (
            .O(N__95508),
            .I(N__95503));
    InMux I__23117 (
            .O(N__95507),
            .I(N__95500));
    InMux I__23116 (
            .O(N__95506),
            .I(N__95497));
    LocalMux I__23115 (
            .O(N__95503),
            .I(\quad_counter1.n2218 ));
    LocalMux I__23114 (
            .O(N__95500),
            .I(\quad_counter1.n2218 ));
    LocalMux I__23113 (
            .O(N__95497),
            .I(\quad_counter1.n2218 ));
    InMux I__23112 (
            .O(N__95490),
            .I(\quad_counter1.n30480 ));
    InMux I__23111 (
            .O(N__95487),
            .I(N__95483));
    InMux I__23110 (
            .O(N__95486),
            .I(N__95480));
    LocalMux I__23109 (
            .O(N__95483),
            .I(\quad_counter1.n2118 ));
    LocalMux I__23108 (
            .O(N__95480),
            .I(\quad_counter1.n2118 ));
    InMux I__23107 (
            .O(N__95475),
            .I(N__95470));
    InMux I__23106 (
            .O(N__95474),
            .I(N__95467));
    InMux I__23105 (
            .O(N__95473),
            .I(N__95464));
    LocalMux I__23104 (
            .O(N__95470),
            .I(\quad_counter1.n2217 ));
    LocalMux I__23103 (
            .O(N__95467),
            .I(\quad_counter1.n2217 ));
    LocalMux I__23102 (
            .O(N__95464),
            .I(\quad_counter1.n2217 ));
    InMux I__23101 (
            .O(N__95457),
            .I(\quad_counter1.n30481 ));
    InMux I__23100 (
            .O(N__95454),
            .I(N__95449));
    InMux I__23099 (
            .O(N__95453),
            .I(N__95446));
    InMux I__23098 (
            .O(N__95452),
            .I(N__95443));
    LocalMux I__23097 (
            .O(N__95449),
            .I(\quad_counter1.n2216 ));
    LocalMux I__23096 (
            .O(N__95446),
            .I(\quad_counter1.n2216 ));
    LocalMux I__23095 (
            .O(N__95443),
            .I(\quad_counter1.n2216 ));
    InMux I__23094 (
            .O(N__95436),
            .I(\quad_counter1.n30482 ));
    InMux I__23093 (
            .O(N__95433),
            .I(N__95428));
    InMux I__23092 (
            .O(N__95432),
            .I(N__95425));
    InMux I__23091 (
            .O(N__95431),
            .I(N__95422));
    LocalMux I__23090 (
            .O(N__95428),
            .I(\quad_counter1.n2215 ));
    LocalMux I__23089 (
            .O(N__95425),
            .I(\quad_counter1.n2215 ));
    LocalMux I__23088 (
            .O(N__95422),
            .I(\quad_counter1.n2215 ));
    InMux I__23087 (
            .O(N__95415),
            .I(\quad_counter1.n30483 ));
    InMux I__23086 (
            .O(N__95412),
            .I(N__95407));
    InMux I__23085 (
            .O(N__95411),
            .I(N__95404));
    InMux I__23084 (
            .O(N__95410),
            .I(N__95401));
    LocalMux I__23083 (
            .O(N__95407),
            .I(\quad_counter1.n2214 ));
    LocalMux I__23082 (
            .O(N__95404),
            .I(\quad_counter1.n2214 ));
    LocalMux I__23081 (
            .O(N__95401),
            .I(\quad_counter1.n2214 ));
    InMux I__23080 (
            .O(N__95394),
            .I(\quad_counter1.n30484 ));
    InMux I__23079 (
            .O(N__95391),
            .I(N__95386));
    InMux I__23078 (
            .O(N__95390),
            .I(N__95383));
    InMux I__23077 (
            .O(N__95389),
            .I(N__95380));
    LocalMux I__23076 (
            .O(N__95386),
            .I(\quad_counter1.n2213 ));
    LocalMux I__23075 (
            .O(N__95383),
            .I(\quad_counter1.n2213 ));
    LocalMux I__23074 (
            .O(N__95380),
            .I(\quad_counter1.n2213 ));
    InMux I__23073 (
            .O(N__95373),
            .I(\quad_counter1.n30485 ));
    InMux I__23072 (
            .O(N__95370),
            .I(N__95367));
    LocalMux I__23071 (
            .O(N__95367),
            .I(N__95362));
    InMux I__23070 (
            .O(N__95366),
            .I(N__95359));
    InMux I__23069 (
            .O(N__95365),
            .I(N__95356));
    Odrv4 I__23068 (
            .O(N__95362),
            .I(\quad_counter1.n2212 ));
    LocalMux I__23067 (
            .O(N__95359),
            .I(\quad_counter1.n2212 ));
    LocalMux I__23066 (
            .O(N__95356),
            .I(\quad_counter1.n2212 ));
    InMux I__23065 (
            .O(N__95349),
            .I(\quad_counter1.n30486 ));
    InMux I__23064 (
            .O(N__95346),
            .I(N__95341));
    InMux I__23063 (
            .O(N__95345),
            .I(N__95338));
    InMux I__23062 (
            .O(N__95344),
            .I(N__95335));
    LocalMux I__23061 (
            .O(N__95341),
            .I(N__95332));
    LocalMux I__23060 (
            .O(N__95338),
            .I(\quad_counter1.n2211 ));
    LocalMux I__23059 (
            .O(N__95335),
            .I(\quad_counter1.n2211 ));
    Odrv4 I__23058 (
            .O(N__95332),
            .I(\quad_counter1.n2211 ));
    InMux I__23057 (
            .O(N__95325),
            .I(bfn_27_12_0_));
    InMux I__23056 (
            .O(N__95322),
            .I(N__95317));
    InMux I__23055 (
            .O(N__95321),
            .I(N__95314));
    InMux I__23054 (
            .O(N__95320),
            .I(N__95311));
    LocalMux I__23053 (
            .O(N__95317),
            .I(N__95308));
    LocalMux I__23052 (
            .O(N__95314),
            .I(N__95304));
    LocalMux I__23051 (
            .O(N__95311),
            .I(N__95299));
    Span4Mux_v I__23050 (
            .O(N__95308),
            .I(N__95299));
    InMux I__23049 (
            .O(N__95307),
            .I(N__95296));
    Span4Mux_v I__23048 (
            .O(N__95304),
            .I(N__95293));
    Span4Mux_h I__23047 (
            .O(N__95299),
            .I(N__95290));
    LocalMux I__23046 (
            .O(N__95296),
            .I(\quad_counter1.millisecond_counter_24 ));
    Odrv4 I__23045 (
            .O(N__95293),
            .I(\quad_counter1.millisecond_counter_24 ));
    Odrv4 I__23044 (
            .O(N__95290),
            .I(\quad_counter1.millisecond_counter_24 ));
    CascadeMux I__23043 (
            .O(N__95283),
            .I(N__95280));
    InMux I__23042 (
            .O(N__95280),
            .I(N__95277));
    LocalMux I__23041 (
            .O(N__95277),
            .I(\quad_counter1.n1987 ));
    CascadeMux I__23040 (
            .O(N__95274),
            .I(\quad_counter1.n2019_cascade_ ));
    CascadeMux I__23039 (
            .O(N__95271),
            .I(\quad_counter1.n28283_cascade_ ));
    InMux I__23038 (
            .O(N__95268),
            .I(N__95265));
    LocalMux I__23037 (
            .O(N__95265),
            .I(\quad_counter1.n9 ));
    CascadeMux I__23036 (
            .O(N__95262),
            .I(\quad_counter1.n10_adj_4432_cascade_ ));
    CascadeMux I__23035 (
            .O(N__95259),
            .I(\quad_counter1.n2045_cascade_ ));
    CascadeMux I__23034 (
            .O(N__95256),
            .I(\quad_counter1.n2118_cascade_ ));
    InMux I__23033 (
            .O(N__95253),
            .I(N__95250));
    LocalMux I__23032 (
            .O(N__95250),
            .I(\quad_counter1.n1986 ));
    InMux I__23031 (
            .O(N__95247),
            .I(N__95243));
    CascadeMux I__23030 (
            .O(N__95246),
            .I(N__95240));
    LocalMux I__23029 (
            .O(N__95243),
            .I(N__95236));
    InMux I__23028 (
            .O(N__95240),
            .I(N__95233));
    InMux I__23027 (
            .O(N__95239),
            .I(N__95230));
    Odrv4 I__23026 (
            .O(N__95236),
            .I(\quad_counter1.n1919 ));
    LocalMux I__23025 (
            .O(N__95233),
            .I(\quad_counter1.n1919 ));
    LocalMux I__23024 (
            .O(N__95230),
            .I(\quad_counter1.n1919 ));
    InMux I__23023 (
            .O(N__95223),
            .I(N__95218));
    InMux I__23022 (
            .O(N__95222),
            .I(N__95215));
    InMux I__23021 (
            .O(N__95221),
            .I(N__95212));
    LocalMux I__23020 (
            .O(N__95218),
            .I(N__95209));
    LocalMux I__23019 (
            .O(N__95215),
            .I(N__95206));
    LocalMux I__23018 (
            .O(N__95212),
            .I(N__95203));
    Span4Mux_v I__23017 (
            .O(N__95209),
            .I(N__95199));
    Span4Mux_v I__23016 (
            .O(N__95206),
            .I(N__95196));
    Span4Mux_h I__23015 (
            .O(N__95203),
            .I(N__95193));
    InMux I__23014 (
            .O(N__95202),
            .I(N__95190));
    Span4Mux_h I__23013 (
            .O(N__95199),
            .I(N__95185));
    Span4Mux_h I__23012 (
            .O(N__95196),
            .I(N__95185));
    Span4Mux_h I__23011 (
            .O(N__95193),
            .I(N__95182));
    LocalMux I__23010 (
            .O(N__95190),
            .I(\quad_counter1.millisecond_counter_22 ));
    Odrv4 I__23009 (
            .O(N__95185),
            .I(\quad_counter1.millisecond_counter_22 ));
    Odrv4 I__23008 (
            .O(N__95182),
            .I(\quad_counter1.millisecond_counter_22 ));
    InMux I__23007 (
            .O(N__95175),
            .I(N__95171));
    InMux I__23006 (
            .O(N__95174),
            .I(N__95168));
    LocalMux I__23005 (
            .O(N__95171),
            .I(\quad_counter1.n1913 ));
    LocalMux I__23004 (
            .O(N__95168),
            .I(\quad_counter1.n1913 ));
    CascadeMux I__23003 (
            .O(N__95163),
            .I(\quad_counter1.n1946_cascade_ ));
    InMux I__23002 (
            .O(N__95160),
            .I(N__95157));
    LocalMux I__23001 (
            .O(N__95157),
            .I(\quad_counter1.n1985 ));
    CascadeMux I__23000 (
            .O(N__95154),
            .I(N__95151));
    InMux I__22999 (
            .O(N__95151),
            .I(N__95148));
    LocalMux I__22998 (
            .O(N__95148),
            .I(\quad_counter1.n1984 ));
    CascadeMux I__22997 (
            .O(N__95145),
            .I(\quad_counter1.n2016_cascade_ ));
    InMux I__22996 (
            .O(N__95142),
            .I(N__95137));
    InMux I__22995 (
            .O(N__95141),
            .I(N__95132));
    InMux I__22994 (
            .O(N__95140),
            .I(N__95132));
    LocalMux I__22993 (
            .O(N__95137),
            .I(\quad_counter1.n1917 ));
    LocalMux I__22992 (
            .O(N__95132),
            .I(\quad_counter1.n1917 ));
    CascadeMux I__22991 (
            .O(N__95127),
            .I(\quad_counter1.n28285_cascade_ ));
    InMux I__22990 (
            .O(N__95124),
            .I(N__95119));
    InMux I__22989 (
            .O(N__95123),
            .I(N__95114));
    InMux I__22988 (
            .O(N__95122),
            .I(N__95114));
    LocalMux I__22987 (
            .O(N__95119),
            .I(\quad_counter1.n1918 ));
    LocalMux I__22986 (
            .O(N__95114),
            .I(\quad_counter1.n1918 ));
    InMux I__22985 (
            .O(N__95109),
            .I(N__95106));
    LocalMux I__22984 (
            .O(N__95106),
            .I(\quad_counter1.n10_adj_4431 ));
    CascadeMux I__22983 (
            .O(N__95103),
            .I(N__95100));
    InMux I__22982 (
            .O(N__95100),
            .I(N__95097));
    LocalMux I__22981 (
            .O(N__95097),
            .I(\quad_counter1.n1983 ));
    CascadeMux I__22980 (
            .O(N__95094),
            .I(N__95091));
    InMux I__22979 (
            .O(N__95091),
            .I(N__95086));
    InMux I__22978 (
            .O(N__95090),
            .I(N__95081));
    InMux I__22977 (
            .O(N__95089),
            .I(N__95081));
    LocalMux I__22976 (
            .O(N__95086),
            .I(\quad_counter1.n1916 ));
    LocalMux I__22975 (
            .O(N__95081),
            .I(\quad_counter1.n1916 ));
    InMux I__22974 (
            .O(N__95076),
            .I(N__95073));
    LocalMux I__22973 (
            .O(N__95073),
            .I(\quad_counter1.n1982 ));
    CascadeMux I__22972 (
            .O(N__95070),
            .I(N__95066));
    InMux I__22971 (
            .O(N__95069),
            .I(N__95060));
    InMux I__22970 (
            .O(N__95066),
            .I(N__95060));
    InMux I__22969 (
            .O(N__95065),
            .I(N__95057));
    LocalMux I__22968 (
            .O(N__95060),
            .I(\quad_counter1.n1915 ));
    LocalMux I__22967 (
            .O(N__95057),
            .I(\quad_counter1.n1915 ));
    InMux I__22966 (
            .O(N__95052),
            .I(N__95046));
    InMux I__22965 (
            .O(N__95051),
            .I(N__95046));
    LocalMux I__22964 (
            .O(N__95046),
            .I(N__95043));
    Span4Mux_h I__22963 (
            .O(N__95043),
            .I(N__95040));
    Odrv4 I__22962 (
            .O(N__95040),
            .I(\c0.n32359 ));
    CascadeMux I__22961 (
            .O(N__95037),
            .I(N__95034));
    InMux I__22960 (
            .O(N__95034),
            .I(N__95030));
    InMux I__22959 (
            .O(N__95033),
            .I(N__95027));
    LocalMux I__22958 (
            .O(N__95030),
            .I(N__95022));
    LocalMux I__22957 (
            .O(N__95027),
            .I(N__95022));
    Span4Mux_h I__22956 (
            .O(N__95022),
            .I(N__95019));
    Span4Mux_h I__22955 (
            .O(N__95019),
            .I(N__95016));
    Odrv4 I__22954 (
            .O(N__95016),
            .I(\c0.n31466 ));
    CascadeMux I__22953 (
            .O(N__95013),
            .I(\c0.n32361_cascade_ ));
    CascadeMux I__22952 (
            .O(N__95010),
            .I(N__95004));
    InMux I__22951 (
            .O(N__95009),
            .I(N__94999));
    InMux I__22950 (
            .O(N__95008),
            .I(N__94999));
    InMux I__22949 (
            .O(N__95007),
            .I(N__94996));
    InMux I__22948 (
            .O(N__95004),
            .I(N__94993));
    LocalMux I__22947 (
            .O(N__94999),
            .I(N__94990));
    LocalMux I__22946 (
            .O(N__94996),
            .I(N__94987));
    LocalMux I__22945 (
            .O(N__94993),
            .I(N__94984));
    Span4Mux_v I__22944 (
            .O(N__94990),
            .I(N__94979));
    Span4Mux_v I__22943 (
            .O(N__94987),
            .I(N__94974));
    Span4Mux_h I__22942 (
            .O(N__94984),
            .I(N__94974));
    InMux I__22941 (
            .O(N__94983),
            .I(N__94969));
    InMux I__22940 (
            .O(N__94982),
            .I(N__94969));
    Odrv4 I__22939 (
            .O(N__94979),
            .I(\c0.n32333 ));
    Odrv4 I__22938 (
            .O(N__94974),
            .I(\c0.n32333 ));
    LocalMux I__22937 (
            .O(N__94969),
            .I(\c0.n32333 ));
    CascadeMux I__22936 (
            .O(N__94962),
            .I(N__94959));
    InMux I__22935 (
            .O(N__94959),
            .I(N__94956));
    LocalMux I__22934 (
            .O(N__94956),
            .I(N__94952));
    InMux I__22933 (
            .O(N__94955),
            .I(N__94949));
    Span4Mux_h I__22932 (
            .O(N__94952),
            .I(N__94946));
    LocalMux I__22931 (
            .O(N__94949),
            .I(\c0.n33861 ));
    Odrv4 I__22930 (
            .O(N__94946),
            .I(\c0.n33861 ));
    InMux I__22929 (
            .O(N__94941),
            .I(N__94938));
    LocalMux I__22928 (
            .O(N__94938),
            .I(N__94935));
    Odrv12 I__22927 (
            .O(N__94935),
            .I(\c0.n21_adj_4551 ));
    CascadeMux I__22926 (
            .O(N__94932),
            .I(\c0.n20_adj_4549_cascade_ ));
    CascadeMux I__22925 (
            .O(N__94929),
            .I(N__94925));
    InMux I__22924 (
            .O(N__94928),
            .I(N__94921));
    InMux I__22923 (
            .O(N__94925),
            .I(N__94918));
    InMux I__22922 (
            .O(N__94924),
            .I(N__94915));
    LocalMux I__22921 (
            .O(N__94921),
            .I(N__94910));
    LocalMux I__22920 (
            .O(N__94918),
            .I(N__94910));
    LocalMux I__22919 (
            .O(N__94915),
            .I(N__94904));
    Span4Mux_h I__22918 (
            .O(N__94910),
            .I(N__94904));
    InMux I__22917 (
            .O(N__94909),
            .I(N__94901));
    Span4Mux_v I__22916 (
            .O(N__94904),
            .I(N__94898));
    LocalMux I__22915 (
            .O(N__94901),
            .I(\c0.n32410 ));
    Odrv4 I__22914 (
            .O(N__94898),
            .I(\c0.n32410 ));
    InMux I__22913 (
            .O(N__94893),
            .I(N__94890));
    LocalMux I__22912 (
            .O(N__94890),
            .I(N__94886));
    InMux I__22911 (
            .O(N__94889),
            .I(N__94883));
    Span4Mux_v I__22910 (
            .O(N__94886),
            .I(N__94877));
    LocalMux I__22909 (
            .O(N__94883),
            .I(N__94877));
    InMux I__22908 (
            .O(N__94882),
            .I(N__94874));
    Span4Mux_h I__22907 (
            .O(N__94877),
            .I(N__94871));
    LocalMux I__22906 (
            .O(N__94874),
            .I(\c0.n32424 ));
    Odrv4 I__22905 (
            .O(N__94871),
            .I(\c0.n32424 ));
    CascadeMux I__22904 (
            .O(N__94866),
            .I(\c0.n34466_cascade_ ));
    InMux I__22903 (
            .O(N__94863),
            .I(N__94859));
    InMux I__22902 (
            .O(N__94862),
            .I(N__94856));
    LocalMux I__22901 (
            .O(N__94859),
            .I(N__94852));
    LocalMux I__22900 (
            .O(N__94856),
            .I(N__94849));
    InMux I__22899 (
            .O(N__94855),
            .I(N__94846));
    Span4Mux_h I__22898 (
            .O(N__94852),
            .I(N__94843));
    Odrv4 I__22897 (
            .O(N__94849),
            .I(\c0.FRAME_MATCHER_i_21 ));
    LocalMux I__22896 (
            .O(N__94846),
            .I(\c0.FRAME_MATCHER_i_21 ));
    Odrv4 I__22895 (
            .O(N__94843),
            .I(\c0.FRAME_MATCHER_i_21 ));
    InMux I__22894 (
            .O(N__94836),
            .I(N__94826));
    InMux I__22893 (
            .O(N__94835),
            .I(N__94826));
    InMux I__22892 (
            .O(N__94834),
            .I(N__94822));
    InMux I__22891 (
            .O(N__94833),
            .I(N__94818));
    InMux I__22890 (
            .O(N__94832),
            .I(N__94811));
    InMux I__22889 (
            .O(N__94831),
            .I(N__94808));
    LocalMux I__22888 (
            .O(N__94826),
            .I(N__94805));
    InMux I__22887 (
            .O(N__94825),
            .I(N__94797));
    LocalMux I__22886 (
            .O(N__94822),
            .I(N__94793));
    InMux I__22885 (
            .O(N__94821),
            .I(N__94790));
    LocalMux I__22884 (
            .O(N__94818),
            .I(N__94787));
    InMux I__22883 (
            .O(N__94817),
            .I(N__94775));
    InMux I__22882 (
            .O(N__94816),
            .I(N__94775));
    InMux I__22881 (
            .O(N__94815),
            .I(N__94770));
    InMux I__22880 (
            .O(N__94814),
            .I(N__94770));
    LocalMux I__22879 (
            .O(N__94811),
            .I(N__94763));
    LocalMux I__22878 (
            .O(N__94808),
            .I(N__94763));
    Span4Mux_v I__22877 (
            .O(N__94805),
            .I(N__94763));
    InMux I__22876 (
            .O(N__94804),
            .I(N__94754));
    InMux I__22875 (
            .O(N__94803),
            .I(N__94754));
    InMux I__22874 (
            .O(N__94802),
            .I(N__94754));
    InMux I__22873 (
            .O(N__94801),
            .I(N__94754));
    InMux I__22872 (
            .O(N__94800),
            .I(N__94751));
    LocalMux I__22871 (
            .O(N__94797),
            .I(N__94744));
    InMux I__22870 (
            .O(N__94796),
            .I(N__94741));
    Span4Mux_v I__22869 (
            .O(N__94793),
            .I(N__94738));
    LocalMux I__22868 (
            .O(N__94790),
            .I(N__94735));
    Span4Mux_v I__22867 (
            .O(N__94787),
            .I(N__94732));
    InMux I__22866 (
            .O(N__94786),
            .I(N__94727));
    InMux I__22865 (
            .O(N__94785),
            .I(N__94727));
    InMux I__22864 (
            .O(N__94784),
            .I(N__94724));
    InMux I__22863 (
            .O(N__94783),
            .I(N__94715));
    InMux I__22862 (
            .O(N__94782),
            .I(N__94715));
    InMux I__22861 (
            .O(N__94781),
            .I(N__94715));
    InMux I__22860 (
            .O(N__94780),
            .I(N__94715));
    LocalMux I__22859 (
            .O(N__94775),
            .I(N__94706));
    LocalMux I__22858 (
            .O(N__94770),
            .I(N__94706));
    Span4Mux_v I__22857 (
            .O(N__94763),
            .I(N__94706));
    LocalMux I__22856 (
            .O(N__94754),
            .I(N__94706));
    LocalMux I__22855 (
            .O(N__94751),
            .I(N__94703));
    InMux I__22854 (
            .O(N__94750),
            .I(N__94700));
    InMux I__22853 (
            .O(N__94749),
            .I(N__94694));
    InMux I__22852 (
            .O(N__94748),
            .I(N__94694));
    InMux I__22851 (
            .O(N__94747),
            .I(N__94691));
    Span4Mux_v I__22850 (
            .O(N__94744),
            .I(N__94684));
    LocalMux I__22849 (
            .O(N__94741),
            .I(N__94684));
    Span4Mux_v I__22848 (
            .O(N__94738),
            .I(N__94681));
    Span4Mux_v I__22847 (
            .O(N__94735),
            .I(N__94678));
    Span4Mux_v I__22846 (
            .O(N__94732),
            .I(N__94675));
    LocalMux I__22845 (
            .O(N__94727),
            .I(N__94666));
    LocalMux I__22844 (
            .O(N__94724),
            .I(N__94666));
    LocalMux I__22843 (
            .O(N__94715),
            .I(N__94666));
    Span4Mux_v I__22842 (
            .O(N__94706),
            .I(N__94666));
    Span4Mux_h I__22841 (
            .O(N__94703),
            .I(N__94663));
    LocalMux I__22840 (
            .O(N__94700),
            .I(N__94660));
    InMux I__22839 (
            .O(N__94699),
            .I(N__94657));
    LocalMux I__22838 (
            .O(N__94694),
            .I(N__94654));
    LocalMux I__22837 (
            .O(N__94691),
            .I(N__94651));
    InMux I__22836 (
            .O(N__94690),
            .I(N__94648));
    InMux I__22835 (
            .O(N__94689),
            .I(N__94645));
    Span4Mux_v I__22834 (
            .O(N__94684),
            .I(N__94640));
    Span4Mux_v I__22833 (
            .O(N__94681),
            .I(N__94640));
    Span4Mux_v I__22832 (
            .O(N__94678),
            .I(N__94633));
    Span4Mux_v I__22831 (
            .O(N__94675),
            .I(N__94633));
    Span4Mux_v I__22830 (
            .O(N__94666),
            .I(N__94633));
    Span4Mux_v I__22829 (
            .O(N__94663),
            .I(N__94630));
    Span4Mux_v I__22828 (
            .O(N__94660),
            .I(N__94627));
    LocalMux I__22827 (
            .O(N__94657),
            .I(N__94624));
    Span12Mux_h I__22826 (
            .O(N__94654),
            .I(N__94621));
    Span12Mux_h I__22825 (
            .O(N__94651),
            .I(N__94618));
    LocalMux I__22824 (
            .O(N__94648),
            .I(N__94609));
    LocalMux I__22823 (
            .O(N__94645),
            .I(N__94609));
    Sp12to4 I__22822 (
            .O(N__94640),
            .I(N__94609));
    Sp12to4 I__22821 (
            .O(N__94633),
            .I(N__94609));
    Span4Mux_v I__22820 (
            .O(N__94630),
            .I(N__94604));
    Span4Mux_h I__22819 (
            .O(N__94627),
            .I(N__94604));
    Span4Mux_h I__22818 (
            .O(N__94624),
            .I(N__94601));
    Span12Mux_v I__22817 (
            .O(N__94621),
            .I(N__94592));
    Span12Mux_v I__22816 (
            .O(N__94618),
            .I(N__94592));
    Span12Mux_h I__22815 (
            .O(N__94609),
            .I(N__94592));
    Sp12to4 I__22814 (
            .O(N__94604),
            .I(N__94592));
    Odrv4 I__22813 (
            .O(N__94601),
            .I(\c0.n2107 ));
    Odrv12 I__22812 (
            .O(N__94592),
            .I(\c0.n2107 ));
    SRMux I__22811 (
            .O(N__94587),
            .I(N__94584));
    LocalMux I__22810 (
            .O(N__94584),
            .I(N__94581));
    Odrv4 I__22809 (
            .O(N__94581),
            .I(\c0.n3_adj_4600 ));
    CascadeMux I__22808 (
            .O(N__94578),
            .I(N__94569));
    InMux I__22807 (
            .O(N__94577),
            .I(N__94564));
    InMux I__22806 (
            .O(N__94576),
            .I(N__94564));
    InMux I__22805 (
            .O(N__94575),
            .I(N__94561));
    InMux I__22804 (
            .O(N__94574),
            .I(N__94556));
    InMux I__22803 (
            .O(N__94573),
            .I(N__94556));
    InMux I__22802 (
            .O(N__94572),
            .I(N__94551));
    InMux I__22801 (
            .O(N__94569),
            .I(N__94551));
    LocalMux I__22800 (
            .O(N__94564),
            .I(N__94542));
    LocalMux I__22799 (
            .O(N__94561),
            .I(N__94542));
    LocalMux I__22798 (
            .O(N__94556),
            .I(N__94542));
    LocalMux I__22797 (
            .O(N__94551),
            .I(N__94542));
    Span4Mux_v I__22796 (
            .O(N__94542),
            .I(N__94539));
    Odrv4 I__22795 (
            .O(N__94539),
            .I(\c0.n18499 ));
    InMux I__22794 (
            .O(N__94536),
            .I(N__94528));
    InMux I__22793 (
            .O(N__94535),
            .I(N__94528));
    CascadeMux I__22792 (
            .O(N__94534),
            .I(N__94524));
    InMux I__22791 (
            .O(N__94533),
            .I(N__94521));
    LocalMux I__22790 (
            .O(N__94528),
            .I(N__94518));
    InMux I__22789 (
            .O(N__94527),
            .I(N__94515));
    InMux I__22788 (
            .O(N__94524),
            .I(N__94510));
    LocalMux I__22787 (
            .O(N__94521),
            .I(N__94507));
    Span4Mux_v I__22786 (
            .O(N__94518),
            .I(N__94504));
    LocalMux I__22785 (
            .O(N__94515),
            .I(N__94501));
    InMux I__22784 (
            .O(N__94514),
            .I(N__94498));
    InMux I__22783 (
            .O(N__94513),
            .I(N__94495));
    LocalMux I__22782 (
            .O(N__94510),
            .I(N__94490));
    Span12Mux_s10_h I__22781 (
            .O(N__94507),
            .I(N__94490));
    Span4Mux_h I__22780 (
            .O(N__94504),
            .I(N__94485));
    Span4Mux_v I__22779 (
            .O(N__94501),
            .I(N__94485));
    LocalMux I__22778 (
            .O(N__94498),
            .I(N__94482));
    LocalMux I__22777 (
            .O(N__94495),
            .I(\c0.n18898 ));
    Odrv12 I__22776 (
            .O(N__94490),
            .I(\c0.n18898 ));
    Odrv4 I__22775 (
            .O(N__94485),
            .I(\c0.n18898 ));
    Odrv12 I__22774 (
            .O(N__94482),
            .I(\c0.n18898 ));
    CascadeMux I__22773 (
            .O(N__94473),
            .I(N__94469));
    InMux I__22772 (
            .O(N__94472),
            .I(N__94464));
    InMux I__22771 (
            .O(N__94469),
            .I(N__94464));
    LocalMux I__22770 (
            .O(N__94464),
            .I(N__94460));
    InMux I__22769 (
            .O(N__94463),
            .I(N__94457));
    Span4Mux_h I__22768 (
            .O(N__94460),
            .I(N__94454));
    LocalMux I__22767 (
            .O(N__94457),
            .I(\c0.FRAME_MATCHER_i_17 ));
    Odrv4 I__22766 (
            .O(N__94454),
            .I(\c0.FRAME_MATCHER_i_17 ));
    SRMux I__22765 (
            .O(N__94449),
            .I(N__94446));
    LocalMux I__22764 (
            .O(N__94446),
            .I(N__94443));
    Span4Mux_h I__22763 (
            .O(N__94443),
            .I(N__94440));
    Odrv4 I__22762 (
            .O(N__94440),
            .I(\c0.n3_adj_4596 ));
    CascadeMux I__22761 (
            .O(N__94437),
            .I(\c0.n17574_cascade_ ));
    InMux I__22760 (
            .O(N__94434),
            .I(N__94431));
    LocalMux I__22759 (
            .O(N__94431),
            .I(N__94428));
    Span4Mux_h I__22758 (
            .O(N__94428),
            .I(N__94425));
    Odrv4 I__22757 (
            .O(N__94425),
            .I(\c0.n35251 ));
    InMux I__22756 (
            .O(N__94422),
            .I(N__94417));
    CascadeMux I__22755 (
            .O(N__94421),
            .I(N__94414));
    InMux I__22754 (
            .O(N__94420),
            .I(N__94411));
    LocalMux I__22753 (
            .O(N__94417),
            .I(N__94408));
    InMux I__22752 (
            .O(N__94414),
            .I(N__94405));
    LocalMux I__22751 (
            .O(N__94411),
            .I(N__94402));
    Span4Mux_v I__22750 (
            .O(N__94408),
            .I(N__94399));
    LocalMux I__22749 (
            .O(N__94405),
            .I(N__94396));
    Odrv4 I__22748 (
            .O(N__94402),
            .I(\c0.n31302 ));
    Odrv4 I__22747 (
            .O(N__94399),
            .I(\c0.n31302 ));
    Odrv4 I__22746 (
            .O(N__94396),
            .I(\c0.n31302 ));
    InMux I__22745 (
            .O(N__94389),
            .I(N__94385));
    InMux I__22744 (
            .O(N__94388),
            .I(N__94382));
    LocalMux I__22743 (
            .O(N__94385),
            .I(N__94379));
    LocalMux I__22742 (
            .O(N__94382),
            .I(N__94374));
    Span4Mux_h I__22741 (
            .O(N__94379),
            .I(N__94374));
    Odrv4 I__22740 (
            .O(N__94374),
            .I(\c0.n32476 ));
    InMux I__22739 (
            .O(N__94371),
            .I(N__94367));
    InMux I__22738 (
            .O(N__94370),
            .I(N__94364));
    LocalMux I__22737 (
            .O(N__94367),
            .I(N__94359));
    LocalMux I__22736 (
            .O(N__94364),
            .I(N__94356));
    InMux I__22735 (
            .O(N__94363),
            .I(N__94351));
    InMux I__22734 (
            .O(N__94362),
            .I(N__94351));
    Span4Mux_h I__22733 (
            .O(N__94359),
            .I(N__94348));
    Odrv12 I__22732 (
            .O(N__94356),
            .I(\c0.n18901 ));
    LocalMux I__22731 (
            .O(N__94351),
            .I(\c0.n18901 ));
    Odrv4 I__22730 (
            .O(N__94348),
            .I(\c0.n18901 ));
    InMux I__22729 (
            .O(N__94341),
            .I(N__94338));
    LocalMux I__22728 (
            .O(N__94338),
            .I(N__94335));
    Span4Mux_h I__22727 (
            .O(N__94335),
            .I(N__94332));
    Odrv4 I__22726 (
            .O(N__94332),
            .I(\c0.n14_adj_4523 ));
    CascadeMux I__22725 (
            .O(N__94329),
            .I(\c0.n31463_cascade_ ));
    InMux I__22724 (
            .O(N__94326),
            .I(N__94318));
    InMux I__22723 (
            .O(N__94325),
            .I(N__94318));
    InMux I__22722 (
            .O(N__94324),
            .I(N__94315));
    CascadeMux I__22721 (
            .O(N__94323),
            .I(N__94312));
    LocalMux I__22720 (
            .O(N__94318),
            .I(N__94307));
    LocalMux I__22719 (
            .O(N__94315),
            .I(N__94304));
    InMux I__22718 (
            .O(N__94312),
            .I(N__94301));
    InMux I__22717 (
            .O(N__94311),
            .I(N__94296));
    InMux I__22716 (
            .O(N__94310),
            .I(N__94296));
    Span4Mux_h I__22715 (
            .O(N__94307),
            .I(N__94292));
    Span4Mux_v I__22714 (
            .O(N__94304),
            .I(N__94287));
    LocalMux I__22713 (
            .O(N__94301),
            .I(N__94287));
    LocalMux I__22712 (
            .O(N__94296),
            .I(N__94284));
    InMux I__22711 (
            .O(N__94295),
            .I(N__94281));
    Span4Mux_h I__22710 (
            .O(N__94292),
            .I(N__94278));
    Span4Mux_h I__22709 (
            .O(N__94287),
            .I(N__94273));
    Span4Mux_h I__22708 (
            .O(N__94284),
            .I(N__94273));
    LocalMux I__22707 (
            .O(N__94281),
            .I(encoder1_position_6));
    Odrv4 I__22706 (
            .O(N__94278),
            .I(encoder1_position_6));
    Odrv4 I__22705 (
            .O(N__94273),
            .I(encoder1_position_6));
    InMux I__22704 (
            .O(N__94266),
            .I(N__94263));
    LocalMux I__22703 (
            .O(N__94263),
            .I(N__94259));
    InMux I__22702 (
            .O(N__94262),
            .I(N__94256));
    Span4Mux_h I__22701 (
            .O(N__94259),
            .I(N__94253));
    LocalMux I__22700 (
            .O(N__94256),
            .I(N__94250));
    Odrv4 I__22699 (
            .O(N__94253),
            .I(\c0.n32361 ));
    Odrv12 I__22698 (
            .O(N__94250),
            .I(\c0.n32361 ));
    CascadeMux I__22697 (
            .O(N__94245),
            .I(\c0.n4_adj_4630_cascade_ ));
    CascadeMux I__22696 (
            .O(N__94242),
            .I(N__94239));
    InMux I__22695 (
            .O(N__94239),
            .I(N__94236));
    LocalMux I__22694 (
            .O(N__94236),
            .I(N__94232));
    InMux I__22693 (
            .O(N__94235),
            .I(N__94229));
    Odrv12 I__22692 (
            .O(N__94232),
            .I(\c0.n4_adj_4630 ));
    LocalMux I__22691 (
            .O(N__94229),
            .I(\c0.n4_adj_4630 ));
    InMux I__22690 (
            .O(N__94224),
            .I(N__94221));
    LocalMux I__22689 (
            .O(N__94221),
            .I(N__94218));
    Odrv4 I__22688 (
            .O(N__94218),
            .I(\c0.data_out_frame_29_5 ));
    InMux I__22687 (
            .O(N__94215),
            .I(N__94212));
    LocalMux I__22686 (
            .O(N__94212),
            .I(N__94209));
    Odrv4 I__22685 (
            .O(N__94209),
            .I(\c0.data_out_frame_28_5 ));
    InMux I__22684 (
            .O(N__94206),
            .I(N__94203));
    LocalMux I__22683 (
            .O(N__94203),
            .I(N__94200));
    Span4Mux_h I__22682 (
            .O(N__94200),
            .I(N__94197));
    Odrv4 I__22681 (
            .O(N__94197),
            .I(\c0.n26_adj_4620 ));
    CascadeMux I__22680 (
            .O(N__94194),
            .I(\c0.n32476_cascade_ ));
    InMux I__22679 (
            .O(N__94191),
            .I(N__94187));
    InMux I__22678 (
            .O(N__94190),
            .I(N__94184));
    LocalMux I__22677 (
            .O(N__94187),
            .I(N__94181));
    LocalMux I__22676 (
            .O(N__94184),
            .I(N__94178));
    Span4Mux_v I__22675 (
            .O(N__94181),
            .I(N__94174));
    Span4Mux_h I__22674 (
            .O(N__94178),
            .I(N__94171));
    InMux I__22673 (
            .O(N__94177),
            .I(N__94168));
    Span4Mux_v I__22672 (
            .O(N__94174),
            .I(N__94165));
    Odrv4 I__22671 (
            .O(N__94171),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__22670 (
            .O(N__94168),
            .I(\c0.FRAME_MATCHER_i_24 ));
    Odrv4 I__22669 (
            .O(N__94165),
            .I(\c0.FRAME_MATCHER_i_24 ));
    InMux I__22668 (
            .O(N__94158),
            .I(N__94155));
    LocalMux I__22667 (
            .O(N__94155),
            .I(N__94152));
    Span4Mux_h I__22666 (
            .O(N__94152),
            .I(N__94148));
    InMux I__22665 (
            .O(N__94151),
            .I(N__94145));
    Span4Mux_v I__22664 (
            .O(N__94148),
            .I(N__94141));
    LocalMux I__22663 (
            .O(N__94145),
            .I(N__94138));
    InMux I__22662 (
            .O(N__94144),
            .I(N__94135));
    Span4Mux_v I__22661 (
            .O(N__94141),
            .I(N__94132));
    Odrv4 I__22660 (
            .O(N__94138),
            .I(\c0.FRAME_MATCHER_i_30 ));
    LocalMux I__22659 (
            .O(N__94135),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__22658 (
            .O(N__94132),
            .I(\c0.FRAME_MATCHER_i_30 ));
    InMux I__22657 (
            .O(N__94125),
            .I(N__94122));
    LocalMux I__22656 (
            .O(N__94122),
            .I(N__94119));
    Span4Mux_h I__22655 (
            .O(N__94119),
            .I(N__94116));
    Odrv4 I__22654 (
            .O(N__94116),
            .I(\c0.n44_adj_4639 ));
    InMux I__22653 (
            .O(N__94113),
            .I(N__94109));
    InMux I__22652 (
            .O(N__94112),
            .I(N__94106));
    LocalMux I__22651 (
            .O(N__94109),
            .I(N__94103));
    LocalMux I__22650 (
            .O(N__94106),
            .I(N__94100));
    Odrv12 I__22649 (
            .O(N__94103),
            .I(\c0.n33572 ));
    Odrv12 I__22648 (
            .O(N__94100),
            .I(\c0.n33572 ));
    InMux I__22647 (
            .O(N__94095),
            .I(N__94091));
    InMux I__22646 (
            .O(N__94094),
            .I(N__94088));
    LocalMux I__22645 (
            .O(N__94091),
            .I(\c0.n32271 ));
    LocalMux I__22644 (
            .O(N__94088),
            .I(\c0.n32271 ));
    CascadeMux I__22643 (
            .O(N__94083),
            .I(\c0.n32300_cascade_ ));
    InMux I__22642 (
            .O(N__94080),
            .I(N__94077));
    LocalMux I__22641 (
            .O(N__94077),
            .I(N__94073));
    InMux I__22640 (
            .O(N__94076),
            .I(N__94070));
    Span4Mux_h I__22639 (
            .O(N__94073),
            .I(N__94067));
    LocalMux I__22638 (
            .O(N__94070),
            .I(N__94064));
    Odrv4 I__22637 (
            .O(N__94067),
            .I(\c0.n31280 ));
    Odrv4 I__22636 (
            .O(N__94064),
            .I(\c0.n31280 ));
    InMux I__22635 (
            .O(N__94059),
            .I(N__94056));
    LocalMux I__22634 (
            .O(N__94056),
            .I(N__94053));
    Span4Mux_h I__22633 (
            .O(N__94053),
            .I(N__94050));
    Span4Mux_v I__22632 (
            .O(N__94050),
            .I(N__94047));
    Odrv4 I__22631 (
            .O(N__94047),
            .I(\c0.n32454 ));
    CascadeMux I__22630 (
            .O(N__94044),
            .I(\c0.n32454_cascade_ ));
    InMux I__22629 (
            .O(N__94041),
            .I(N__94038));
    LocalMux I__22628 (
            .O(N__94038),
            .I(\c0.n32445 ));
    InMux I__22627 (
            .O(N__94035),
            .I(N__94031));
    InMux I__22626 (
            .O(N__94034),
            .I(N__94028));
    LocalMux I__22625 (
            .O(N__94031),
            .I(\c0.n32331 ));
    LocalMux I__22624 (
            .O(N__94028),
            .I(\c0.n32331 ));
    InMux I__22623 (
            .O(N__94023),
            .I(N__94016));
    InMux I__22622 (
            .O(N__94022),
            .I(N__94016));
    CascadeMux I__22621 (
            .O(N__94021),
            .I(N__94012));
    LocalMux I__22620 (
            .O(N__94016),
            .I(N__94009));
    InMux I__22619 (
            .O(N__94015),
            .I(N__94004));
    InMux I__22618 (
            .O(N__94012),
            .I(N__94004));
    Span4Mux_v I__22617 (
            .O(N__94009),
            .I(N__93999));
    LocalMux I__22616 (
            .O(N__94004),
            .I(N__93999));
    Odrv4 I__22615 (
            .O(N__93999),
            .I(\c0.n32377 ));
    InMux I__22614 (
            .O(N__93996),
            .I(N__93993));
    LocalMux I__22613 (
            .O(N__93993),
            .I(N__93989));
    CascadeMux I__22612 (
            .O(N__93992),
            .I(N__93985));
    Span4Mux_h I__22611 (
            .O(N__93989),
            .I(N__93982));
    InMux I__22610 (
            .O(N__93988),
            .I(N__93977));
    InMux I__22609 (
            .O(N__93985),
            .I(N__93977));
    Odrv4 I__22608 (
            .O(N__93982),
            .I(\c0.n32300 ));
    LocalMux I__22607 (
            .O(N__93977),
            .I(\c0.n32300 ));
    CascadeMux I__22606 (
            .O(N__93972),
            .I(\c0.n32331_cascade_ ));
    InMux I__22605 (
            .O(N__93969),
            .I(N__93966));
    LocalMux I__22604 (
            .O(N__93966),
            .I(N__93963));
    Span4Mux_h I__22603 (
            .O(N__93963),
            .I(N__93960));
    Odrv4 I__22602 (
            .O(N__93960),
            .I(n35623));
    InMux I__22601 (
            .O(N__93957),
            .I(N__93953));
    InMux I__22600 (
            .O(N__93956),
            .I(N__93950));
    LocalMux I__22599 (
            .O(N__93953),
            .I(N__93945));
    LocalMux I__22598 (
            .O(N__93950),
            .I(N__93945));
    Span4Mux_v I__22597 (
            .O(N__93945),
            .I(N__93941));
    InMux I__22596 (
            .O(N__93944),
            .I(N__93938));
    Odrv4 I__22595 (
            .O(N__93941),
            .I(\quad_counter1.n2309 ));
    LocalMux I__22594 (
            .O(N__93938),
            .I(\quad_counter1.n2309 ));
    InMux I__22593 (
            .O(N__93933),
            .I(N__93929));
    InMux I__22592 (
            .O(N__93932),
            .I(N__93926));
    LocalMux I__22591 (
            .O(N__93929),
            .I(N__93921));
    LocalMux I__22590 (
            .O(N__93926),
            .I(N__93921));
    Span4Mux_h I__22589 (
            .O(N__93921),
            .I(N__93917));
    InMux I__22588 (
            .O(N__93920),
            .I(N__93914));
    Odrv4 I__22587 (
            .O(N__93917),
            .I(\quad_counter1.n2312 ));
    LocalMux I__22586 (
            .O(N__93914),
            .I(\quad_counter1.n2312 ));
    InMux I__22585 (
            .O(N__93909),
            .I(N__93906));
    LocalMux I__22584 (
            .O(N__93906),
            .I(N__93903));
    Span4Mux_h I__22583 (
            .O(N__93903),
            .I(N__93900));
    Odrv4 I__22582 (
            .O(N__93900),
            .I(\quad_counter1.n8_adj_4438 ));
    CascadeMux I__22581 (
            .O(N__93897),
            .I(\c0.n6_adj_4533_cascade_ ));
    InMux I__22580 (
            .O(N__93894),
            .I(N__93891));
    LocalMux I__22579 (
            .O(N__93891),
            .I(\c0.data_out_frame_28_2 ));
    InMux I__22578 (
            .O(N__93888),
            .I(N__93885));
    LocalMux I__22577 (
            .O(N__93885),
            .I(N__93882));
    Span4Mux_h I__22576 (
            .O(N__93882),
            .I(N__93879));
    Span4Mux_h I__22575 (
            .O(N__93879),
            .I(N__93876));
    Span4Mux_h I__22574 (
            .O(N__93876),
            .I(N__93873));
    Odrv4 I__22573 (
            .O(N__93873),
            .I(\c0.n26_adj_4512 ));
    CascadeMux I__22572 (
            .O(N__93870),
            .I(\c0.n32271_cascade_ ));
    InMux I__22571 (
            .O(N__93867),
            .I(N__93864));
    LocalMux I__22570 (
            .O(N__93864),
            .I(\c0.data_out_frame_28_1 ));
    InMux I__22569 (
            .O(N__93861),
            .I(N__93858));
    LocalMux I__22568 (
            .O(N__93858),
            .I(N__93855));
    Span4Mux_h I__22567 (
            .O(N__93855),
            .I(N__93852));
    Span4Mux_h I__22566 (
            .O(N__93852),
            .I(N__93849));
    Odrv4 I__22565 (
            .O(N__93849),
            .I(\c0.n26_adj_4506 ));
    InMux I__22564 (
            .O(N__93846),
            .I(N__93843));
    LocalMux I__22563 (
            .O(N__93843),
            .I(N__93840));
    Sp12to4 I__22562 (
            .O(N__93840),
            .I(N__93837));
    Span12Mux_v I__22561 (
            .O(N__93837),
            .I(N__93834));
    Odrv12 I__22560 (
            .O(N__93834),
            .I(\c0.data_out_frame_28_4 ));
    InMux I__22559 (
            .O(N__93831),
            .I(N__93827));
    InMux I__22558 (
            .O(N__93830),
            .I(N__93824));
    LocalMux I__22557 (
            .O(N__93827),
            .I(N__93821));
    LocalMux I__22556 (
            .O(N__93824),
            .I(N__93818));
    Span4Mux_h I__22555 (
            .O(N__93821),
            .I(N__93815));
    Odrv4 I__22554 (
            .O(N__93818),
            .I(\c0.n33607 ));
    Odrv4 I__22553 (
            .O(N__93815),
            .I(\c0.n33607 ));
    CascadeMux I__22552 (
            .O(N__93810),
            .I(N__93807));
    InMux I__22551 (
            .O(N__93807),
            .I(N__93804));
    LocalMux I__22550 (
            .O(N__93804),
            .I(N__93800));
    CascadeMux I__22549 (
            .O(N__93803),
            .I(N__93797));
    Span4Mux_v I__22548 (
            .O(N__93800),
            .I(N__93794));
    InMux I__22547 (
            .O(N__93797),
            .I(N__93791));
    Span4Mux_h I__22546 (
            .O(N__93794),
            .I(N__93788));
    LocalMux I__22545 (
            .O(N__93791),
            .I(\c0.n33379 ));
    Odrv4 I__22544 (
            .O(N__93788),
            .I(\c0.n33379 ));
    InMux I__22543 (
            .O(N__93783),
            .I(N__93779));
    InMux I__22542 (
            .O(N__93782),
            .I(N__93776));
    LocalMux I__22541 (
            .O(N__93779),
            .I(N__93770));
    LocalMux I__22540 (
            .O(N__93776),
            .I(N__93770));
    InMux I__22539 (
            .O(N__93775),
            .I(N__93767));
    Span4Mux_v I__22538 (
            .O(N__93770),
            .I(N__93762));
    LocalMux I__22537 (
            .O(N__93767),
            .I(N__93762));
    Odrv4 I__22536 (
            .O(N__93762),
            .I(\quad_counter1.n2316 ));
    InMux I__22535 (
            .O(N__93759),
            .I(\quad_counter1.n30491 ));
    InMux I__22534 (
            .O(N__93756),
            .I(N__93752));
    InMux I__22533 (
            .O(N__93755),
            .I(N__93749));
    LocalMux I__22532 (
            .O(N__93752),
            .I(N__93743));
    LocalMux I__22531 (
            .O(N__93749),
            .I(N__93743));
    InMux I__22530 (
            .O(N__93748),
            .I(N__93740));
    Span4Mux_v I__22529 (
            .O(N__93743),
            .I(N__93735));
    LocalMux I__22528 (
            .O(N__93740),
            .I(N__93735));
    Odrv4 I__22527 (
            .O(N__93735),
            .I(\quad_counter1.n2315 ));
    InMux I__22526 (
            .O(N__93732),
            .I(\quad_counter1.n30492 ));
    InMux I__22525 (
            .O(N__93729),
            .I(N__93725));
    InMux I__22524 (
            .O(N__93728),
            .I(N__93722));
    LocalMux I__22523 (
            .O(N__93725),
            .I(N__93716));
    LocalMux I__22522 (
            .O(N__93722),
            .I(N__93716));
    InMux I__22521 (
            .O(N__93721),
            .I(N__93713));
    Span4Mux_v I__22520 (
            .O(N__93716),
            .I(N__93708));
    LocalMux I__22519 (
            .O(N__93713),
            .I(N__93708));
    Odrv4 I__22518 (
            .O(N__93708),
            .I(\quad_counter1.n2314 ));
    InMux I__22517 (
            .O(N__93705),
            .I(\quad_counter1.n30493 ));
    CascadeMux I__22516 (
            .O(N__93702),
            .I(N__93694));
    CascadeMux I__22515 (
            .O(N__93701),
            .I(N__93691));
    CascadeMux I__22514 (
            .O(N__93700),
            .I(N__93688));
    CascadeMux I__22513 (
            .O(N__93699),
            .I(N__93685));
    CascadeMux I__22512 (
            .O(N__93698),
            .I(N__93682));
    CascadeMux I__22511 (
            .O(N__93697),
            .I(N__93679));
    InMux I__22510 (
            .O(N__93694),
            .I(N__93674));
    InMux I__22509 (
            .O(N__93691),
            .I(N__93674));
    InMux I__22508 (
            .O(N__93688),
            .I(N__93665));
    InMux I__22507 (
            .O(N__93685),
            .I(N__93665));
    InMux I__22506 (
            .O(N__93682),
            .I(N__93665));
    InMux I__22505 (
            .O(N__93679),
            .I(N__93665));
    LocalMux I__22504 (
            .O(N__93674),
            .I(\quad_counter1.n36136 ));
    LocalMux I__22503 (
            .O(N__93665),
            .I(\quad_counter1.n36136 ));
    InMux I__22502 (
            .O(N__93660),
            .I(N__93657));
    LocalMux I__22501 (
            .O(N__93657),
            .I(N__93653));
    InMux I__22500 (
            .O(N__93656),
            .I(N__93650));
    Span4Mux_v I__22499 (
            .O(N__93653),
            .I(N__93646));
    LocalMux I__22498 (
            .O(N__93650),
            .I(N__93643));
    InMux I__22497 (
            .O(N__93649),
            .I(N__93640));
    Span4Mux_h I__22496 (
            .O(N__93646),
            .I(N__93635));
    Span4Mux_v I__22495 (
            .O(N__93643),
            .I(N__93635));
    LocalMux I__22494 (
            .O(N__93640),
            .I(N__93632));
    Odrv4 I__22493 (
            .O(N__93635),
            .I(\quad_counter1.n2313 ));
    Odrv4 I__22492 (
            .O(N__93632),
            .I(\quad_counter1.n2313 ));
    InMux I__22491 (
            .O(N__93627),
            .I(\quad_counter1.n30494 ));
    InMux I__22490 (
            .O(N__93624),
            .I(\quad_counter1.n30495 ));
    InMux I__22489 (
            .O(N__93621),
            .I(N__93616));
    InMux I__22488 (
            .O(N__93620),
            .I(N__93613));
    InMux I__22487 (
            .O(N__93619),
            .I(N__93610));
    LocalMux I__22486 (
            .O(N__93616),
            .I(N__93603));
    LocalMux I__22485 (
            .O(N__93613),
            .I(N__93603));
    LocalMux I__22484 (
            .O(N__93610),
            .I(N__93603));
    Span4Mux_v I__22483 (
            .O(N__93603),
            .I(N__93600));
    Span4Mux_h I__22482 (
            .O(N__93600),
            .I(N__93597));
    Odrv4 I__22481 (
            .O(N__93597),
            .I(\quad_counter1.n2311 ));
    InMux I__22480 (
            .O(N__93594),
            .I(bfn_26_12_0_));
    InMux I__22479 (
            .O(N__93591),
            .I(N__93586));
    InMux I__22478 (
            .O(N__93590),
            .I(N__93583));
    InMux I__22477 (
            .O(N__93589),
            .I(N__93580));
    LocalMux I__22476 (
            .O(N__93586),
            .I(N__93573));
    LocalMux I__22475 (
            .O(N__93583),
            .I(N__93573));
    LocalMux I__22474 (
            .O(N__93580),
            .I(N__93573));
    Span4Mux_v I__22473 (
            .O(N__93573),
            .I(N__93570));
    Odrv4 I__22472 (
            .O(N__93570),
            .I(\quad_counter1.n2310 ));
    InMux I__22471 (
            .O(N__93567),
            .I(\quad_counter1.n30497 ));
    CascadeMux I__22470 (
            .O(N__93564),
            .I(N__93559));
    CascadeMux I__22469 (
            .O(N__93563),
            .I(N__93556));
    CascadeMux I__22468 (
            .O(N__93562),
            .I(N__93553));
    InMux I__22467 (
            .O(N__93559),
            .I(N__93548));
    InMux I__22466 (
            .O(N__93556),
            .I(N__93543));
    InMux I__22465 (
            .O(N__93553),
            .I(N__93543));
    CascadeMux I__22464 (
            .O(N__93552),
            .I(N__93540));
    CascadeMux I__22463 (
            .O(N__93551),
            .I(N__93537));
    LocalMux I__22462 (
            .O(N__93548),
            .I(N__93532));
    LocalMux I__22461 (
            .O(N__93543),
            .I(N__93532));
    InMux I__22460 (
            .O(N__93540),
            .I(N__93527));
    InMux I__22459 (
            .O(N__93537),
            .I(N__93527));
    Odrv4 I__22458 (
            .O(N__93532),
            .I(\quad_counter1.n2243 ));
    LocalMux I__22457 (
            .O(N__93527),
            .I(\quad_counter1.n2243 ));
    InMux I__22456 (
            .O(N__93522),
            .I(\quad_counter1.n30498 ));
    InMux I__22455 (
            .O(N__93519),
            .I(\quad_counter1.n30471 ));
    CascadeMux I__22454 (
            .O(N__93516),
            .I(\quad_counter1.n28279_cascade_ ));
    CascadeMux I__22453 (
            .O(N__93513),
            .I(\quad_counter1.n10_adj_4435_cascade_ ));
    CascadeMux I__22452 (
            .O(N__93510),
            .I(\quad_counter1.n7_adj_4436_cascade_ ));
    CascadeMux I__22451 (
            .O(N__93507),
            .I(\quad_counter1.n2243_cascade_ ));
    InMux I__22450 (
            .O(N__93504),
            .I(N__93499));
    InMux I__22449 (
            .O(N__93503),
            .I(N__93496));
    InMux I__22448 (
            .O(N__93502),
            .I(N__93493));
    LocalMux I__22447 (
            .O(N__93499),
            .I(N__93486));
    LocalMux I__22446 (
            .O(N__93496),
            .I(N__93486));
    LocalMux I__22445 (
            .O(N__93493),
            .I(N__93486));
    Span4Mux_v I__22444 (
            .O(N__93486),
            .I(N__93482));
    InMux I__22443 (
            .O(N__93485),
            .I(N__93479));
    Span4Mux_h I__22442 (
            .O(N__93482),
            .I(N__93476));
    LocalMux I__22441 (
            .O(N__93479),
            .I(\quad_counter1.millisecond_counter_21 ));
    Odrv4 I__22440 (
            .O(N__93476),
            .I(\quad_counter1.millisecond_counter_21 ));
    InMux I__22439 (
            .O(N__93471),
            .I(N__93467));
    InMux I__22438 (
            .O(N__93470),
            .I(N__93464));
    LocalMux I__22437 (
            .O(N__93467),
            .I(N__93458));
    LocalMux I__22436 (
            .O(N__93464),
            .I(N__93458));
    InMux I__22435 (
            .O(N__93463),
            .I(N__93455));
    Span4Mux_h I__22434 (
            .O(N__93458),
            .I(N__93452));
    LocalMux I__22433 (
            .O(N__93455),
            .I(N__93449));
    Odrv4 I__22432 (
            .O(N__93452),
            .I(\quad_counter1.n2319 ));
    Odrv12 I__22431 (
            .O(N__93449),
            .I(\quad_counter1.n2319 ));
    InMux I__22430 (
            .O(N__93444),
            .I(bfn_26_11_0_));
    InMux I__22429 (
            .O(N__93441),
            .I(N__93436));
    InMux I__22428 (
            .O(N__93440),
            .I(N__93433));
    InMux I__22427 (
            .O(N__93439),
            .I(N__93430));
    LocalMux I__22426 (
            .O(N__93436),
            .I(N__93425));
    LocalMux I__22425 (
            .O(N__93433),
            .I(N__93425));
    LocalMux I__22424 (
            .O(N__93430),
            .I(N__93422));
    Span4Mux_h I__22423 (
            .O(N__93425),
            .I(N__93419));
    Span4Mux_h I__22422 (
            .O(N__93422),
            .I(N__93416));
    Odrv4 I__22421 (
            .O(N__93419),
            .I(\quad_counter1.n2318 ));
    Odrv4 I__22420 (
            .O(N__93416),
            .I(\quad_counter1.n2318 ));
    InMux I__22419 (
            .O(N__93411),
            .I(\quad_counter1.n30489 ));
    InMux I__22418 (
            .O(N__93408),
            .I(N__93404));
    InMux I__22417 (
            .O(N__93407),
            .I(N__93401));
    LocalMux I__22416 (
            .O(N__93404),
            .I(N__93395));
    LocalMux I__22415 (
            .O(N__93401),
            .I(N__93395));
    InMux I__22414 (
            .O(N__93400),
            .I(N__93392));
    Span4Mux_v I__22413 (
            .O(N__93395),
            .I(N__93387));
    LocalMux I__22412 (
            .O(N__93392),
            .I(N__93387));
    Odrv4 I__22411 (
            .O(N__93387),
            .I(\quad_counter1.n2317 ));
    InMux I__22410 (
            .O(N__93384),
            .I(\quad_counter1.n30490 ));
    InMux I__22409 (
            .O(N__93381),
            .I(N__93376));
    InMux I__22408 (
            .O(N__93380),
            .I(N__93373));
    InMux I__22407 (
            .O(N__93379),
            .I(N__93370));
    LocalMux I__22406 (
            .O(N__93376),
            .I(N__93364));
    LocalMux I__22405 (
            .O(N__93373),
            .I(N__93364));
    LocalMux I__22404 (
            .O(N__93370),
            .I(N__93361));
    InMux I__22403 (
            .O(N__93369),
            .I(N__93358));
    Span4Mux_h I__22402 (
            .O(N__93364),
            .I(N__93355));
    Span4Mux_h I__22401 (
            .O(N__93361),
            .I(N__93352));
    LocalMux I__22400 (
            .O(N__93358),
            .I(\quad_counter1.millisecond_counter_30 ));
    Odrv4 I__22399 (
            .O(N__93355),
            .I(\quad_counter1.millisecond_counter_30 ));
    Odrv4 I__22398 (
            .O(N__93352),
            .I(\quad_counter1.millisecond_counter_30 ));
    InMux I__22397 (
            .O(N__93345),
            .I(\quad_counter1.n30463 ));
    InMux I__22396 (
            .O(N__93342),
            .I(N__93337));
    InMux I__22395 (
            .O(N__93341),
            .I(N__93334));
    InMux I__22394 (
            .O(N__93340),
            .I(N__93331));
    LocalMux I__22393 (
            .O(N__93337),
            .I(N__93325));
    LocalMux I__22392 (
            .O(N__93334),
            .I(N__93325));
    LocalMux I__22391 (
            .O(N__93331),
            .I(N__93322));
    InMux I__22390 (
            .O(N__93330),
            .I(N__93319));
    Span4Mux_h I__22389 (
            .O(N__93325),
            .I(N__93316));
    Span4Mux_h I__22388 (
            .O(N__93322),
            .I(N__93313));
    LocalMux I__22387 (
            .O(N__93319),
            .I(\quad_counter1.millisecond_counter_31 ));
    Odrv4 I__22386 (
            .O(N__93316),
            .I(\quad_counter1.millisecond_counter_31 ));
    Odrv4 I__22385 (
            .O(N__93313),
            .I(\quad_counter1.millisecond_counter_31 ));
    CascadeMux I__22384 (
            .O(N__93306),
            .I(N__93298));
    CascadeMux I__22383 (
            .O(N__93305),
            .I(N__93295));
    CascadeMux I__22382 (
            .O(N__93304),
            .I(N__93292));
    CascadeMux I__22381 (
            .O(N__93303),
            .I(N__93289));
    CascadeMux I__22380 (
            .O(N__93302),
            .I(N__93286));
    CascadeMux I__22379 (
            .O(N__93301),
            .I(N__93283));
    InMux I__22378 (
            .O(N__93298),
            .I(N__93278));
    InMux I__22377 (
            .O(N__93295),
            .I(N__93278));
    InMux I__22376 (
            .O(N__93292),
            .I(N__93269));
    InMux I__22375 (
            .O(N__93289),
            .I(N__93269));
    InMux I__22374 (
            .O(N__93286),
            .I(N__93269));
    InMux I__22373 (
            .O(N__93283),
            .I(N__93269));
    LocalMux I__22372 (
            .O(N__93278),
            .I(\quad_counter1.n36138 ));
    LocalMux I__22371 (
            .O(N__93269),
            .I(\quad_counter1.n36138 ));
    InMux I__22370 (
            .O(N__93264),
            .I(\quad_counter1.n30464 ));
    InMux I__22369 (
            .O(N__93261),
            .I(bfn_26_9_0_));
    InMux I__22368 (
            .O(N__93258),
            .I(\quad_counter1.n30465 ));
    InMux I__22367 (
            .O(N__93255),
            .I(\quad_counter1.n30466 ));
    InMux I__22366 (
            .O(N__93252),
            .I(\quad_counter1.n30467 ));
    InMux I__22365 (
            .O(N__93249),
            .I(\quad_counter1.n30468 ));
    InMux I__22364 (
            .O(N__93246),
            .I(\quad_counter1.n30469 ));
    InMux I__22363 (
            .O(N__93243),
            .I(\quad_counter1.n30470 ));
    CascadeMux I__22362 (
            .O(N__93240),
            .I(\quad_counter1.n10_adj_4430_cascade_ ));
    CascadeMux I__22361 (
            .O(N__93237),
            .I(\quad_counter1.n1847_cascade_ ));
    CascadeMux I__22360 (
            .O(N__93234),
            .I(N__93231));
    InMux I__22359 (
            .O(N__93231),
            .I(N__93228));
    LocalMux I__22358 (
            .O(N__93228),
            .I(N__93220));
    InMux I__22357 (
            .O(N__93227),
            .I(N__93216));
    InMux I__22356 (
            .O(N__93226),
            .I(N__93209));
    InMux I__22355 (
            .O(N__93225),
            .I(N__93209));
    InMux I__22354 (
            .O(N__93224),
            .I(N__93209));
    InMux I__22353 (
            .O(N__93223),
            .I(N__93206));
    Span4Mux_v I__22352 (
            .O(N__93220),
            .I(N__93203));
    InMux I__22351 (
            .O(N__93219),
            .I(N__93199));
    LocalMux I__22350 (
            .O(N__93216),
            .I(N__93195));
    LocalMux I__22349 (
            .O(N__93209),
            .I(N__93192));
    LocalMux I__22348 (
            .O(N__93206),
            .I(N__93189));
    Span4Mux_h I__22347 (
            .O(N__93203),
            .I(N__93186));
    InMux I__22346 (
            .O(N__93202),
            .I(N__93182));
    LocalMux I__22345 (
            .O(N__93199),
            .I(N__93179));
    InMux I__22344 (
            .O(N__93198),
            .I(N__93176));
    Span4Mux_h I__22343 (
            .O(N__93195),
            .I(N__93171));
    Span4Mux_h I__22342 (
            .O(N__93192),
            .I(N__93171));
    Span4Mux_v I__22341 (
            .O(N__93189),
            .I(N__93166));
    Span4Mux_h I__22340 (
            .O(N__93186),
            .I(N__93166));
    InMux I__22339 (
            .O(N__93185),
            .I(N__93163));
    LocalMux I__22338 (
            .O(N__93182),
            .I(N__93160));
    Span4Mux_h I__22337 (
            .O(N__93179),
            .I(N__93155));
    LocalMux I__22336 (
            .O(N__93176),
            .I(N__93155));
    Sp12to4 I__22335 (
            .O(N__93171),
            .I(N__93152));
    Span4Mux_v I__22334 (
            .O(N__93166),
            .I(N__93149));
    LocalMux I__22333 (
            .O(N__93163),
            .I(N__93146));
    Span12Mux_h I__22332 (
            .O(N__93160),
            .I(N__93143));
    Sp12to4 I__22331 (
            .O(N__93155),
            .I(N__93134));
    Span12Mux_v I__22330 (
            .O(N__93152),
            .I(N__93134));
    Sp12to4 I__22329 (
            .O(N__93149),
            .I(N__93134));
    Span12Mux_h I__22328 (
            .O(N__93146),
            .I(N__93134));
    Span12Mux_v I__22327 (
            .O(N__93143),
            .I(N__93130));
    Span12Mux_v I__22326 (
            .O(N__93134),
            .I(N__93127));
    InMux I__22325 (
            .O(N__93133),
            .I(N__93124));
    Odrv12 I__22324 (
            .O(N__93130),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv12 I__22323 (
            .O(N__93127),
            .I(\c0.FRAME_MATCHER_i_0 ));
    LocalMux I__22322 (
            .O(N__93124),
            .I(\c0.FRAME_MATCHER_i_0 ));
    SRMux I__22321 (
            .O(N__93117),
            .I(N__93114));
    LocalMux I__22320 (
            .O(N__93114),
            .I(N__93111));
    Span12Mux_s6_v I__22319 (
            .O(N__93111),
            .I(N__93108));
    Odrv12 I__22318 (
            .O(N__93108),
            .I(\c0.n3 ));
    InMux I__22317 (
            .O(N__93105),
            .I(N__93100));
    InMux I__22316 (
            .O(N__93104),
            .I(N__93097));
    InMux I__22315 (
            .O(N__93103),
            .I(N__93094));
    LocalMux I__22314 (
            .O(N__93100),
            .I(N__93088));
    LocalMux I__22313 (
            .O(N__93097),
            .I(N__93088));
    LocalMux I__22312 (
            .O(N__93094),
            .I(N__93085));
    InMux I__22311 (
            .O(N__93093),
            .I(N__93082));
    Span4Mux_h I__22310 (
            .O(N__93088),
            .I(N__93079));
    Span4Mux_h I__22309 (
            .O(N__93085),
            .I(N__93076));
    LocalMux I__22308 (
            .O(N__93082),
            .I(\quad_counter1.millisecond_counter_25 ));
    Odrv4 I__22307 (
            .O(N__93079),
            .I(\quad_counter1.millisecond_counter_25 ));
    Odrv4 I__22306 (
            .O(N__93076),
            .I(\quad_counter1.millisecond_counter_25 ));
    InMux I__22305 (
            .O(N__93069),
            .I(bfn_26_8_0_));
    InMux I__22304 (
            .O(N__93066),
            .I(N__93061));
    InMux I__22303 (
            .O(N__93065),
            .I(N__93058));
    InMux I__22302 (
            .O(N__93064),
            .I(N__93055));
    LocalMux I__22301 (
            .O(N__93061),
            .I(N__93047));
    LocalMux I__22300 (
            .O(N__93058),
            .I(N__93047));
    LocalMux I__22299 (
            .O(N__93055),
            .I(N__93047));
    InMux I__22298 (
            .O(N__93054),
            .I(N__93044));
    Span4Mux_v I__22297 (
            .O(N__93047),
            .I(N__93041));
    LocalMux I__22296 (
            .O(N__93044),
            .I(\quad_counter1.millisecond_counter_26 ));
    Odrv4 I__22295 (
            .O(N__93041),
            .I(\quad_counter1.millisecond_counter_26 ));
    CascadeMux I__22294 (
            .O(N__93036),
            .I(N__93033));
    InMux I__22293 (
            .O(N__93033),
            .I(N__93030));
    LocalMux I__22292 (
            .O(N__93030),
            .I(\quad_counter1.n1847 ));
    InMux I__22291 (
            .O(N__93027),
            .I(\quad_counter1.n30459 ));
    InMux I__22290 (
            .O(N__93024),
            .I(N__93019));
    InMux I__22289 (
            .O(N__93023),
            .I(N__93016));
    InMux I__22288 (
            .O(N__93022),
            .I(N__93013));
    LocalMux I__22287 (
            .O(N__93019),
            .I(N__93007));
    LocalMux I__22286 (
            .O(N__93016),
            .I(N__93007));
    LocalMux I__22285 (
            .O(N__93013),
            .I(N__93004));
    InMux I__22284 (
            .O(N__93012),
            .I(N__93001));
    Span4Mux_v I__22283 (
            .O(N__93007),
            .I(N__92998));
    Span4Mux_h I__22282 (
            .O(N__93004),
            .I(N__92995));
    LocalMux I__22281 (
            .O(N__93001),
            .I(\quad_counter1.millisecond_counter_27 ));
    Odrv4 I__22280 (
            .O(N__92998),
            .I(\quad_counter1.millisecond_counter_27 ));
    Odrv4 I__22279 (
            .O(N__92995),
            .I(\quad_counter1.millisecond_counter_27 ));
    InMux I__22278 (
            .O(N__92988),
            .I(\quad_counter1.n30460 ));
    InMux I__22277 (
            .O(N__92985),
            .I(N__92980));
    InMux I__22276 (
            .O(N__92984),
            .I(N__92977));
    InMux I__22275 (
            .O(N__92983),
            .I(N__92974));
    LocalMux I__22274 (
            .O(N__92980),
            .I(N__92966));
    LocalMux I__22273 (
            .O(N__92977),
            .I(N__92966));
    LocalMux I__22272 (
            .O(N__92974),
            .I(N__92966));
    InMux I__22271 (
            .O(N__92973),
            .I(N__92963));
    Span4Mux_v I__22270 (
            .O(N__92966),
            .I(N__92960));
    LocalMux I__22269 (
            .O(N__92963),
            .I(\quad_counter1.millisecond_counter_28 ));
    Odrv4 I__22268 (
            .O(N__92960),
            .I(\quad_counter1.millisecond_counter_28 ));
    InMux I__22267 (
            .O(N__92955),
            .I(\quad_counter1.n30461 ));
    CascadeMux I__22266 (
            .O(N__92952),
            .I(N__92947));
    InMux I__22265 (
            .O(N__92951),
            .I(N__92944));
    InMux I__22264 (
            .O(N__92950),
            .I(N__92941));
    InMux I__22263 (
            .O(N__92947),
            .I(N__92938));
    LocalMux I__22262 (
            .O(N__92944),
            .I(N__92930));
    LocalMux I__22261 (
            .O(N__92941),
            .I(N__92930));
    LocalMux I__22260 (
            .O(N__92938),
            .I(N__92930));
    InMux I__22259 (
            .O(N__92937),
            .I(N__92927));
    Span4Mux_v I__22258 (
            .O(N__92930),
            .I(N__92924));
    LocalMux I__22257 (
            .O(N__92927),
            .I(\quad_counter1.millisecond_counter_29 ));
    Odrv4 I__22256 (
            .O(N__92924),
            .I(\quad_counter1.millisecond_counter_29 ));
    InMux I__22255 (
            .O(N__92919),
            .I(\quad_counter1.n30462 ));
    InMux I__22254 (
            .O(N__92916),
            .I(N__92911));
    InMux I__22253 (
            .O(N__92915),
            .I(N__92908));
    InMux I__22252 (
            .O(N__92914),
            .I(N__92905));
    LocalMux I__22251 (
            .O(N__92911),
            .I(N__92887));
    LocalMux I__22250 (
            .O(N__92908),
            .I(N__92887));
    LocalMux I__22249 (
            .O(N__92905),
            .I(N__92887));
    InMux I__22248 (
            .O(N__92904),
            .I(N__92884));
    InMux I__22247 (
            .O(N__92903),
            .I(N__92881));
    InMux I__22246 (
            .O(N__92902),
            .I(N__92878));
    InMux I__22245 (
            .O(N__92901),
            .I(N__92867));
    InMux I__22244 (
            .O(N__92900),
            .I(N__92861));
    InMux I__22243 (
            .O(N__92899),
            .I(N__92858));
    InMux I__22242 (
            .O(N__92898),
            .I(N__92855));
    InMux I__22241 (
            .O(N__92897),
            .I(N__92852));
    InMux I__22240 (
            .O(N__92896),
            .I(N__92849));
    InMux I__22239 (
            .O(N__92895),
            .I(N__92846));
    InMux I__22238 (
            .O(N__92894),
            .I(N__92834));
    Span4Mux_v I__22237 (
            .O(N__92887),
            .I(N__92831));
    LocalMux I__22236 (
            .O(N__92884),
            .I(N__92826));
    LocalMux I__22235 (
            .O(N__92881),
            .I(N__92826));
    LocalMux I__22234 (
            .O(N__92878),
            .I(N__92823));
    InMux I__22233 (
            .O(N__92877),
            .I(N__92820));
    InMux I__22232 (
            .O(N__92876),
            .I(N__92817));
    InMux I__22231 (
            .O(N__92875),
            .I(N__92814));
    InMux I__22230 (
            .O(N__92874),
            .I(N__92811));
    InMux I__22229 (
            .O(N__92873),
            .I(N__92808));
    InMux I__22228 (
            .O(N__92872),
            .I(N__92805));
    InMux I__22227 (
            .O(N__92871),
            .I(N__92802));
    InMux I__22226 (
            .O(N__92870),
            .I(N__92799));
    LocalMux I__22225 (
            .O(N__92867),
            .I(N__92796));
    InMux I__22224 (
            .O(N__92866),
            .I(N__92793));
    InMux I__22223 (
            .O(N__92865),
            .I(N__92790));
    InMux I__22222 (
            .O(N__92864),
            .I(N__92787));
    LocalMux I__22221 (
            .O(N__92861),
            .I(N__92778));
    LocalMux I__22220 (
            .O(N__92858),
            .I(N__92778));
    LocalMux I__22219 (
            .O(N__92855),
            .I(N__92778));
    LocalMux I__22218 (
            .O(N__92852),
            .I(N__92778));
    LocalMux I__22217 (
            .O(N__92849),
            .I(N__92775));
    LocalMux I__22216 (
            .O(N__92846),
            .I(N__92772));
    InMux I__22215 (
            .O(N__92845),
            .I(N__92769));
    InMux I__22214 (
            .O(N__92844),
            .I(N__92766));
    InMux I__22213 (
            .O(N__92843),
            .I(N__92763));
    InMux I__22212 (
            .O(N__92842),
            .I(N__92760));
    InMux I__22211 (
            .O(N__92841),
            .I(N__92757));
    InMux I__22210 (
            .O(N__92840),
            .I(N__92754));
    InMux I__22209 (
            .O(N__92839),
            .I(N__92751));
    InMux I__22208 (
            .O(N__92838),
            .I(N__92747));
    InMux I__22207 (
            .O(N__92837),
            .I(N__92744));
    LocalMux I__22206 (
            .O(N__92834),
            .I(N__92735));
    Span4Mux_v I__22205 (
            .O(N__92831),
            .I(N__92735));
    Span4Mux_v I__22204 (
            .O(N__92826),
            .I(N__92735));
    Span4Mux_v I__22203 (
            .O(N__92823),
            .I(N__92735));
    LocalMux I__22202 (
            .O(N__92820),
            .I(N__92724));
    LocalMux I__22201 (
            .O(N__92817),
            .I(N__92724));
    LocalMux I__22200 (
            .O(N__92814),
            .I(N__92724));
    LocalMux I__22199 (
            .O(N__92811),
            .I(N__92724));
    LocalMux I__22198 (
            .O(N__92808),
            .I(N__92724));
    LocalMux I__22197 (
            .O(N__92805),
            .I(N__92707));
    LocalMux I__22196 (
            .O(N__92802),
            .I(N__92707));
    LocalMux I__22195 (
            .O(N__92799),
            .I(N__92707));
    Sp12to4 I__22194 (
            .O(N__92796),
            .I(N__92707));
    LocalMux I__22193 (
            .O(N__92793),
            .I(N__92707));
    LocalMux I__22192 (
            .O(N__92790),
            .I(N__92707));
    LocalMux I__22191 (
            .O(N__92787),
            .I(N__92707));
    Sp12to4 I__22190 (
            .O(N__92778),
            .I(N__92707));
    Span4Mux_v I__22189 (
            .O(N__92775),
            .I(N__92702));
    Span4Mux_v I__22188 (
            .O(N__92772),
            .I(N__92702));
    LocalMux I__22187 (
            .O(N__92769),
            .I(N__92687));
    LocalMux I__22186 (
            .O(N__92766),
            .I(N__92687));
    LocalMux I__22185 (
            .O(N__92763),
            .I(N__92687));
    LocalMux I__22184 (
            .O(N__92760),
            .I(N__92687));
    LocalMux I__22183 (
            .O(N__92757),
            .I(N__92687));
    LocalMux I__22182 (
            .O(N__92754),
            .I(N__92687));
    LocalMux I__22181 (
            .O(N__92751),
            .I(N__92687));
    InMux I__22180 (
            .O(N__92750),
            .I(N__92684));
    LocalMux I__22179 (
            .O(N__92747),
            .I(N__92681));
    LocalMux I__22178 (
            .O(N__92744),
            .I(N__92675));
    Sp12to4 I__22177 (
            .O(N__92735),
            .I(N__92670));
    Span12Mux_s9_v I__22176 (
            .O(N__92724),
            .I(N__92670));
    Span12Mux_s10_v I__22175 (
            .O(N__92707),
            .I(N__92661));
    Sp12to4 I__22174 (
            .O(N__92702),
            .I(N__92661));
    Span12Mux_v I__22173 (
            .O(N__92687),
            .I(N__92661));
    LocalMux I__22172 (
            .O(N__92684),
            .I(N__92661));
    Span4Mux_v I__22171 (
            .O(N__92681),
            .I(N__92658));
    InMux I__22170 (
            .O(N__92680),
            .I(N__92655));
    InMux I__22169 (
            .O(N__92679),
            .I(N__92650));
    InMux I__22168 (
            .O(N__92678),
            .I(N__92650));
    Span4Mux_v I__22167 (
            .O(N__92675),
            .I(N__92647));
    Span12Mux_h I__22166 (
            .O(N__92670),
            .I(N__92642));
    Span12Mux_h I__22165 (
            .O(N__92661),
            .I(N__92642));
    Span4Mux_h I__22164 (
            .O(N__92658),
            .I(N__92637));
    LocalMux I__22163 (
            .O(N__92655),
            .I(N__92637));
    LocalMux I__22162 (
            .O(N__92650),
            .I(N__92634));
    Odrv4 I__22161 (
            .O(N__92647),
            .I(\c0.n1286 ));
    Odrv12 I__22160 (
            .O(N__92642),
            .I(\c0.n1286 ));
    Odrv4 I__22159 (
            .O(N__92637),
            .I(\c0.n1286 ));
    Odrv4 I__22158 (
            .O(N__92634),
            .I(\c0.n1286 ));
    InMux I__22157 (
            .O(N__92625),
            .I(bfn_24_32_0_));
    InMux I__22156 (
            .O(N__92622),
            .I(N__92619));
    LocalMux I__22155 (
            .O(N__92619),
            .I(N__92610));
    InMux I__22154 (
            .O(N__92618),
            .I(N__92607));
    CascadeMux I__22153 (
            .O(N__92617),
            .I(N__92604));
    CascadeMux I__22152 (
            .O(N__92616),
            .I(N__92601));
    CascadeMux I__22151 (
            .O(N__92615),
            .I(N__92596));
    InMux I__22150 (
            .O(N__92614),
            .I(N__92591));
    InMux I__22149 (
            .O(N__92613),
            .I(N__92591));
    Span4Mux_v I__22148 (
            .O(N__92610),
            .I(N__92586));
    LocalMux I__22147 (
            .O(N__92607),
            .I(N__92586));
    InMux I__22146 (
            .O(N__92604),
            .I(N__92583));
    InMux I__22145 (
            .O(N__92601),
            .I(N__92580));
    InMux I__22144 (
            .O(N__92600),
            .I(N__92577));
    InMux I__22143 (
            .O(N__92599),
            .I(N__92574));
    InMux I__22142 (
            .O(N__92596),
            .I(N__92571));
    LocalMux I__22141 (
            .O(N__92591),
            .I(N__92564));
    Span4Mux_h I__22140 (
            .O(N__92586),
            .I(N__92564));
    LocalMux I__22139 (
            .O(N__92583),
            .I(N__92564));
    LocalMux I__22138 (
            .O(N__92580),
            .I(N__92561));
    LocalMux I__22137 (
            .O(N__92577),
            .I(N__92558));
    LocalMux I__22136 (
            .O(N__92574),
            .I(N__92555));
    LocalMux I__22135 (
            .O(N__92571),
            .I(N__92550));
    Span4Mux_v I__22134 (
            .O(N__92564),
            .I(N__92550));
    Span4Mux_v I__22133 (
            .O(N__92561),
            .I(N__92547));
    Span4Mux_v I__22132 (
            .O(N__92558),
            .I(N__92544));
    Span4Mux_h I__22131 (
            .O(N__92555),
            .I(N__92541));
    Span4Mux_v I__22130 (
            .O(N__92550),
            .I(N__92538));
    Span4Mux_v I__22129 (
            .O(N__92547),
            .I(N__92533));
    Span4Mux_v I__22128 (
            .O(N__92544),
            .I(N__92533));
    Span4Mux_h I__22127 (
            .O(N__92541),
            .I(N__92530));
    Sp12to4 I__22126 (
            .O(N__92538),
            .I(N__92525));
    Sp12to4 I__22125 (
            .O(N__92533),
            .I(N__92525));
    Sp12to4 I__22124 (
            .O(N__92530),
            .I(N__92518));
    Span12Mux_h I__22123 (
            .O(N__92525),
            .I(N__92518));
    InMux I__22122 (
            .O(N__92524),
            .I(N__92513));
    InMux I__22121 (
            .O(N__92523),
            .I(N__92513));
    Span12Mux_v I__22120 (
            .O(N__92518),
            .I(N__92510));
    LocalMux I__22119 (
            .O(N__92513),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv12 I__22118 (
            .O(N__92510),
            .I(\c0.FRAME_MATCHER_i_31 ));
    SRMux I__22117 (
            .O(N__92505),
            .I(N__92502));
    LocalMux I__22116 (
            .O(N__92502),
            .I(N__92499));
    Span4Mux_h I__22115 (
            .O(N__92499),
            .I(N__92496));
    Odrv4 I__22114 (
            .O(N__92496),
            .I(\c0.n3_adj_4610 ));
    InMux I__22113 (
            .O(N__92493),
            .I(N__92490));
    LocalMux I__22112 (
            .O(N__92490),
            .I(N__92486));
    InMux I__22111 (
            .O(N__92489),
            .I(N__92483));
    Span4Mux_v I__22110 (
            .O(N__92486),
            .I(N__92479));
    LocalMux I__22109 (
            .O(N__92483),
            .I(N__92476));
    InMux I__22108 (
            .O(N__92482),
            .I(N__92473));
    Span4Mux_v I__22107 (
            .O(N__92479),
            .I(N__92470));
    Odrv12 I__22106 (
            .O(N__92476),
            .I(\c0.FRAME_MATCHER_i_28 ));
    LocalMux I__22105 (
            .O(N__92473),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__22104 (
            .O(N__92470),
            .I(\c0.FRAME_MATCHER_i_28 ));
    SRMux I__22103 (
            .O(N__92463),
            .I(N__92460));
    LocalMux I__22102 (
            .O(N__92460),
            .I(N__92457));
    Odrv4 I__22101 (
            .O(N__92457),
            .I(\c0.n3_adj_4607 ));
    SRMux I__22100 (
            .O(N__92454),
            .I(N__92451));
    LocalMux I__22099 (
            .O(N__92451),
            .I(N__92448));
    Span4Mux_v I__22098 (
            .O(N__92448),
            .I(N__92445));
    Odrv4 I__22097 (
            .O(N__92445),
            .I(\c0.n3_adj_4608 ));
    InMux I__22096 (
            .O(N__92442),
            .I(bfn_24_31_0_));
    SRMux I__22095 (
            .O(N__92439),
            .I(N__92436));
    LocalMux I__22094 (
            .O(N__92436),
            .I(N__92433));
    Span4Mux_s2_v I__22093 (
            .O(N__92433),
            .I(N__92430));
    Odrv4 I__22092 (
            .O(N__92430),
            .I(\c0.n3_adj_4609 ));
    InMux I__22091 (
            .O(N__92427),
            .I(bfn_24_29_0_));
    InMux I__22090 (
            .O(N__92424),
            .I(N__92420));
    InMux I__22089 (
            .O(N__92423),
            .I(N__92417));
    LocalMux I__22088 (
            .O(N__92420),
            .I(N__92411));
    LocalMux I__22087 (
            .O(N__92417),
            .I(N__92411));
    InMux I__22086 (
            .O(N__92416),
            .I(N__92408));
    Sp12to4 I__22085 (
            .O(N__92411),
            .I(N__92405));
    LocalMux I__22084 (
            .O(N__92408),
            .I(\c0.FRAME_MATCHER_i_29 ));
    Odrv12 I__22083 (
            .O(N__92405),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__22082 (
            .O(N__92400),
            .I(bfn_24_30_0_));
    InMux I__22081 (
            .O(N__92397),
            .I(N__92394));
    LocalMux I__22080 (
            .O(N__92394),
            .I(N__92391));
    Span4Mux_h I__22079 (
            .O(N__92391),
            .I(N__92386));
    InMux I__22078 (
            .O(N__92390),
            .I(N__92383));
    InMux I__22077 (
            .O(N__92389),
            .I(N__92380));
    Span4Mux_v I__22076 (
            .O(N__92386),
            .I(N__92377));
    LocalMux I__22075 (
            .O(N__92383),
            .I(\c0.FRAME_MATCHER_i_27 ));
    LocalMux I__22074 (
            .O(N__92380),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv4 I__22073 (
            .O(N__92377),
            .I(\c0.FRAME_MATCHER_i_27 ));
    InMux I__22072 (
            .O(N__92370),
            .I(bfn_24_28_0_));
    SRMux I__22071 (
            .O(N__92367),
            .I(N__92364));
    LocalMux I__22070 (
            .O(N__92364),
            .I(N__92361));
    Odrv4 I__22069 (
            .O(N__92361),
            .I(\c0.n3_adj_4606 ));
    InMux I__22068 (
            .O(N__92358),
            .I(N__92355));
    LocalMux I__22067 (
            .O(N__92355),
            .I(N__92350));
    InMux I__22066 (
            .O(N__92354),
            .I(N__92347));
    InMux I__22065 (
            .O(N__92353),
            .I(N__92344));
    Span4Mux_v I__22064 (
            .O(N__92350),
            .I(N__92341));
    LocalMux I__22063 (
            .O(N__92347),
            .I(\c0.FRAME_MATCHER_i_26 ));
    LocalMux I__22062 (
            .O(N__92344),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__22061 (
            .O(N__92341),
            .I(\c0.FRAME_MATCHER_i_26 ));
    InMux I__22060 (
            .O(N__92334),
            .I(bfn_24_27_0_));
    SRMux I__22059 (
            .O(N__92331),
            .I(N__92328));
    LocalMux I__22058 (
            .O(N__92328),
            .I(N__92325));
    Odrv4 I__22057 (
            .O(N__92325),
            .I(\c0.n3_adj_4605 ));
    InMux I__22056 (
            .O(N__92322),
            .I(N__92319));
    LocalMux I__22055 (
            .O(N__92319),
            .I(N__92314));
    InMux I__22054 (
            .O(N__92318),
            .I(N__92311));
    InMux I__22053 (
            .O(N__92317),
            .I(N__92308));
    Sp12to4 I__22052 (
            .O(N__92314),
            .I(N__92305));
    LocalMux I__22051 (
            .O(N__92311),
            .I(\c0.FRAME_MATCHER_i_25 ));
    LocalMux I__22050 (
            .O(N__92308),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv12 I__22049 (
            .O(N__92305),
            .I(\c0.FRAME_MATCHER_i_25 ));
    InMux I__22048 (
            .O(N__92298),
            .I(bfn_24_26_0_));
    SRMux I__22047 (
            .O(N__92295),
            .I(N__92292));
    LocalMux I__22046 (
            .O(N__92292),
            .I(\c0.n3_adj_4604 ));
    InMux I__22045 (
            .O(N__92289),
            .I(bfn_24_25_0_));
    SRMux I__22044 (
            .O(N__92286),
            .I(N__92283));
    LocalMux I__22043 (
            .O(N__92283),
            .I(N__92280));
    Span4Mux_h I__22042 (
            .O(N__92280),
            .I(N__92277));
    Odrv4 I__22041 (
            .O(N__92277),
            .I(\c0.n3_adj_4603 ));
    InMux I__22040 (
            .O(N__92274),
            .I(N__92269));
    InMux I__22039 (
            .O(N__92273),
            .I(N__92266));
    InMux I__22038 (
            .O(N__92272),
            .I(N__92263));
    LocalMux I__22037 (
            .O(N__92269),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__22036 (
            .O(N__92266),
            .I(\c0.FRAME_MATCHER_i_23 ));
    LocalMux I__22035 (
            .O(N__92263),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__22034 (
            .O(N__92256),
            .I(bfn_24_24_0_));
    SRMux I__22033 (
            .O(N__92253),
            .I(N__92250));
    LocalMux I__22032 (
            .O(N__92250),
            .I(N__92247));
    Span4Mux_v I__22031 (
            .O(N__92247),
            .I(N__92244));
    Odrv4 I__22030 (
            .O(N__92244),
            .I(\c0.n3_adj_4602 ));
    InMux I__22029 (
            .O(N__92241),
            .I(N__92236));
    InMux I__22028 (
            .O(N__92240),
            .I(N__92233));
    InMux I__22027 (
            .O(N__92239),
            .I(N__92230));
    LocalMux I__22026 (
            .O(N__92236),
            .I(N__92227));
    LocalMux I__22025 (
            .O(N__92233),
            .I(\c0.FRAME_MATCHER_i_22 ));
    LocalMux I__22024 (
            .O(N__92230),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__22023 (
            .O(N__92227),
            .I(\c0.FRAME_MATCHER_i_22 ));
    InMux I__22022 (
            .O(N__92220),
            .I(bfn_24_23_0_));
    SRMux I__22021 (
            .O(N__92217),
            .I(N__92214));
    LocalMux I__22020 (
            .O(N__92214),
            .I(N__92211));
    Odrv4 I__22019 (
            .O(N__92211),
            .I(\c0.n3_adj_4601 ));
    InMux I__22018 (
            .O(N__92208),
            .I(bfn_24_22_0_));
    SRMux I__22017 (
            .O(N__92205),
            .I(N__92202));
    LocalMux I__22016 (
            .O(N__92202),
            .I(N__92199));
    Odrv4 I__22015 (
            .O(N__92199),
            .I(\c0.n3_adj_4598 ));
    InMux I__22014 (
            .O(N__92196),
            .I(N__92191));
    InMux I__22013 (
            .O(N__92195),
            .I(N__92186));
    InMux I__22012 (
            .O(N__92194),
            .I(N__92186));
    LocalMux I__22011 (
            .O(N__92191),
            .I(\c0.FRAME_MATCHER_i_20 ));
    LocalMux I__22010 (
            .O(N__92186),
            .I(\c0.FRAME_MATCHER_i_20 ));
    InMux I__22009 (
            .O(N__92181),
            .I(bfn_24_21_0_));
    SRMux I__22008 (
            .O(N__92178),
            .I(N__92175));
    LocalMux I__22007 (
            .O(N__92175),
            .I(N__92172));
    Span4Mux_h I__22006 (
            .O(N__92172),
            .I(N__92169));
    Span4Mux_h I__22005 (
            .O(N__92169),
            .I(N__92166));
    Odrv4 I__22004 (
            .O(N__92166),
            .I(\c0.n3_adj_4599 ));
    InMux I__22003 (
            .O(N__92163),
            .I(N__92157));
    InMux I__22002 (
            .O(N__92162),
            .I(N__92157));
    LocalMux I__22001 (
            .O(N__92157),
            .I(N__92153));
    InMux I__22000 (
            .O(N__92156),
            .I(N__92150));
    Span4Mux_v I__21999 (
            .O(N__92153),
            .I(N__92147));
    LocalMux I__21998 (
            .O(N__92150),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__21997 (
            .O(N__92147),
            .I(\c0.FRAME_MATCHER_i_18 ));
    InMux I__21996 (
            .O(N__92142),
            .I(bfn_24_19_0_));
    SRMux I__21995 (
            .O(N__92139),
            .I(N__92136));
    LocalMux I__21994 (
            .O(N__92136),
            .I(N__92133));
    Span4Mux_v I__21993 (
            .O(N__92133),
            .I(N__92130));
    Odrv4 I__21992 (
            .O(N__92130),
            .I(\c0.n3_adj_4597 ));
    CascadeMux I__21991 (
            .O(N__92127),
            .I(N__92124));
    InMux I__21990 (
            .O(N__92124),
            .I(N__92121));
    LocalMux I__21989 (
            .O(N__92121),
            .I(N__92116));
    InMux I__21988 (
            .O(N__92120),
            .I(N__92113));
    InMux I__21987 (
            .O(N__92119),
            .I(N__92110));
    Span4Mux_h I__21986 (
            .O(N__92116),
            .I(N__92107));
    LocalMux I__21985 (
            .O(N__92113),
            .I(\c0.FRAME_MATCHER_i_19 ));
    LocalMux I__21984 (
            .O(N__92110),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv4 I__21983 (
            .O(N__92107),
            .I(\c0.FRAME_MATCHER_i_19 ));
    InMux I__21982 (
            .O(N__92100),
            .I(bfn_24_20_0_));
    InMux I__21981 (
            .O(N__92097),
            .I(bfn_24_18_0_));
    InMux I__21980 (
            .O(N__92094),
            .I(N__92090));
    CascadeMux I__21979 (
            .O(N__92093),
            .I(N__92087));
    LocalMux I__21978 (
            .O(N__92090),
            .I(N__92084));
    InMux I__21977 (
            .O(N__92087),
            .I(N__92081));
    Span4Mux_h I__21976 (
            .O(N__92084),
            .I(N__92075));
    LocalMux I__21975 (
            .O(N__92081),
            .I(N__92075));
    InMux I__21974 (
            .O(N__92080),
            .I(N__92072));
    Span4Mux_v I__21973 (
            .O(N__92075),
            .I(N__92069));
    LocalMux I__21972 (
            .O(N__92072),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__21971 (
            .O(N__92069),
            .I(\c0.FRAME_MATCHER_i_16 ));
    InMux I__21970 (
            .O(N__92064),
            .I(bfn_24_17_0_));
    SRMux I__21969 (
            .O(N__92061),
            .I(N__92058));
    LocalMux I__21968 (
            .O(N__92058),
            .I(N__92055));
    Span4Mux_h I__21967 (
            .O(N__92055),
            .I(N__92052));
    Odrv4 I__21966 (
            .O(N__92052),
            .I(\c0.n3_adj_4595 ));
    InMux I__21965 (
            .O(N__92049),
            .I(N__92045));
    InMux I__21964 (
            .O(N__92048),
            .I(N__92042));
    LocalMux I__21963 (
            .O(N__92045),
            .I(N__92038));
    LocalMux I__21962 (
            .O(N__92042),
            .I(N__92035));
    InMux I__21961 (
            .O(N__92041),
            .I(N__92032));
    Span4Mux_v I__21960 (
            .O(N__92038),
            .I(N__92029));
    Odrv4 I__21959 (
            .O(N__92035),
            .I(\c0.FRAME_MATCHER_i_15 ));
    LocalMux I__21958 (
            .O(N__92032),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__21957 (
            .O(N__92029),
            .I(\c0.FRAME_MATCHER_i_15 ));
    InMux I__21956 (
            .O(N__92022),
            .I(bfn_24_16_0_));
    SRMux I__21955 (
            .O(N__92019),
            .I(N__92016));
    LocalMux I__21954 (
            .O(N__92016),
            .I(N__92013));
    Odrv12 I__21953 (
            .O(N__92013),
            .I(\c0.n3_adj_4594 ));
    CascadeMux I__21952 (
            .O(N__92010),
            .I(N__92006));
    InMux I__21951 (
            .O(N__92009),
            .I(N__92003));
    InMux I__21950 (
            .O(N__92006),
            .I(N__92000));
    LocalMux I__21949 (
            .O(N__92003),
            .I(N__91994));
    LocalMux I__21948 (
            .O(N__92000),
            .I(N__91994));
    InMux I__21947 (
            .O(N__91999),
            .I(N__91991));
    Span4Mux_v I__21946 (
            .O(N__91994),
            .I(N__91988));
    LocalMux I__21945 (
            .O(N__91991),
            .I(\c0.FRAME_MATCHER_i_14 ));
    Odrv4 I__21944 (
            .O(N__91988),
            .I(\c0.FRAME_MATCHER_i_14 ));
    InMux I__21943 (
            .O(N__91983),
            .I(bfn_24_15_0_));
    SRMux I__21942 (
            .O(N__91980),
            .I(N__91977));
    LocalMux I__21941 (
            .O(N__91977),
            .I(N__91974));
    Span4Mux_v I__21940 (
            .O(N__91974),
            .I(N__91971));
    Odrv4 I__21939 (
            .O(N__91971),
            .I(\c0.n3_adj_4593 ));
    InMux I__21938 (
            .O(N__91968),
            .I(N__91964));
    InMux I__21937 (
            .O(N__91967),
            .I(N__91961));
    LocalMux I__21936 (
            .O(N__91964),
            .I(N__91955));
    LocalMux I__21935 (
            .O(N__91961),
            .I(N__91955));
    InMux I__21934 (
            .O(N__91960),
            .I(N__91952));
    Span4Mux_v I__21933 (
            .O(N__91955),
            .I(N__91949));
    LocalMux I__21932 (
            .O(N__91952),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv4 I__21931 (
            .O(N__91949),
            .I(\c0.FRAME_MATCHER_i_13 ));
    InMux I__21930 (
            .O(N__91944),
            .I(bfn_24_14_0_));
    SRMux I__21929 (
            .O(N__91941),
            .I(N__91938));
    LocalMux I__21928 (
            .O(N__91938),
            .I(N__91935));
    Span4Mux_h I__21927 (
            .O(N__91935),
            .I(N__91932));
    Odrv4 I__21926 (
            .O(N__91932),
            .I(\c0.n3_adj_4592 ));
    InMux I__21925 (
            .O(N__91929),
            .I(N__91925));
    InMux I__21924 (
            .O(N__91928),
            .I(N__91922));
    LocalMux I__21923 (
            .O(N__91925),
            .I(N__91917));
    LocalMux I__21922 (
            .O(N__91922),
            .I(N__91917));
    Span4Mux_v I__21921 (
            .O(N__91917),
            .I(N__91914));
    Span4Mux_v I__21920 (
            .O(N__91914),
            .I(N__91910));
    InMux I__21919 (
            .O(N__91913),
            .I(N__91907));
    Odrv4 I__21918 (
            .O(N__91910),
            .I(\c0.FRAME_MATCHER_i_12 ));
    LocalMux I__21917 (
            .O(N__91907),
            .I(\c0.FRAME_MATCHER_i_12 ));
    InMux I__21916 (
            .O(N__91902),
            .I(bfn_24_13_0_));
    SRMux I__21915 (
            .O(N__91899),
            .I(N__91896));
    LocalMux I__21914 (
            .O(N__91896),
            .I(N__91893));
    Span4Mux_v I__21913 (
            .O(N__91893),
            .I(N__91890));
    Odrv4 I__21912 (
            .O(N__91890),
            .I(\c0.n3_adj_4591 ));
    InMux I__21911 (
            .O(N__91887),
            .I(N__91883));
    InMux I__21910 (
            .O(N__91886),
            .I(N__91880));
    LocalMux I__21909 (
            .O(N__91883),
            .I(N__91874));
    LocalMux I__21908 (
            .O(N__91880),
            .I(N__91874));
    InMux I__21907 (
            .O(N__91879),
            .I(N__91871));
    Sp12to4 I__21906 (
            .O(N__91874),
            .I(N__91868));
    LocalMux I__21905 (
            .O(N__91871),
            .I(\c0.FRAME_MATCHER_i_11 ));
    Odrv12 I__21904 (
            .O(N__91868),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__21903 (
            .O(N__91863),
            .I(bfn_24_12_0_));
    SRMux I__21902 (
            .O(N__91860),
            .I(N__91857));
    LocalMux I__21901 (
            .O(N__91857),
            .I(N__91854));
    Span4Mux_v I__21900 (
            .O(N__91854),
            .I(N__91851));
    Odrv4 I__21899 (
            .O(N__91851),
            .I(\c0.n3_adj_4590 ));
    SRMux I__21898 (
            .O(N__91848),
            .I(N__91845));
    LocalMux I__21897 (
            .O(N__91845),
            .I(\c0.n3_adj_4588 ));
    CascadeMux I__21896 (
            .O(N__91842),
            .I(N__91838));
    InMux I__21895 (
            .O(N__91841),
            .I(N__91835));
    InMux I__21894 (
            .O(N__91838),
            .I(N__91832));
    LocalMux I__21893 (
            .O(N__91835),
            .I(N__91829));
    LocalMux I__21892 (
            .O(N__91832),
            .I(N__91826));
    Span4Mux_h I__21891 (
            .O(N__91829),
            .I(N__91823));
    Span4Mux_v I__21890 (
            .O(N__91826),
            .I(N__91819));
    Span4Mux_v I__21889 (
            .O(N__91823),
            .I(N__91816));
    InMux I__21888 (
            .O(N__91822),
            .I(N__91813));
    Span4Mux_v I__21887 (
            .O(N__91819),
            .I(N__91810));
    Odrv4 I__21886 (
            .O(N__91816),
            .I(\c0.FRAME_MATCHER_i_10 ));
    LocalMux I__21885 (
            .O(N__91813),
            .I(\c0.FRAME_MATCHER_i_10 ));
    Odrv4 I__21884 (
            .O(N__91810),
            .I(\c0.FRAME_MATCHER_i_10 ));
    InMux I__21883 (
            .O(N__91803),
            .I(bfn_24_11_0_));
    SRMux I__21882 (
            .O(N__91800),
            .I(N__91797));
    LocalMux I__21881 (
            .O(N__91797),
            .I(N__91794));
    Span4Mux_v I__21880 (
            .O(N__91794),
            .I(N__91791));
    Span4Mux_v I__21879 (
            .O(N__91791),
            .I(N__91788));
    Odrv4 I__21878 (
            .O(N__91788),
            .I(\c0.n3_adj_4589 ));
    InMux I__21877 (
            .O(N__91785),
            .I(N__91779));
    InMux I__21876 (
            .O(N__91784),
            .I(N__91779));
    LocalMux I__21875 (
            .O(N__91779),
            .I(N__91775));
    InMux I__21874 (
            .O(N__91778),
            .I(N__91772));
    Span12Mux_h I__21873 (
            .O(N__91775),
            .I(N__91769));
    LocalMux I__21872 (
            .O(N__91772),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv12 I__21871 (
            .O(N__91769),
            .I(\c0.FRAME_MATCHER_i_8 ));
    InMux I__21870 (
            .O(N__91764),
            .I(bfn_24_9_0_));
    SRMux I__21869 (
            .O(N__91761),
            .I(N__91758));
    LocalMux I__21868 (
            .O(N__91758),
            .I(N__91755));
    Span4Mux_h I__21867 (
            .O(N__91755),
            .I(N__91752));
    Span4Mux_v I__21866 (
            .O(N__91752),
            .I(N__91749));
    Odrv4 I__21865 (
            .O(N__91749),
            .I(\c0.n3_adj_4587 ));
    InMux I__21864 (
            .O(N__91746),
            .I(N__91743));
    LocalMux I__21863 (
            .O(N__91743),
            .I(N__91740));
    Span4Mux_h I__21862 (
            .O(N__91740),
            .I(N__91737));
    Span4Mux_v I__21861 (
            .O(N__91737),
            .I(N__91732));
    InMux I__21860 (
            .O(N__91736),
            .I(N__91729));
    InMux I__21859 (
            .O(N__91735),
            .I(N__91726));
    Span4Mux_v I__21858 (
            .O(N__91732),
            .I(N__91723));
    LocalMux I__21857 (
            .O(N__91729),
            .I(\c0.FRAME_MATCHER_i_9 ));
    LocalMux I__21856 (
            .O(N__91726),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv4 I__21855 (
            .O(N__91723),
            .I(\c0.FRAME_MATCHER_i_9 ));
    InMux I__21854 (
            .O(N__91716),
            .I(bfn_24_10_0_));
    InMux I__21853 (
            .O(N__91713),
            .I(N__91710));
    LocalMux I__21852 (
            .O(N__91710),
            .I(N__91706));
    InMux I__21851 (
            .O(N__91709),
            .I(N__91703));
    Sp12to4 I__21850 (
            .O(N__91706),
            .I(N__91700));
    LocalMux I__21849 (
            .O(N__91703),
            .I(N__91697));
    Span12Mux_v I__21848 (
            .O(N__91700),
            .I(N__91694));
    Sp12to4 I__21847 (
            .O(N__91697),
            .I(N__91690));
    Span12Mux_h I__21846 (
            .O(N__91694),
            .I(N__91687));
    InMux I__21845 (
            .O(N__91693),
            .I(N__91684));
    Span12Mux_v I__21844 (
            .O(N__91690),
            .I(N__91681));
    Odrv12 I__21843 (
            .O(N__91687),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__21842 (
            .O(N__91684),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv12 I__21841 (
            .O(N__91681),
            .I(\c0.FRAME_MATCHER_i_7 ));
    InMux I__21840 (
            .O(N__91674),
            .I(bfn_24_8_0_));
    SRMux I__21839 (
            .O(N__91671),
            .I(N__91668));
    LocalMux I__21838 (
            .O(N__91668),
            .I(N__91665));
    Sp12to4 I__21837 (
            .O(N__91665),
            .I(N__91662));
    Span12Mux_h I__21836 (
            .O(N__91662),
            .I(N__91659));
    Span12Mux_h I__21835 (
            .O(N__91659),
            .I(N__91656));
    Odrv12 I__21834 (
            .O(N__91656),
            .I(\c0.n3_adj_4586 ));
    InMux I__21833 (
            .O(N__91653),
            .I(N__91650));
    LocalMux I__21832 (
            .O(N__91650),
            .I(N__91645));
    InMux I__21831 (
            .O(N__91649),
            .I(N__91640));
    InMux I__21830 (
            .O(N__91648),
            .I(N__91640));
    Span4Mux_h I__21829 (
            .O(N__91645),
            .I(N__91635));
    LocalMux I__21828 (
            .O(N__91640),
            .I(N__91632));
    CascadeMux I__21827 (
            .O(N__91639),
            .I(N__91629));
    InMux I__21826 (
            .O(N__91638),
            .I(N__91625));
    Span4Mux_h I__21825 (
            .O(N__91635),
            .I(N__91622));
    Span4Mux_h I__21824 (
            .O(N__91632),
            .I(N__91619));
    InMux I__21823 (
            .O(N__91629),
            .I(N__91616));
    InMux I__21822 (
            .O(N__91628),
            .I(N__91613));
    LocalMux I__21821 (
            .O(N__91625),
            .I(N__91610));
    Span4Mux_h I__21820 (
            .O(N__91622),
            .I(N__91607));
    Span4Mux_h I__21819 (
            .O(N__91619),
            .I(N__91602));
    LocalMux I__21818 (
            .O(N__91616),
            .I(N__91602));
    LocalMux I__21817 (
            .O(N__91613),
            .I(N__91599));
    Sp12to4 I__21816 (
            .O(N__91610),
            .I(N__91592));
    Sp12to4 I__21815 (
            .O(N__91607),
            .I(N__91592));
    Sp12to4 I__21814 (
            .O(N__91602),
            .I(N__91592));
    Span12Mux_h I__21813 (
            .O(N__91599),
            .I(N__91586));
    Span12Mux_v I__21812 (
            .O(N__91592),
            .I(N__91586));
    InMux I__21811 (
            .O(N__91591),
            .I(N__91583));
    Odrv12 I__21810 (
            .O(N__91586),
            .I(\c0.FRAME_MATCHER_i_6 ));
    LocalMux I__21809 (
            .O(N__91583),
            .I(\c0.FRAME_MATCHER_i_6 ));
    InMux I__21808 (
            .O(N__91578),
            .I(bfn_24_7_0_));
    SRMux I__21807 (
            .O(N__91575),
            .I(N__91572));
    LocalMux I__21806 (
            .O(N__91572),
            .I(N__91569));
    Span4Mux_v I__21805 (
            .O(N__91569),
            .I(N__91566));
    Span4Mux_v I__21804 (
            .O(N__91566),
            .I(N__91563));
    Odrv4 I__21803 (
            .O(N__91563),
            .I(\c0.n3_adj_4585 ));
    InMux I__21802 (
            .O(N__91560),
            .I(N__91557));
    LocalMux I__21801 (
            .O(N__91557),
            .I(N__91551));
    InMux I__21800 (
            .O(N__91556),
            .I(N__91546));
    InMux I__21799 (
            .O(N__91555),
            .I(N__91546));
    InMux I__21798 (
            .O(N__91554),
            .I(N__91543));
    Span4Mux_v I__21797 (
            .O(N__91551),
            .I(N__91540));
    LocalMux I__21796 (
            .O(N__91546),
            .I(N__91537));
    LocalMux I__21795 (
            .O(N__91543),
            .I(N__91534));
    Span4Mux_h I__21794 (
            .O(N__91540),
            .I(N__91529));
    Span4Mux_v I__21793 (
            .O(N__91537),
            .I(N__91529));
    Span4Mux_v I__21792 (
            .O(N__91534),
            .I(N__91523));
    Span4Mux_v I__21791 (
            .O(N__91529),
            .I(N__91523));
    InMux I__21790 (
            .O(N__91528),
            .I(N__91520));
    Span4Mux_h I__21789 (
            .O(N__91523),
            .I(N__91514));
    LocalMux I__21788 (
            .O(N__91520),
            .I(N__91514));
    InMux I__21787 (
            .O(N__91519),
            .I(N__91511));
    Span4Mux_v I__21786 (
            .O(N__91514),
            .I(N__91508));
    LocalMux I__21785 (
            .O(N__91511),
            .I(N__91505));
    Span4Mux_v I__21784 (
            .O(N__91508),
            .I(N__91502));
    Span4Mux_h I__21783 (
            .O(N__91505),
            .I(N__91498));
    Span4Mux_v I__21782 (
            .O(N__91502),
            .I(N__91495));
    InMux I__21781 (
            .O(N__91501),
            .I(N__91492));
    Odrv4 I__21780 (
            .O(N__91498),
            .I(\c0.FRAME_MATCHER_i_5 ));
    Odrv4 I__21779 (
            .O(N__91495),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__21778 (
            .O(N__91492),
            .I(\c0.FRAME_MATCHER_i_5 ));
    InMux I__21777 (
            .O(N__91485),
            .I(bfn_24_6_0_));
    SRMux I__21776 (
            .O(N__91482),
            .I(N__91479));
    LocalMux I__21775 (
            .O(N__91479),
            .I(N__91476));
    Span12Mux_s7_v I__21774 (
            .O(N__91476),
            .I(N__91473));
    Odrv12 I__21773 (
            .O(N__91473),
            .I(\c0.n3_adj_4584 ));
    InMux I__21772 (
            .O(N__91470),
            .I(N__91464));
    InMux I__21771 (
            .O(N__91469),
            .I(N__91457));
    InMux I__21770 (
            .O(N__91468),
            .I(N__91457));
    InMux I__21769 (
            .O(N__91467),
            .I(N__91457));
    LocalMux I__21768 (
            .O(N__91464),
            .I(N__91453));
    LocalMux I__21767 (
            .O(N__91457),
            .I(N__91449));
    InMux I__21766 (
            .O(N__91456),
            .I(N__91446));
    Span4Mux_h I__21765 (
            .O(N__91453),
            .I(N__91443));
    InMux I__21764 (
            .O(N__91452),
            .I(N__91440));
    Span4Mux_h I__21763 (
            .O(N__91449),
            .I(N__91436));
    LocalMux I__21762 (
            .O(N__91446),
            .I(N__91433));
    Span4Mux_v I__21761 (
            .O(N__91443),
            .I(N__91428));
    LocalMux I__21760 (
            .O(N__91440),
            .I(N__91428));
    InMux I__21759 (
            .O(N__91439),
            .I(N__91425));
    Span4Mux_v I__21758 (
            .O(N__91436),
            .I(N__91422));
    Span4Mux_h I__21757 (
            .O(N__91433),
            .I(N__91419));
    Span4Mux_v I__21756 (
            .O(N__91428),
            .I(N__91416));
    LocalMux I__21755 (
            .O(N__91425),
            .I(N__91409));
    Span4Mux_v I__21754 (
            .O(N__91422),
            .I(N__91409));
    Span4Mux_h I__21753 (
            .O(N__91419),
            .I(N__91409));
    Span4Mux_h I__21752 (
            .O(N__91416),
            .I(N__91406));
    Sp12to4 I__21751 (
            .O(N__91409),
            .I(N__91399));
    Sp12to4 I__21750 (
            .O(N__91406),
            .I(N__91399));
    InMux I__21749 (
            .O(N__91405),
            .I(N__91396));
    InMux I__21748 (
            .O(N__91404),
            .I(N__91393));
    Span12Mux_v I__21747 (
            .O(N__91399),
            .I(N__91390));
    LocalMux I__21746 (
            .O(N__91396),
            .I(\c0.FRAME_MATCHER_i_4 ));
    LocalMux I__21745 (
            .O(N__91393),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv12 I__21744 (
            .O(N__91390),
            .I(\c0.FRAME_MATCHER_i_4 ));
    InMux I__21743 (
            .O(N__91383),
            .I(bfn_24_5_0_));
    SRMux I__21742 (
            .O(N__91380),
            .I(N__91377));
    LocalMux I__21741 (
            .O(N__91377),
            .I(N__91374));
    Odrv12 I__21740 (
            .O(N__91374),
            .I(\c0.n3_adj_4583 ));
    CascadeMux I__21739 (
            .O(N__91371),
            .I(N__91368));
    InMux I__21738 (
            .O(N__91368),
            .I(N__91362));
    CascadeMux I__21737 (
            .O(N__91367),
            .I(N__91359));
    CascadeMux I__21736 (
            .O(N__91366),
            .I(N__91356));
    CascadeMux I__21735 (
            .O(N__91365),
            .I(N__91353));
    LocalMux I__21734 (
            .O(N__91362),
            .I(N__91349));
    InMux I__21733 (
            .O(N__91359),
            .I(N__91346));
    InMux I__21732 (
            .O(N__91356),
            .I(N__91339));
    InMux I__21731 (
            .O(N__91353),
            .I(N__91339));
    InMux I__21730 (
            .O(N__91352),
            .I(N__91339));
    Span4Mux_v I__21729 (
            .O(N__91349),
            .I(N__91336));
    LocalMux I__21728 (
            .O(N__91346),
            .I(N__91333));
    LocalMux I__21727 (
            .O(N__91339),
            .I(N__91330));
    Span4Mux_h I__21726 (
            .O(N__91336),
            .I(N__91322));
    Span4Mux_v I__21725 (
            .O(N__91333),
            .I(N__91322));
    Span4Mux_v I__21724 (
            .O(N__91330),
            .I(N__91322));
    CascadeMux I__21723 (
            .O(N__91329),
            .I(N__91318));
    Span4Mux_v I__21722 (
            .O(N__91322),
            .I(N__91315));
    InMux I__21721 (
            .O(N__91321),
            .I(N__91312));
    InMux I__21720 (
            .O(N__91318),
            .I(N__91309));
    Span4Mux_h I__21719 (
            .O(N__91315),
            .I(N__91302));
    LocalMux I__21718 (
            .O(N__91312),
            .I(N__91302));
    LocalMux I__21717 (
            .O(N__91309),
            .I(N__91302));
    Span4Mux_v I__21716 (
            .O(N__91302),
            .I(N__91299));
    Sp12to4 I__21715 (
            .O(N__91299),
            .I(N__91295));
    InMux I__21714 (
            .O(N__91298),
            .I(N__91291));
    Span12Mux_h I__21713 (
            .O(N__91295),
            .I(N__91288));
    InMux I__21712 (
            .O(N__91294),
            .I(N__91285));
    LocalMux I__21711 (
            .O(N__91291),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv12 I__21710 (
            .O(N__91288),
            .I(\c0.FRAME_MATCHER_i_3 ));
    LocalMux I__21709 (
            .O(N__91285),
            .I(\c0.FRAME_MATCHER_i_3 ));
    InMux I__21708 (
            .O(N__91278),
            .I(bfn_24_4_0_));
    SRMux I__21707 (
            .O(N__91275),
            .I(N__91272));
    LocalMux I__21706 (
            .O(N__91272),
            .I(N__91269));
    Span4Mux_h I__21705 (
            .O(N__91269),
            .I(N__91266));
    Odrv4 I__21704 (
            .O(N__91266),
            .I(\c0.n3_adj_4581 ));
    InMux I__21703 (
            .O(N__91263),
            .I(N__91260));
    LocalMux I__21702 (
            .O(N__91260),
            .I(N__91255));
    InMux I__21701 (
            .O(N__91259),
            .I(N__91252));
    CascadeMux I__21700 (
            .O(N__91258),
            .I(N__91247));
    Span4Mux_h I__21699 (
            .O(N__91255),
            .I(N__91241));
    LocalMux I__21698 (
            .O(N__91252),
            .I(N__91241));
    InMux I__21697 (
            .O(N__91251),
            .I(N__91236));
    InMux I__21696 (
            .O(N__91250),
            .I(N__91231));
    InMux I__21695 (
            .O(N__91247),
            .I(N__91231));
    InMux I__21694 (
            .O(N__91246),
            .I(N__91228));
    Span4Mux_v I__21693 (
            .O(N__91241),
            .I(N__91225));
    InMux I__21692 (
            .O(N__91240),
            .I(N__91222));
    InMux I__21691 (
            .O(N__91239),
            .I(N__91218));
    LocalMux I__21690 (
            .O(N__91236),
            .I(N__91215));
    LocalMux I__21689 (
            .O(N__91231),
            .I(N__91210));
    LocalMux I__21688 (
            .O(N__91228),
            .I(N__91210));
    Span4Mux_v I__21687 (
            .O(N__91225),
            .I(N__91206));
    LocalMux I__21686 (
            .O(N__91222),
            .I(N__91203));
    InMux I__21685 (
            .O(N__91221),
            .I(N__91199));
    LocalMux I__21684 (
            .O(N__91218),
            .I(N__91192));
    Span4Mux_h I__21683 (
            .O(N__91215),
            .I(N__91192));
    Span4Mux_h I__21682 (
            .O(N__91210),
            .I(N__91192));
    InMux I__21681 (
            .O(N__91209),
            .I(N__91189));
    Span4Mux_h I__21680 (
            .O(N__91206),
            .I(N__91184));
    Span4Mux_h I__21679 (
            .O(N__91203),
            .I(N__91184));
    InMux I__21678 (
            .O(N__91202),
            .I(N__91181));
    LocalMux I__21677 (
            .O(N__91199),
            .I(N__91178));
    Span4Mux_v I__21676 (
            .O(N__91192),
            .I(N__91175));
    LocalMux I__21675 (
            .O(N__91189),
            .I(N__91172));
    Sp12to4 I__21674 (
            .O(N__91184),
            .I(N__91169));
    LocalMux I__21673 (
            .O(N__91181),
            .I(N__91166));
    Sp12to4 I__21672 (
            .O(N__91178),
            .I(N__91159));
    Sp12to4 I__21671 (
            .O(N__91175),
            .I(N__91159));
    Span12Mux_h I__21670 (
            .O(N__91172),
            .I(N__91159));
    Span12Mux_v I__21669 (
            .O(N__91169),
            .I(N__91156));
    Sp12to4 I__21668 (
            .O(N__91166),
            .I(N__91150));
    Span12Mux_v I__21667 (
            .O(N__91159),
            .I(N__91150));
    Span12Mux_h I__21666 (
            .O(N__91156),
            .I(N__91147));
    InMux I__21665 (
            .O(N__91155),
            .I(N__91144));
    Odrv12 I__21664 (
            .O(N__91150),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv12 I__21663 (
            .O(N__91147),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__21662 (
            .O(N__91144),
            .I(\c0.FRAME_MATCHER_i_2 ));
    InMux I__21661 (
            .O(N__91137),
            .I(bfn_24_3_0_));
    SRMux I__21660 (
            .O(N__91134),
            .I(N__91131));
    LocalMux I__21659 (
            .O(N__91131),
            .I(N__91128));
    Sp12to4 I__21658 (
            .O(N__91128),
            .I(N__91125));
    Span12Mux_s10_v I__21657 (
            .O(N__91125),
            .I(N__91122));
    Span12Mux_v I__21656 (
            .O(N__91122),
            .I(N__91119));
    Odrv12 I__21655 (
            .O(N__91119),
            .I(\c0.n3_adj_4580 ));
    CascadeMux I__21654 (
            .O(N__91116),
            .I(N__91112));
    InMux I__21653 (
            .O(N__91115),
            .I(N__91107));
    InMux I__21652 (
            .O(N__91112),
            .I(N__91104));
    InMux I__21651 (
            .O(N__91111),
            .I(N__91098));
    InMux I__21650 (
            .O(N__91110),
            .I(N__91094));
    LocalMux I__21649 (
            .O(N__91107),
            .I(N__91089));
    LocalMux I__21648 (
            .O(N__91104),
            .I(N__91089));
    InMux I__21647 (
            .O(N__91103),
            .I(N__91082));
    InMux I__21646 (
            .O(N__91102),
            .I(N__91082));
    InMux I__21645 (
            .O(N__91101),
            .I(N__91082));
    LocalMux I__21644 (
            .O(N__91098),
            .I(N__91079));
    InMux I__21643 (
            .O(N__91097),
            .I(N__91075));
    LocalMux I__21642 (
            .O(N__91094),
            .I(N__91072));
    Span4Mux_v I__21641 (
            .O(N__91089),
            .I(N__91066));
    LocalMux I__21640 (
            .O(N__91082),
            .I(N__91066));
    Span4Mux_v I__21639 (
            .O(N__91079),
            .I(N__91063));
    InMux I__21638 (
            .O(N__91078),
            .I(N__91060));
    LocalMux I__21637 (
            .O(N__91075),
            .I(N__91057));
    Span4Mux_v I__21636 (
            .O(N__91072),
            .I(N__91054));
    InMux I__21635 (
            .O(N__91071),
            .I(N__91051));
    Span4Mux_v I__21634 (
            .O(N__91066),
            .I(N__91048));
    Span4Mux_v I__21633 (
            .O(N__91063),
            .I(N__91045));
    LocalMux I__21632 (
            .O(N__91060),
            .I(N__91042));
    Span4Mux_v I__21631 (
            .O(N__91057),
            .I(N__91039));
    Span4Mux_h I__21630 (
            .O(N__91054),
            .I(N__91036));
    LocalMux I__21629 (
            .O(N__91051),
            .I(N__91033));
    Sp12to4 I__21628 (
            .O(N__91048),
            .I(N__91029));
    Span4Mux_h I__21627 (
            .O(N__91045),
            .I(N__91026));
    Span4Mux_v I__21626 (
            .O(N__91042),
            .I(N__91023));
    Span4Mux_h I__21625 (
            .O(N__91039),
            .I(N__91018));
    Span4Mux_v I__21624 (
            .O(N__91036),
            .I(N__91018));
    Span4Mux_v I__21623 (
            .O(N__91033),
            .I(N__91015));
    InMux I__21622 (
            .O(N__91032),
            .I(N__91012));
    Span12Mux_h I__21621 (
            .O(N__91029),
            .I(N__91009));
    Sp12to4 I__21620 (
            .O(N__91026),
            .I(N__91006));
    Span4Mux_h I__21619 (
            .O(N__91023),
            .I(N__91003));
    Span4Mux_v I__21618 (
            .O(N__91018),
            .I(N__91000));
    Sp12to4 I__21617 (
            .O(N__91015),
            .I(N__90997));
    LocalMux I__21616 (
            .O(N__91012),
            .I(N__90994));
    Span12Mux_v I__21615 (
            .O(N__91009),
            .I(N__90991));
    Span12Mux_h I__21614 (
            .O(N__91006),
            .I(N__90982));
    Sp12to4 I__21613 (
            .O(N__91003),
            .I(N__90982));
    Sp12to4 I__21612 (
            .O(N__91000),
            .I(N__90982));
    Span12Mux_h I__21611 (
            .O(N__90997),
            .I(N__90982));
    Span4Mux_v I__21610 (
            .O(N__90994),
            .I(N__90978));
    Span12Mux_v I__21609 (
            .O(N__90991),
            .I(N__90973));
    Span12Mux_v I__21608 (
            .O(N__90982),
            .I(N__90973));
    InMux I__21607 (
            .O(N__90981),
            .I(N__90970));
    Odrv4 I__21606 (
            .O(N__90978),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv12 I__21605 (
            .O(N__90973),
            .I(\c0.FRAME_MATCHER_i_1 ));
    LocalMux I__21604 (
            .O(N__90970),
            .I(\c0.FRAME_MATCHER_i_1 ));
    InMux I__21603 (
            .O(N__90963),
            .I(bfn_24_2_0_));
    SRMux I__21602 (
            .O(N__90960),
            .I(N__90957));
    LocalMux I__21601 (
            .O(N__90957),
            .I(N__90954));
    Sp12to4 I__21600 (
            .O(N__90954),
            .I(N__90951));
    Span12Mux_s11_h I__21599 (
            .O(N__90951),
            .I(N__90948));
    Span12Mux_v I__21598 (
            .O(N__90948),
            .I(N__90945));
    Odrv12 I__21597 (
            .O(N__90945),
            .I(\c0.n3_adj_4579 ));
    InMux I__21596 (
            .O(N__90942),
            .I(N__90937));
    InMux I__21595 (
            .O(N__90941),
            .I(N__90934));
    InMux I__21594 (
            .O(N__90940),
            .I(N__90931));
    LocalMux I__21593 (
            .O(N__90937),
            .I(N__90922));
    LocalMux I__21592 (
            .O(N__90934),
            .I(N__90922));
    LocalMux I__21591 (
            .O(N__90931),
            .I(N__90922));
    InMux I__21590 (
            .O(N__90930),
            .I(N__90917));
    InMux I__21589 (
            .O(N__90929),
            .I(N__90917));
    Odrv4 I__21588 (
            .O(N__90922),
            .I(\c0.n18469 ));
    LocalMux I__21587 (
            .O(N__90917),
            .I(\c0.n18469 ));
    CascadeMux I__21586 (
            .O(N__90912),
            .I(N__90909));
    InMux I__21585 (
            .O(N__90909),
            .I(N__90906));
    LocalMux I__21584 (
            .O(N__90906),
            .I(N__90903));
    Span4Mux_s0_v I__21583 (
            .O(N__90903),
            .I(N__90900));
    Span4Mux_h I__21582 (
            .O(N__90900),
            .I(N__90897));
    Sp12to4 I__21581 (
            .O(N__90897),
            .I(N__90894));
    Span12Mux_s5_v I__21580 (
            .O(N__90894),
            .I(N__90891));
    Span12Mux_v I__21579 (
            .O(N__90891),
            .I(N__90888));
    Odrv12 I__21578 (
            .O(N__90888),
            .I(\c0.n161 ));
    CascadeMux I__21577 (
            .O(N__90885),
            .I(N__90881));
    InMux I__21576 (
            .O(N__90884),
            .I(N__90878));
    InMux I__21575 (
            .O(N__90881),
            .I(N__90874));
    LocalMux I__21574 (
            .O(N__90878),
            .I(N__90867));
    InMux I__21573 (
            .O(N__90877),
            .I(N__90864));
    LocalMux I__21572 (
            .O(N__90874),
            .I(N__90861));
    InMux I__21571 (
            .O(N__90873),
            .I(N__90858));
    InMux I__21570 (
            .O(N__90872),
            .I(N__90855));
    CascadeMux I__21569 (
            .O(N__90871),
            .I(N__90852));
    InMux I__21568 (
            .O(N__90870),
            .I(N__90849));
    Span4Mux_v I__21567 (
            .O(N__90867),
            .I(N__90846));
    LocalMux I__21566 (
            .O(N__90864),
            .I(N__90843));
    Span4Mux_v I__21565 (
            .O(N__90861),
            .I(N__90840));
    LocalMux I__21564 (
            .O(N__90858),
            .I(N__90835));
    LocalMux I__21563 (
            .O(N__90855),
            .I(N__90835));
    InMux I__21562 (
            .O(N__90852),
            .I(N__90832));
    LocalMux I__21561 (
            .O(N__90849),
            .I(N__90829));
    Span4Mux_h I__21560 (
            .O(N__90846),
            .I(N__90826));
    Span4Mux_v I__21559 (
            .O(N__90843),
            .I(N__90819));
    Span4Mux_h I__21558 (
            .O(N__90840),
            .I(N__90819));
    Span4Mux_v I__21557 (
            .O(N__90835),
            .I(N__90819));
    LocalMux I__21556 (
            .O(N__90832),
            .I(N__90814));
    Span4Mux_h I__21555 (
            .O(N__90829),
            .I(N__90814));
    Odrv4 I__21554 (
            .O(N__90826),
            .I(n17453));
    Odrv4 I__21553 (
            .O(N__90819),
            .I(n17453));
    Odrv4 I__21552 (
            .O(N__90814),
            .I(n17453));
    InMux I__21551 (
            .O(N__90807),
            .I(N__90804));
    LocalMux I__21550 (
            .O(N__90804),
            .I(N__90801));
    Odrv4 I__21549 (
            .O(N__90801),
            .I(n36101));
    CascadeMux I__21548 (
            .O(N__90798),
            .I(n26_cascade_));
    InMux I__21547 (
            .O(N__90795),
            .I(N__90790));
    CascadeMux I__21546 (
            .O(N__90794),
            .I(N__90786));
    InMux I__21545 (
            .O(N__90793),
            .I(N__90782));
    LocalMux I__21544 (
            .O(N__90790),
            .I(N__90779));
    InMux I__21543 (
            .O(N__90789),
            .I(N__90775));
    InMux I__21542 (
            .O(N__90786),
            .I(N__90771));
    CascadeMux I__21541 (
            .O(N__90785),
            .I(N__90768));
    LocalMux I__21540 (
            .O(N__90782),
            .I(N__90764));
    Span4Mux_v I__21539 (
            .O(N__90779),
            .I(N__90761));
    InMux I__21538 (
            .O(N__90778),
            .I(N__90755));
    LocalMux I__21537 (
            .O(N__90775),
            .I(N__90752));
    InMux I__21536 (
            .O(N__90774),
            .I(N__90749));
    LocalMux I__21535 (
            .O(N__90771),
            .I(N__90746));
    InMux I__21534 (
            .O(N__90768),
            .I(N__90743));
    InMux I__21533 (
            .O(N__90767),
            .I(N__90740));
    Span4Mux_h I__21532 (
            .O(N__90764),
            .I(N__90735));
    Span4Mux_v I__21531 (
            .O(N__90761),
            .I(N__90735));
    InMux I__21530 (
            .O(N__90760),
            .I(N__90732));
    InMux I__21529 (
            .O(N__90759),
            .I(N__90729));
    InMux I__21528 (
            .O(N__90758),
            .I(N__90725));
    LocalMux I__21527 (
            .O(N__90755),
            .I(N__90721));
    Span4Mux_v I__21526 (
            .O(N__90752),
            .I(N__90718));
    LocalMux I__21525 (
            .O(N__90749),
            .I(N__90711));
    Span4Mux_h I__21524 (
            .O(N__90746),
            .I(N__90711));
    LocalMux I__21523 (
            .O(N__90743),
            .I(N__90711));
    LocalMux I__21522 (
            .O(N__90740),
            .I(N__90702));
    Span4Mux_h I__21521 (
            .O(N__90735),
            .I(N__90702));
    LocalMux I__21520 (
            .O(N__90732),
            .I(N__90702));
    LocalMux I__21519 (
            .O(N__90729),
            .I(N__90702));
    InMux I__21518 (
            .O(N__90728),
            .I(N__90699));
    LocalMux I__21517 (
            .O(N__90725),
            .I(N__90696));
    InMux I__21516 (
            .O(N__90724),
            .I(N__90689));
    Span4Mux_v I__21515 (
            .O(N__90721),
            .I(N__90686));
    Span4Mux_v I__21514 (
            .O(N__90718),
            .I(N__90683));
    Span4Mux_v I__21513 (
            .O(N__90711),
            .I(N__90678));
    Span4Mux_v I__21512 (
            .O(N__90702),
            .I(N__90678));
    LocalMux I__21511 (
            .O(N__90699),
            .I(N__90675));
    Span4Mux_v I__21510 (
            .O(N__90696),
            .I(N__90672));
    InMux I__21509 (
            .O(N__90695),
            .I(N__90669));
    InMux I__21508 (
            .O(N__90694),
            .I(N__90666));
    InMux I__21507 (
            .O(N__90693),
            .I(N__90663));
    InMux I__21506 (
            .O(N__90692),
            .I(N__90660));
    LocalMux I__21505 (
            .O(N__90689),
            .I(N__90657));
    Sp12to4 I__21504 (
            .O(N__90686),
            .I(N__90650));
    Sp12to4 I__21503 (
            .O(N__90683),
            .I(N__90650));
    Sp12to4 I__21502 (
            .O(N__90678),
            .I(N__90650));
    Span4Mux_v I__21501 (
            .O(N__90675),
            .I(N__90643));
    Span4Mux_h I__21500 (
            .O(N__90672),
            .I(N__90643));
    LocalMux I__21499 (
            .O(N__90669),
            .I(N__90643));
    LocalMux I__21498 (
            .O(N__90666),
            .I(byte_transmit_counter_4));
    LocalMux I__21497 (
            .O(N__90663),
            .I(byte_transmit_counter_4));
    LocalMux I__21496 (
            .O(N__90660),
            .I(byte_transmit_counter_4));
    Odrv4 I__21495 (
            .O(N__90657),
            .I(byte_transmit_counter_4));
    Odrv12 I__21494 (
            .O(N__90650),
            .I(byte_transmit_counter_4));
    Odrv4 I__21493 (
            .O(N__90643),
            .I(byte_transmit_counter_4));
    InMux I__21492 (
            .O(N__90630),
            .I(N__90627));
    LocalMux I__21491 (
            .O(N__90627),
            .I(N__90624));
    Span4Mux_v I__21490 (
            .O(N__90624),
            .I(N__90621));
    Sp12to4 I__21489 (
            .O(N__90621),
            .I(N__90618));
    Span12Mux_s5_h I__21488 (
            .O(N__90618),
            .I(N__90615));
    Span12Mux_h I__21487 (
            .O(N__90615),
            .I(N__90612));
    Odrv12 I__21486 (
            .O(N__90612),
            .I(n36102));
    InMux I__21485 (
            .O(N__90609),
            .I(N__90606));
    LocalMux I__21484 (
            .O(N__90606),
            .I(N__90603));
    Span4Mux_v I__21483 (
            .O(N__90603),
            .I(N__90599));
    InMux I__21482 (
            .O(N__90602),
            .I(N__90596));
    Odrv4 I__21481 (
            .O(N__90599),
            .I(\c0.n17570 ));
    LocalMux I__21480 (
            .O(N__90596),
            .I(\c0.n17570 ));
    CascadeMux I__21479 (
            .O(N__90591),
            .I(\c0.n14_adj_4522_cascade_ ));
    CascadeMux I__21478 (
            .O(N__90588),
            .I(\c0.n9_adj_4524_cascade_ ));
    InMux I__21477 (
            .O(N__90585),
            .I(N__90582));
    LocalMux I__21476 (
            .O(N__90582),
            .I(\c0.data_out_frame_29_4 ));
    InMux I__21475 (
            .O(N__90579),
            .I(N__90575));
    InMux I__21474 (
            .O(N__90578),
            .I(N__90570));
    LocalMux I__21473 (
            .O(N__90575),
            .I(N__90567));
    InMux I__21472 (
            .O(N__90574),
            .I(N__90562));
    InMux I__21471 (
            .O(N__90573),
            .I(N__90562));
    LocalMux I__21470 (
            .O(N__90570),
            .I(N__90559));
    Span4Mux_v I__21469 (
            .O(N__90567),
            .I(N__90554));
    LocalMux I__21468 (
            .O(N__90562),
            .I(N__90554));
    Span4Mux_v I__21467 (
            .O(N__90559),
            .I(N__90551));
    Span4Mux_h I__21466 (
            .O(N__90554),
            .I(N__90548));
    Odrv4 I__21465 (
            .O(N__90551),
            .I(\c0.n33795 ));
    Odrv4 I__21464 (
            .O(N__90548),
            .I(\c0.n33795 ));
    InMux I__21463 (
            .O(N__90543),
            .I(N__90540));
    LocalMux I__21462 (
            .O(N__90540),
            .I(N__90537));
    Odrv4 I__21461 (
            .O(N__90537),
            .I(\c0.n42_adj_4640 ));
    CascadeMux I__21460 (
            .O(N__90534),
            .I(\c0.n41_adj_4642_cascade_ ));
    InMux I__21459 (
            .O(N__90531),
            .I(N__90528));
    LocalMux I__21458 (
            .O(N__90528),
            .I(\c0.n43_adj_4641 ));
    InMux I__21457 (
            .O(N__90525),
            .I(N__90522));
    LocalMux I__21456 (
            .O(N__90522),
            .I(\c0.n40_adj_4643 ));
    InMux I__21455 (
            .O(N__90519),
            .I(N__90516));
    LocalMux I__21454 (
            .O(N__90516),
            .I(N__90513));
    Odrv4 I__21453 (
            .O(N__90513),
            .I(\c0.n39_adj_4644 ));
    CascadeMux I__21452 (
            .O(N__90510),
            .I(\c0.n50_cascade_ ));
    InMux I__21451 (
            .O(N__90507),
            .I(N__90504));
    LocalMux I__21450 (
            .O(N__90504),
            .I(N__90501));
    Odrv4 I__21449 (
            .O(N__90501),
            .I(\c0.n45_adj_4645 ));
    InMux I__21448 (
            .O(N__90498),
            .I(N__90494));
    CascadeMux I__21447 (
            .O(N__90497),
            .I(N__90490));
    LocalMux I__21446 (
            .O(N__90494),
            .I(N__90487));
    InMux I__21445 (
            .O(N__90493),
            .I(N__90484));
    InMux I__21444 (
            .O(N__90490),
            .I(N__90481));
    Span4Mux_h I__21443 (
            .O(N__90487),
            .I(N__90476));
    LocalMux I__21442 (
            .O(N__90484),
            .I(N__90476));
    LocalMux I__21441 (
            .O(N__90481),
            .I(N__90473));
    Span4Mux_v I__21440 (
            .O(N__90476),
            .I(N__90470));
    Span4Mux_h I__21439 (
            .O(N__90473),
            .I(N__90467));
    Sp12to4 I__21438 (
            .O(N__90470),
            .I(N__90464));
    Span4Mux_h I__21437 (
            .O(N__90467),
            .I(N__90461));
    Span12Mux_h I__21436 (
            .O(N__90464),
            .I(N__90458));
    Odrv4 I__21435 (
            .O(N__90461),
            .I(\c0.n18083 ));
    Odrv12 I__21434 (
            .O(N__90458),
            .I(\c0.n18083 ));
    CascadeMux I__21433 (
            .O(N__90453),
            .I(N__90450));
    InMux I__21432 (
            .O(N__90450),
            .I(N__90445));
    InMux I__21431 (
            .O(N__90449),
            .I(N__90442));
    InMux I__21430 (
            .O(N__90448),
            .I(N__90439));
    LocalMux I__21429 (
            .O(N__90445),
            .I(N__90434));
    LocalMux I__21428 (
            .O(N__90442),
            .I(N__90434));
    LocalMux I__21427 (
            .O(N__90439),
            .I(\c0.n17669 ));
    Odrv12 I__21426 (
            .O(N__90434),
            .I(\c0.n17669 ));
    InMux I__21425 (
            .O(N__90429),
            .I(N__90426));
    LocalMux I__21424 (
            .O(N__90426),
            .I(\c0.n31299 ));
    CascadeMux I__21423 (
            .O(N__90423),
            .I(\c0.n31299_cascade_ ));
    InMux I__21422 (
            .O(N__90420),
            .I(N__90417));
    LocalMux I__21421 (
            .O(N__90417),
            .I(N__90414));
    Span4Mux_h I__21420 (
            .O(N__90414),
            .I(N__90411));
    Odrv4 I__21419 (
            .O(N__90411),
            .I(\c0.data_out_frame_28_6 ));
    InMux I__21418 (
            .O(N__90408),
            .I(N__90405));
    LocalMux I__21417 (
            .O(N__90405),
            .I(N__90402));
    Odrv4 I__21416 (
            .O(N__90402),
            .I(\c0.n32238 ));
    CascadeMux I__21415 (
            .O(N__90399),
            .I(\c0.n32238_cascade_ ));
    InMux I__21414 (
            .O(N__90396),
            .I(N__90388));
    CascadeMux I__21413 (
            .O(N__90395),
            .I(N__90382));
    CascadeMux I__21412 (
            .O(N__90394),
            .I(N__90367));
    CascadeMux I__21411 (
            .O(N__90393),
            .I(N__90364));
    InMux I__21410 (
            .O(N__90392),
            .I(N__90361));
    CascadeMux I__21409 (
            .O(N__90391),
            .I(N__90358));
    LocalMux I__21408 (
            .O(N__90388),
            .I(N__90355));
    InMux I__21407 (
            .O(N__90387),
            .I(N__90348));
    InMux I__21406 (
            .O(N__90386),
            .I(N__90348));
    InMux I__21405 (
            .O(N__90385),
            .I(N__90348));
    InMux I__21404 (
            .O(N__90382),
            .I(N__90345));
    InMux I__21403 (
            .O(N__90381),
            .I(N__90340));
    CascadeMux I__21402 (
            .O(N__90380),
            .I(N__90336));
    CascadeMux I__21401 (
            .O(N__90379),
            .I(N__90332));
    CascadeMux I__21400 (
            .O(N__90378),
            .I(N__90329));
    CascadeMux I__21399 (
            .O(N__90377),
            .I(N__90326));
    InMux I__21398 (
            .O(N__90376),
            .I(N__90323));
    CascadeMux I__21397 (
            .O(N__90375),
            .I(N__90311));
    InMux I__21396 (
            .O(N__90374),
            .I(N__90304));
    InMux I__21395 (
            .O(N__90373),
            .I(N__90304));
    InMux I__21394 (
            .O(N__90372),
            .I(N__90304));
    CascadeMux I__21393 (
            .O(N__90371),
            .I(N__90301));
    InMux I__21392 (
            .O(N__90370),
            .I(N__90298));
    InMux I__21391 (
            .O(N__90367),
            .I(N__90295));
    InMux I__21390 (
            .O(N__90364),
            .I(N__90292));
    LocalMux I__21389 (
            .O(N__90361),
            .I(N__90289));
    InMux I__21388 (
            .O(N__90358),
            .I(N__90286));
    Span4Mux_v I__21387 (
            .O(N__90355),
            .I(N__90279));
    LocalMux I__21386 (
            .O(N__90348),
            .I(N__90279));
    LocalMux I__21385 (
            .O(N__90345),
            .I(N__90279));
    InMux I__21384 (
            .O(N__90344),
            .I(N__90276));
    InMux I__21383 (
            .O(N__90343),
            .I(N__90273));
    LocalMux I__21382 (
            .O(N__90340),
            .I(N__90270));
    InMux I__21381 (
            .O(N__90339),
            .I(N__90267));
    InMux I__21380 (
            .O(N__90336),
            .I(N__90264));
    InMux I__21379 (
            .O(N__90335),
            .I(N__90259));
    InMux I__21378 (
            .O(N__90332),
            .I(N__90259));
    InMux I__21377 (
            .O(N__90329),
            .I(N__90254));
    InMux I__21376 (
            .O(N__90326),
            .I(N__90254));
    LocalMux I__21375 (
            .O(N__90323),
            .I(N__90251));
    InMux I__21374 (
            .O(N__90322),
            .I(N__90244));
    InMux I__21373 (
            .O(N__90321),
            .I(N__90244));
    InMux I__21372 (
            .O(N__90320),
            .I(N__90244));
    InMux I__21371 (
            .O(N__90319),
            .I(N__90239));
    InMux I__21370 (
            .O(N__90318),
            .I(N__90239));
    InMux I__21369 (
            .O(N__90317),
            .I(N__90232));
    InMux I__21368 (
            .O(N__90316),
            .I(N__90232));
    InMux I__21367 (
            .O(N__90315),
            .I(N__90232));
    CascadeMux I__21366 (
            .O(N__90314),
            .I(N__90228));
    InMux I__21365 (
            .O(N__90311),
            .I(N__90225));
    LocalMux I__21364 (
            .O(N__90304),
            .I(N__90222));
    InMux I__21363 (
            .O(N__90301),
            .I(N__90219));
    LocalMux I__21362 (
            .O(N__90298),
            .I(N__90212));
    LocalMux I__21361 (
            .O(N__90295),
            .I(N__90212));
    LocalMux I__21360 (
            .O(N__90292),
            .I(N__90212));
    Span4Mux_v I__21359 (
            .O(N__90289),
            .I(N__90209));
    LocalMux I__21358 (
            .O(N__90286),
            .I(N__90201));
    Span4Mux_v I__21357 (
            .O(N__90279),
            .I(N__90201));
    LocalMux I__21356 (
            .O(N__90276),
            .I(N__90194));
    LocalMux I__21355 (
            .O(N__90273),
            .I(N__90194));
    Span4Mux_v I__21354 (
            .O(N__90270),
            .I(N__90194));
    LocalMux I__21353 (
            .O(N__90267),
            .I(N__90183));
    LocalMux I__21352 (
            .O(N__90264),
            .I(N__90183));
    LocalMux I__21351 (
            .O(N__90259),
            .I(N__90183));
    LocalMux I__21350 (
            .O(N__90254),
            .I(N__90183));
    Span4Mux_v I__21349 (
            .O(N__90251),
            .I(N__90180));
    LocalMux I__21348 (
            .O(N__90244),
            .I(N__90173));
    LocalMux I__21347 (
            .O(N__90239),
            .I(N__90173));
    LocalMux I__21346 (
            .O(N__90232),
            .I(N__90173));
    InMux I__21345 (
            .O(N__90231),
            .I(N__90170));
    InMux I__21344 (
            .O(N__90228),
            .I(N__90167));
    LocalMux I__21343 (
            .O(N__90225),
            .I(N__90156));
    Span4Mux_v I__21342 (
            .O(N__90222),
            .I(N__90156));
    LocalMux I__21341 (
            .O(N__90219),
            .I(N__90156));
    Span4Mux_v I__21340 (
            .O(N__90212),
            .I(N__90156));
    Span4Mux_h I__21339 (
            .O(N__90209),
            .I(N__90156));
    InMux I__21338 (
            .O(N__90208),
            .I(N__90149));
    InMux I__21337 (
            .O(N__90207),
            .I(N__90149));
    InMux I__21336 (
            .O(N__90206),
            .I(N__90149));
    Span4Mux_v I__21335 (
            .O(N__90201),
            .I(N__90144));
    Span4Mux_h I__21334 (
            .O(N__90194),
            .I(N__90144));
    InMux I__21333 (
            .O(N__90193),
            .I(N__90141));
    InMux I__21332 (
            .O(N__90192),
            .I(N__90138));
    Span4Mux_v I__21331 (
            .O(N__90183),
            .I(N__90133));
    Span4Mux_h I__21330 (
            .O(N__90180),
            .I(N__90133));
    Span4Mux_v I__21329 (
            .O(N__90173),
            .I(N__90128));
    LocalMux I__21328 (
            .O(N__90170),
            .I(N__90128));
    LocalMux I__21327 (
            .O(N__90167),
            .I(N__90123));
    Span4Mux_h I__21326 (
            .O(N__90156),
            .I(N__90123));
    LocalMux I__21325 (
            .O(N__90149),
            .I(N__90118));
    Span4Mux_h I__21324 (
            .O(N__90144),
            .I(N__90118));
    LocalMux I__21323 (
            .O(N__90141),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__21322 (
            .O(N__90138),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__21321 (
            .O(N__90133),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__21320 (
            .O(N__90128),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__21319 (
            .O(N__90123),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__21318 (
            .O(N__90118),
            .I(\c0.byte_transmit_counter_1 ));
    InMux I__21317 (
            .O(N__90105),
            .I(N__90097));
    CascadeMux I__21316 (
            .O(N__90104),
            .I(N__90090));
    CascadeMux I__21315 (
            .O(N__90103),
            .I(N__90087));
    InMux I__21314 (
            .O(N__90102),
            .I(N__90079));
    InMux I__21313 (
            .O(N__90101),
            .I(N__90079));
    InMux I__21312 (
            .O(N__90100),
            .I(N__90076));
    LocalMux I__21311 (
            .O(N__90097),
            .I(N__90071));
    InMux I__21310 (
            .O(N__90096),
            .I(N__90068));
    InMux I__21309 (
            .O(N__90095),
            .I(N__90065));
    InMux I__21308 (
            .O(N__90094),
            .I(N__90055));
    InMux I__21307 (
            .O(N__90093),
            .I(N__90055));
    InMux I__21306 (
            .O(N__90090),
            .I(N__90055));
    InMux I__21305 (
            .O(N__90087),
            .I(N__90055));
    InMux I__21304 (
            .O(N__90086),
            .I(N__90052));
    InMux I__21303 (
            .O(N__90085),
            .I(N__90048));
    InMux I__21302 (
            .O(N__90084),
            .I(N__90041));
    LocalMux I__21301 (
            .O(N__90079),
            .I(N__90034));
    LocalMux I__21300 (
            .O(N__90076),
            .I(N__90034));
    InMux I__21299 (
            .O(N__90075),
            .I(N__90031));
    CascadeMux I__21298 (
            .O(N__90074),
            .I(N__90028));
    Span4Mux_h I__21297 (
            .O(N__90071),
            .I(N__90024));
    LocalMux I__21296 (
            .O(N__90068),
            .I(N__90019));
    LocalMux I__21295 (
            .O(N__90065),
            .I(N__90019));
    InMux I__21294 (
            .O(N__90064),
            .I(N__90014));
    LocalMux I__21293 (
            .O(N__90055),
            .I(N__90009));
    LocalMux I__21292 (
            .O(N__90052),
            .I(N__90009));
    InMux I__21291 (
            .O(N__90051),
            .I(N__90006));
    LocalMux I__21290 (
            .O(N__90048),
            .I(N__90001));
    InMux I__21289 (
            .O(N__90047),
            .I(N__89998));
    InMux I__21288 (
            .O(N__90046),
            .I(N__89995));
    InMux I__21287 (
            .O(N__90045),
            .I(N__89992));
    InMux I__21286 (
            .O(N__90044),
            .I(N__89989));
    LocalMux I__21285 (
            .O(N__90041),
            .I(N__89986));
    InMux I__21284 (
            .O(N__90040),
            .I(N__89983));
    InMux I__21283 (
            .O(N__90039),
            .I(N__89980));
    Span4Mux_v I__21282 (
            .O(N__90034),
            .I(N__89975));
    LocalMux I__21281 (
            .O(N__90031),
            .I(N__89975));
    InMux I__21280 (
            .O(N__90028),
            .I(N__89971));
    InMux I__21279 (
            .O(N__90027),
            .I(N__89968));
    Span4Mux_v I__21278 (
            .O(N__90024),
            .I(N__89963));
    Span4Mux_v I__21277 (
            .O(N__90019),
            .I(N__89963));
    InMux I__21276 (
            .O(N__90018),
            .I(N__89960));
    InMux I__21275 (
            .O(N__90017),
            .I(N__89957));
    LocalMux I__21274 (
            .O(N__90014),
            .I(N__89950));
    Span4Mux_v I__21273 (
            .O(N__90009),
            .I(N__89950));
    LocalMux I__21272 (
            .O(N__90006),
            .I(N__89950));
    InMux I__21271 (
            .O(N__90005),
            .I(N__89946));
    InMux I__21270 (
            .O(N__90004),
            .I(N__89943));
    Span4Mux_h I__21269 (
            .O(N__90001),
            .I(N__89936));
    LocalMux I__21268 (
            .O(N__89998),
            .I(N__89936));
    LocalMux I__21267 (
            .O(N__89995),
            .I(N__89936));
    LocalMux I__21266 (
            .O(N__89992),
            .I(N__89933));
    LocalMux I__21265 (
            .O(N__89989),
            .I(N__89928));
    Span4Mux_v I__21264 (
            .O(N__89986),
            .I(N__89928));
    LocalMux I__21263 (
            .O(N__89983),
            .I(N__89921));
    LocalMux I__21262 (
            .O(N__89980),
            .I(N__89921));
    Span4Mux_h I__21261 (
            .O(N__89975),
            .I(N__89921));
    InMux I__21260 (
            .O(N__89974),
            .I(N__89918));
    LocalMux I__21259 (
            .O(N__89971),
            .I(N__89911));
    LocalMux I__21258 (
            .O(N__89968),
            .I(N__89911));
    Span4Mux_h I__21257 (
            .O(N__89963),
            .I(N__89911));
    LocalMux I__21256 (
            .O(N__89960),
            .I(N__89904));
    LocalMux I__21255 (
            .O(N__89957),
            .I(N__89904));
    Span4Mux_h I__21254 (
            .O(N__89950),
            .I(N__89904));
    InMux I__21253 (
            .O(N__89949),
            .I(N__89901));
    LocalMux I__21252 (
            .O(N__89946),
            .I(N__89892));
    LocalMux I__21251 (
            .O(N__89943),
            .I(N__89892));
    Span4Mux_h I__21250 (
            .O(N__89936),
            .I(N__89892));
    Span4Mux_v I__21249 (
            .O(N__89933),
            .I(N__89892));
    Span4Mux_v I__21248 (
            .O(N__89928),
            .I(N__89885));
    Span4Mux_v I__21247 (
            .O(N__89921),
            .I(N__89885));
    LocalMux I__21246 (
            .O(N__89918),
            .I(N__89885));
    Span4Mux_h I__21245 (
            .O(N__89911),
            .I(N__89880));
    Span4Mux_v I__21244 (
            .O(N__89904),
            .I(N__89880));
    LocalMux I__21243 (
            .O(N__89901),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__21242 (
            .O(N__89892),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__21241 (
            .O(N__89885),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__21240 (
            .O(N__89880),
            .I(\c0.byte_transmit_counter_2 ));
    InMux I__21239 (
            .O(N__89871),
            .I(N__89868));
    LocalMux I__21238 (
            .O(N__89868),
            .I(N__89864));
    CascadeMux I__21237 (
            .O(N__89867),
            .I(N__89861));
    Span4Mux_v I__21236 (
            .O(N__89864),
            .I(N__89858));
    InMux I__21235 (
            .O(N__89861),
            .I(N__89855));
    Span4Mux_v I__21234 (
            .O(N__89858),
            .I(N__89852));
    LocalMux I__21233 (
            .O(N__89855),
            .I(data_out_frame_21_0));
    Odrv4 I__21232 (
            .O(N__89852),
            .I(data_out_frame_21_0));
    CascadeMux I__21231 (
            .O(N__89847),
            .I(\c0.n14078_cascade_ ));
    InMux I__21230 (
            .O(N__89844),
            .I(N__89841));
    LocalMux I__21229 (
            .O(N__89841),
            .I(N__89837));
    InMux I__21228 (
            .O(N__89840),
            .I(N__89834));
    Span4Mux_h I__21227 (
            .O(N__89837),
            .I(N__89831));
    LocalMux I__21226 (
            .O(N__89834),
            .I(data_out_frame_17_0));
    Odrv4 I__21225 (
            .O(N__89831),
            .I(data_out_frame_17_0));
    CascadeMux I__21224 (
            .O(N__89826),
            .I(N__89820));
    InMux I__21223 (
            .O(N__89825),
            .I(N__89812));
    InMux I__21222 (
            .O(N__89824),
            .I(N__89812));
    InMux I__21221 (
            .O(N__89823),
            .I(N__89812));
    InMux I__21220 (
            .O(N__89820),
            .I(N__89809));
    CascadeMux I__21219 (
            .O(N__89819),
            .I(N__89804));
    LocalMux I__21218 (
            .O(N__89812),
            .I(N__89799));
    LocalMux I__21217 (
            .O(N__89809),
            .I(N__89799));
    CascadeMux I__21216 (
            .O(N__89808),
            .I(N__89791));
    CascadeMux I__21215 (
            .O(N__89807),
            .I(N__89788));
    InMux I__21214 (
            .O(N__89804),
            .I(N__89785));
    Span4Mux_v I__21213 (
            .O(N__89799),
            .I(N__89781));
    InMux I__21212 (
            .O(N__89798),
            .I(N__89778));
    InMux I__21211 (
            .O(N__89797),
            .I(N__89775));
    InMux I__21210 (
            .O(N__89796),
            .I(N__89768));
    InMux I__21209 (
            .O(N__89795),
            .I(N__89765));
    CascadeMux I__21208 (
            .O(N__89794),
            .I(N__89762));
    InMux I__21207 (
            .O(N__89791),
            .I(N__89753));
    InMux I__21206 (
            .O(N__89788),
            .I(N__89753));
    LocalMux I__21205 (
            .O(N__89785),
            .I(N__89749));
    InMux I__21204 (
            .O(N__89784),
            .I(N__89746));
    Span4Mux_h I__21203 (
            .O(N__89781),
            .I(N__89739));
    LocalMux I__21202 (
            .O(N__89778),
            .I(N__89739));
    LocalMux I__21201 (
            .O(N__89775),
            .I(N__89739));
    InMux I__21200 (
            .O(N__89774),
            .I(N__89736));
    InMux I__21199 (
            .O(N__89773),
            .I(N__89730));
    InMux I__21198 (
            .O(N__89772),
            .I(N__89730));
    InMux I__21197 (
            .O(N__89771),
            .I(N__89727));
    LocalMux I__21196 (
            .O(N__89768),
            .I(N__89724));
    LocalMux I__21195 (
            .O(N__89765),
            .I(N__89721));
    InMux I__21194 (
            .O(N__89762),
            .I(N__89718));
    InMux I__21193 (
            .O(N__89761),
            .I(N__89713));
    InMux I__21192 (
            .O(N__89760),
            .I(N__89713));
    InMux I__21191 (
            .O(N__89759),
            .I(N__89707));
    InMux I__21190 (
            .O(N__89758),
            .I(N__89707));
    LocalMux I__21189 (
            .O(N__89753),
            .I(N__89704));
    InMux I__21188 (
            .O(N__89752),
            .I(N__89701));
    Span4Mux_v I__21187 (
            .O(N__89749),
            .I(N__89696));
    LocalMux I__21186 (
            .O(N__89746),
            .I(N__89696));
    Span4Mux_v I__21185 (
            .O(N__89739),
            .I(N__89693));
    LocalMux I__21184 (
            .O(N__89736),
            .I(N__89690));
    InMux I__21183 (
            .O(N__89735),
            .I(N__89687));
    LocalMux I__21182 (
            .O(N__89730),
            .I(N__89682));
    LocalMux I__21181 (
            .O(N__89727),
            .I(N__89682));
    Span4Mux_h I__21180 (
            .O(N__89724),
            .I(N__89679));
    Span4Mux_h I__21179 (
            .O(N__89721),
            .I(N__89672));
    LocalMux I__21178 (
            .O(N__89718),
            .I(N__89672));
    LocalMux I__21177 (
            .O(N__89713),
            .I(N__89672));
    InMux I__21176 (
            .O(N__89712),
            .I(N__89669));
    LocalMux I__21175 (
            .O(N__89707),
            .I(N__89666));
    Span4Mux_h I__21174 (
            .O(N__89704),
            .I(N__89663));
    LocalMux I__21173 (
            .O(N__89701),
            .I(N__89660));
    Span4Mux_h I__21172 (
            .O(N__89696),
            .I(N__89657));
    Span4Mux_h I__21171 (
            .O(N__89693),
            .I(N__89652));
    Span4Mux_v I__21170 (
            .O(N__89690),
            .I(N__89652));
    LocalMux I__21169 (
            .O(N__89687),
            .I(N__89645));
    Span4Mux_v I__21168 (
            .O(N__89682),
            .I(N__89645));
    Span4Mux_h I__21167 (
            .O(N__89679),
            .I(N__89645));
    Span4Mux_v I__21166 (
            .O(N__89672),
            .I(N__89640));
    LocalMux I__21165 (
            .O(N__89669),
            .I(N__89640));
    Span4Mux_h I__21164 (
            .O(N__89666),
            .I(N__89637));
    Sp12to4 I__21163 (
            .O(N__89663),
            .I(N__89634));
    Span4Mux_v I__21162 (
            .O(N__89660),
            .I(N__89629));
    Span4Mux_v I__21161 (
            .O(N__89657),
            .I(N__89629));
    Span4Mux_h I__21160 (
            .O(N__89652),
            .I(N__89626));
    Span4Mux_h I__21159 (
            .O(N__89645),
            .I(N__89623));
    Span4Mux_h I__21158 (
            .O(N__89640),
            .I(N__89620));
    Span4Mux_h I__21157 (
            .O(N__89637),
            .I(N__89617));
    Span12Mux_v I__21156 (
            .O(N__89634),
            .I(N__89614));
    Sp12to4 I__21155 (
            .O(N__89629),
            .I(N__89611));
    Span4Mux_v I__21154 (
            .O(N__89626),
            .I(N__89608));
    Span4Mux_h I__21153 (
            .O(N__89623),
            .I(N__89605));
    Sp12to4 I__21152 (
            .O(N__89620),
            .I(N__89596));
    Sp12to4 I__21151 (
            .O(N__89617),
            .I(N__89596));
    Span12Mux_h I__21150 (
            .O(N__89614),
            .I(N__89596));
    Span12Mux_h I__21149 (
            .O(N__89611),
            .I(N__89596));
    Odrv4 I__21148 (
            .O(N__89608),
            .I(\c0.n9_adj_4552 ));
    Odrv4 I__21147 (
            .O(N__89605),
            .I(\c0.n9_adj_4552 ));
    Odrv12 I__21146 (
            .O(N__89596),
            .I(\c0.n9_adj_4552 ));
    CascadeMux I__21145 (
            .O(N__89589),
            .I(\quad_counter1.n29_adj_4428_cascade_ ));
    InMux I__21144 (
            .O(N__89586),
            .I(N__89583));
    LocalMux I__21143 (
            .O(N__89583),
            .I(\quad_counter1.n27_adj_4429 ));
    CascadeMux I__21142 (
            .O(N__89580),
            .I(N__89561));
    CascadeMux I__21141 (
            .O(N__89579),
            .I(N__89558));
    CascadeMux I__21140 (
            .O(N__89578),
            .I(N__89555));
    CascadeMux I__21139 (
            .O(N__89577),
            .I(N__89552));
    CascadeMux I__21138 (
            .O(N__89576),
            .I(N__89549));
    CascadeMux I__21137 (
            .O(N__89575),
            .I(N__89546));
    CascadeMux I__21136 (
            .O(N__89574),
            .I(N__89543));
    CascadeMux I__21135 (
            .O(N__89573),
            .I(N__89540));
    CascadeMux I__21134 (
            .O(N__89572),
            .I(N__89537));
    CascadeMux I__21133 (
            .O(N__89571),
            .I(N__89534));
    CascadeMux I__21132 (
            .O(N__89570),
            .I(N__89531));
    CascadeMux I__21131 (
            .O(N__89569),
            .I(N__89528));
    CascadeMux I__21130 (
            .O(N__89568),
            .I(N__89525));
    CascadeMux I__21129 (
            .O(N__89567),
            .I(N__89522));
    CascadeMux I__21128 (
            .O(N__89566),
            .I(N__89519));
    CascadeMux I__21127 (
            .O(N__89565),
            .I(N__89516));
    CascadeMux I__21126 (
            .O(N__89564),
            .I(N__89513));
    InMux I__21125 (
            .O(N__89561),
            .I(N__89506));
    InMux I__21124 (
            .O(N__89558),
            .I(N__89506));
    InMux I__21123 (
            .O(N__89555),
            .I(N__89506));
    InMux I__21122 (
            .O(N__89552),
            .I(N__89497));
    InMux I__21121 (
            .O(N__89549),
            .I(N__89497));
    InMux I__21120 (
            .O(N__89546),
            .I(N__89497));
    InMux I__21119 (
            .O(N__89543),
            .I(N__89497));
    InMux I__21118 (
            .O(N__89540),
            .I(N__89488));
    InMux I__21117 (
            .O(N__89537),
            .I(N__89488));
    InMux I__21116 (
            .O(N__89534),
            .I(N__89488));
    InMux I__21115 (
            .O(N__89531),
            .I(N__89488));
    InMux I__21114 (
            .O(N__89528),
            .I(N__89483));
    InMux I__21113 (
            .O(N__89525),
            .I(N__89483));
    InMux I__21112 (
            .O(N__89522),
            .I(N__89474));
    InMux I__21111 (
            .O(N__89519),
            .I(N__89474));
    InMux I__21110 (
            .O(N__89516),
            .I(N__89474));
    InMux I__21109 (
            .O(N__89513),
            .I(N__89474));
    LocalMux I__21108 (
            .O(N__89506),
            .I(N__89467));
    LocalMux I__21107 (
            .O(N__89497),
            .I(N__89467));
    LocalMux I__21106 (
            .O(N__89488),
            .I(N__89467));
    LocalMux I__21105 (
            .O(N__89483),
            .I(N__89464));
    LocalMux I__21104 (
            .O(N__89474),
            .I(\quad_counter1.n3431 ));
    Odrv4 I__21103 (
            .O(N__89467),
            .I(\quad_counter1.n3431 ));
    Odrv4 I__21102 (
            .O(N__89464),
            .I(\quad_counter1.n3431 ));
    CascadeMux I__21101 (
            .O(N__89457),
            .I(\quad_counter1.n3431_cascade_ ));
    CascadeMux I__21100 (
            .O(N__89454),
            .I(N__89446));
    CascadeMux I__21099 (
            .O(N__89453),
            .I(N__89443));
    CascadeMux I__21098 (
            .O(N__89452),
            .I(N__89440));
    CascadeMux I__21097 (
            .O(N__89451),
            .I(N__89437));
    CascadeMux I__21096 (
            .O(N__89450),
            .I(N__89434));
    CascadeMux I__21095 (
            .O(N__89449),
            .I(N__89431));
    InMux I__21094 (
            .O(N__89446),
            .I(N__89426));
    InMux I__21093 (
            .O(N__89443),
            .I(N__89426));
    InMux I__21092 (
            .O(N__89440),
            .I(N__89417));
    InMux I__21091 (
            .O(N__89437),
            .I(N__89417));
    InMux I__21090 (
            .O(N__89434),
            .I(N__89417));
    InMux I__21089 (
            .O(N__89431),
            .I(N__89417));
    LocalMux I__21088 (
            .O(N__89426),
            .I(N__89412));
    LocalMux I__21087 (
            .O(N__89417),
            .I(N__89412));
    Odrv12 I__21086 (
            .O(N__89412),
            .I(\quad_counter1.n36142 ));
    CascadeMux I__21085 (
            .O(N__89409),
            .I(N__89406));
    InMux I__21084 (
            .O(N__89406),
            .I(N__89403));
    LocalMux I__21083 (
            .O(N__89403),
            .I(N__89399));
    InMux I__21082 (
            .O(N__89402),
            .I(N__89396));
    Span4Mux_v I__21081 (
            .O(N__89399),
            .I(N__89391));
    LocalMux I__21080 (
            .O(N__89396),
            .I(N__89388));
    InMux I__21079 (
            .O(N__89395),
            .I(N__89385));
    InMux I__21078 (
            .O(N__89394),
            .I(N__89382));
    Span4Mux_v I__21077 (
            .O(N__89391),
            .I(N__89379));
    Span12Mux_s10_h I__21076 (
            .O(N__89388),
            .I(N__89374));
    LocalMux I__21075 (
            .O(N__89385),
            .I(N__89374));
    LocalMux I__21074 (
            .O(N__89382),
            .I(\quad_counter1.millisecond_counter_8 ));
    Odrv4 I__21073 (
            .O(N__89379),
            .I(\quad_counter1.millisecond_counter_8 ));
    Odrv12 I__21072 (
            .O(N__89374),
            .I(\quad_counter1.millisecond_counter_8 ));
    InMux I__21071 (
            .O(N__89367),
            .I(N__89362));
    InMux I__21070 (
            .O(N__89366),
            .I(N__89359));
    CascadeMux I__21069 (
            .O(N__89365),
            .I(N__89356));
    LocalMux I__21068 (
            .O(N__89362),
            .I(N__89351));
    LocalMux I__21067 (
            .O(N__89359),
            .I(N__89351));
    InMux I__21066 (
            .O(N__89356),
            .I(N__89348));
    Odrv12 I__21065 (
            .O(N__89351),
            .I(\quad_counter1.n3519 ));
    LocalMux I__21064 (
            .O(N__89348),
            .I(\quad_counter1.n3519 ));
    InMux I__21063 (
            .O(N__89343),
            .I(N__89339));
    InMux I__21062 (
            .O(N__89342),
            .I(N__89335));
    LocalMux I__21061 (
            .O(N__89339),
            .I(N__89332));
    InMux I__21060 (
            .O(N__89338),
            .I(N__89329));
    LocalMux I__21059 (
            .O(N__89335),
            .I(N__89326));
    Odrv4 I__21058 (
            .O(N__89332),
            .I(\quad_counter1.n3514 ));
    LocalMux I__21057 (
            .O(N__89329),
            .I(\quad_counter1.n3514 ));
    Odrv12 I__21056 (
            .O(N__89326),
            .I(\quad_counter1.n3514 ));
    InMux I__21055 (
            .O(N__89319),
            .I(N__89314));
    InMux I__21054 (
            .O(N__89318),
            .I(N__89311));
    CascadeMux I__21053 (
            .O(N__89317),
            .I(N__89308));
    LocalMux I__21052 (
            .O(N__89314),
            .I(N__89303));
    LocalMux I__21051 (
            .O(N__89311),
            .I(N__89303));
    InMux I__21050 (
            .O(N__89308),
            .I(N__89300));
    Odrv12 I__21049 (
            .O(N__89303),
            .I(\quad_counter1.n3517 ));
    LocalMux I__21048 (
            .O(N__89300),
            .I(\quad_counter1.n3517 ));
    CascadeMux I__21047 (
            .O(N__89295),
            .I(\quad_counter1.n28415_cascade_ ));
    InMux I__21046 (
            .O(N__89292),
            .I(N__89287));
    InMux I__21045 (
            .O(N__89291),
            .I(N__89284));
    CascadeMux I__21044 (
            .O(N__89290),
            .I(N__89281));
    LocalMux I__21043 (
            .O(N__89287),
            .I(N__89276));
    LocalMux I__21042 (
            .O(N__89284),
            .I(N__89276));
    InMux I__21041 (
            .O(N__89281),
            .I(N__89273));
    Odrv12 I__21040 (
            .O(N__89276),
            .I(\quad_counter1.n3518 ));
    LocalMux I__21039 (
            .O(N__89273),
            .I(\quad_counter1.n3518 ));
    InMux I__21038 (
            .O(N__89268),
            .I(N__89264));
    InMux I__21037 (
            .O(N__89267),
            .I(N__89260));
    LocalMux I__21036 (
            .O(N__89264),
            .I(N__89257));
    InMux I__21035 (
            .O(N__89263),
            .I(N__89254));
    LocalMux I__21034 (
            .O(N__89260),
            .I(N__89251));
    Odrv4 I__21033 (
            .O(N__89257),
            .I(\quad_counter1.n3515 ));
    LocalMux I__21032 (
            .O(N__89254),
            .I(\quad_counter1.n3515 ));
    Odrv12 I__21031 (
            .O(N__89251),
            .I(\quad_counter1.n3515 ));
    InMux I__21030 (
            .O(N__89244),
            .I(N__89241));
    LocalMux I__21029 (
            .O(N__89241),
            .I(N__89238));
    Odrv4 I__21028 (
            .O(N__89238),
            .I(\quad_counter1.n3509 ));
    CascadeMux I__21027 (
            .O(N__89235),
            .I(\quad_counter1.n10_adj_4462_cascade_ ));
    InMux I__21026 (
            .O(N__89232),
            .I(N__89227));
    InMux I__21025 (
            .O(N__89231),
            .I(N__89224));
    CascadeMux I__21024 (
            .O(N__89230),
            .I(N__89221));
    LocalMux I__21023 (
            .O(N__89227),
            .I(N__89216));
    LocalMux I__21022 (
            .O(N__89224),
            .I(N__89216));
    InMux I__21021 (
            .O(N__89221),
            .I(N__89213));
    Odrv12 I__21020 (
            .O(N__89216),
            .I(\quad_counter1.n3516 ));
    LocalMux I__21019 (
            .O(N__89213),
            .I(\quad_counter1.n3516 ));
    InMux I__21018 (
            .O(N__89208),
            .I(N__89205));
    LocalMux I__21017 (
            .O(N__89205),
            .I(\quad_counter1.n21 ));
    InMux I__21016 (
            .O(N__89202),
            .I(N__89199));
    LocalMux I__21015 (
            .O(N__89199),
            .I(N__89195));
    InMux I__21014 (
            .O(N__89198),
            .I(N__89192));
    Span4Mux_h I__21013 (
            .O(N__89195),
            .I(N__89189));
    LocalMux I__21012 (
            .O(N__89192),
            .I(data_out_frame_13_2));
    Odrv4 I__21011 (
            .O(N__89189),
            .I(data_out_frame_13_2));
    InMux I__21010 (
            .O(N__89184),
            .I(N__89181));
    LocalMux I__21009 (
            .O(N__89181),
            .I(N__89177));
    InMux I__21008 (
            .O(N__89180),
            .I(N__89174));
    Span4Mux_v I__21007 (
            .O(N__89177),
            .I(N__89171));
    LocalMux I__21006 (
            .O(N__89174),
            .I(data_out_frame_12_2));
    Odrv4 I__21005 (
            .O(N__89171),
            .I(data_out_frame_12_2));
    InMux I__21004 (
            .O(N__89166),
            .I(N__89163));
    LocalMux I__21003 (
            .O(N__89163),
            .I(N__89160));
    Span4Mux_v I__21002 (
            .O(N__89160),
            .I(N__89157));
    Span4Mux_h I__21001 (
            .O(N__89157),
            .I(N__89154));
    Span4Mux_h I__21000 (
            .O(N__89154),
            .I(N__89151));
    Odrv4 I__20999 (
            .O(N__89151),
            .I(\c0.n11_adj_4513 ));
    InMux I__20998 (
            .O(N__89148),
            .I(\quad_counter1.n30693 ));
    CascadeMux I__20997 (
            .O(N__89145),
            .I(N__89140));
    InMux I__20996 (
            .O(N__89144),
            .I(N__89137));
    InMux I__20995 (
            .O(N__89143),
            .I(N__89134));
    InMux I__20994 (
            .O(N__89140),
            .I(N__89131));
    LocalMux I__20993 (
            .O(N__89137),
            .I(\quad_counter1.n3400 ));
    LocalMux I__20992 (
            .O(N__89134),
            .I(\quad_counter1.n3400 ));
    LocalMux I__20991 (
            .O(N__89131),
            .I(\quad_counter1.n3400 ));
    InMux I__20990 (
            .O(N__89124),
            .I(N__89121));
    LocalMux I__20989 (
            .O(N__89121),
            .I(N__89118));
    Odrv4 I__20988 (
            .O(N__89118),
            .I(\quad_counter1.n3499 ));
    InMux I__20987 (
            .O(N__89115),
            .I(\quad_counter1.n30694 ));
    InMux I__20986 (
            .O(N__89112),
            .I(N__89107));
    InMux I__20985 (
            .O(N__89111),
            .I(N__89104));
    InMux I__20984 (
            .O(N__89110),
            .I(N__89101));
    LocalMux I__20983 (
            .O(N__89107),
            .I(\quad_counter1.n3399 ));
    LocalMux I__20982 (
            .O(N__89104),
            .I(\quad_counter1.n3399 ));
    LocalMux I__20981 (
            .O(N__89101),
            .I(\quad_counter1.n3399 ));
    InMux I__20980 (
            .O(N__89094),
            .I(N__89091));
    LocalMux I__20979 (
            .O(N__89091),
            .I(N__89088));
    Odrv4 I__20978 (
            .O(N__89088),
            .I(\quad_counter1.n3498 ));
    InMux I__20977 (
            .O(N__89085),
            .I(\quad_counter1.n30695 ));
    InMux I__20976 (
            .O(N__89082),
            .I(N__89077));
    InMux I__20975 (
            .O(N__89081),
            .I(N__89074));
    InMux I__20974 (
            .O(N__89080),
            .I(N__89071));
    LocalMux I__20973 (
            .O(N__89077),
            .I(\quad_counter1.n3398 ));
    LocalMux I__20972 (
            .O(N__89074),
            .I(\quad_counter1.n3398 ));
    LocalMux I__20971 (
            .O(N__89071),
            .I(\quad_counter1.n3398 ));
    InMux I__20970 (
            .O(N__89064),
            .I(\quad_counter1.n30696 ));
    InMux I__20969 (
            .O(N__89061),
            .I(N__89058));
    LocalMux I__20968 (
            .O(N__89058),
            .I(\quad_counter1.n3506 ));
    InMux I__20967 (
            .O(N__89055),
            .I(N__89052));
    LocalMux I__20966 (
            .O(N__89052),
            .I(\quad_counter1.n3511 ));
    CascadeMux I__20965 (
            .O(N__89049),
            .I(\quad_counter1.n3497_cascade_ ));
    InMux I__20964 (
            .O(N__89046),
            .I(N__89043));
    LocalMux I__20963 (
            .O(N__89043),
            .I(\quad_counter1.n3505 ));
    InMux I__20962 (
            .O(N__89040),
            .I(N__89037));
    LocalMux I__20961 (
            .O(N__89037),
            .I(N__89034));
    Odrv4 I__20960 (
            .O(N__89034),
            .I(\quad_counter1.n30_adj_4463 ));
    CascadeMux I__20959 (
            .O(N__89031),
            .I(\quad_counter1.n12_adj_4464_cascade_ ));
    InMux I__20958 (
            .O(N__89028),
            .I(N__89025));
    LocalMux I__20957 (
            .O(N__89025),
            .I(N__89022));
    Odrv4 I__20956 (
            .O(N__89022),
            .I(\quad_counter1.n35985 ));
    InMux I__20955 (
            .O(N__89019),
            .I(N__89014));
    InMux I__20954 (
            .O(N__89018),
            .I(N__89011));
    InMux I__20953 (
            .O(N__89017),
            .I(N__89008));
    LocalMux I__20952 (
            .O(N__89014),
            .I(\quad_counter1.n3407 ));
    LocalMux I__20951 (
            .O(N__89011),
            .I(\quad_counter1.n3407 ));
    LocalMux I__20950 (
            .O(N__89008),
            .I(\quad_counter1.n3407 ));
    InMux I__20949 (
            .O(N__89001),
            .I(N__88996));
    InMux I__20948 (
            .O(N__89000),
            .I(N__88993));
    InMux I__20947 (
            .O(N__88999),
            .I(N__88990));
    LocalMux I__20946 (
            .O(N__88996),
            .I(\quad_counter1.n3405 ));
    LocalMux I__20945 (
            .O(N__88993),
            .I(\quad_counter1.n3405 ));
    LocalMux I__20944 (
            .O(N__88990),
            .I(\quad_counter1.n3405 ));
    CascadeMux I__20943 (
            .O(N__88983),
            .I(N__88978));
    InMux I__20942 (
            .O(N__88982),
            .I(N__88975));
    InMux I__20941 (
            .O(N__88981),
            .I(N__88972));
    InMux I__20940 (
            .O(N__88978),
            .I(N__88969));
    LocalMux I__20939 (
            .O(N__88975),
            .I(\quad_counter1.n3411 ));
    LocalMux I__20938 (
            .O(N__88972),
            .I(\quad_counter1.n3411 ));
    LocalMux I__20937 (
            .O(N__88969),
            .I(\quad_counter1.n3411 ));
    InMux I__20936 (
            .O(N__88962),
            .I(N__88959));
    LocalMux I__20935 (
            .O(N__88959),
            .I(N__88954));
    InMux I__20934 (
            .O(N__88958),
            .I(N__88951));
    InMux I__20933 (
            .O(N__88957),
            .I(N__88948));
    Span4Mux_v I__20932 (
            .O(N__88954),
            .I(N__88945));
    LocalMux I__20931 (
            .O(N__88951),
            .I(\quad_counter1.n3413 ));
    LocalMux I__20930 (
            .O(N__88948),
            .I(\quad_counter1.n3413 ));
    Odrv4 I__20929 (
            .O(N__88945),
            .I(\quad_counter1.n3413 ));
    InMux I__20928 (
            .O(N__88938),
            .I(N__88935));
    LocalMux I__20927 (
            .O(N__88935),
            .I(N__88932));
    Span4Mux_v I__20926 (
            .O(N__88932),
            .I(N__88929));
    Odrv4 I__20925 (
            .O(N__88929),
            .I(\quad_counter1.n30_adj_4426 ));
    InMux I__20924 (
            .O(N__88926),
            .I(N__88923));
    LocalMux I__20923 (
            .O(N__88923),
            .I(\quad_counter1.n28_adj_4427 ));
    InMux I__20922 (
            .O(N__88920),
            .I(N__88917));
    LocalMux I__20921 (
            .O(N__88917),
            .I(\quad_counter1.n3508 ));
    InMux I__20920 (
            .O(N__88914),
            .I(\quad_counter1.n30685 ));
    InMux I__20919 (
            .O(N__88911),
            .I(N__88907));
    InMux I__20918 (
            .O(N__88910),
            .I(N__88903));
    LocalMux I__20917 (
            .O(N__88907),
            .I(N__88900));
    InMux I__20916 (
            .O(N__88906),
            .I(N__88897));
    LocalMux I__20915 (
            .O(N__88903),
            .I(\quad_counter1.n3408 ));
    Odrv4 I__20914 (
            .O(N__88900),
            .I(\quad_counter1.n3408 ));
    LocalMux I__20913 (
            .O(N__88897),
            .I(\quad_counter1.n3408 ));
    InMux I__20912 (
            .O(N__88890),
            .I(N__88887));
    LocalMux I__20911 (
            .O(N__88887),
            .I(N__88884));
    Odrv4 I__20910 (
            .O(N__88884),
            .I(\quad_counter1.n3507 ));
    InMux I__20909 (
            .O(N__88881),
            .I(\quad_counter1.n30686 ));
    InMux I__20908 (
            .O(N__88878),
            .I(\quad_counter1.n30687 ));
    CascadeMux I__20907 (
            .O(N__88875),
            .I(N__88870));
    InMux I__20906 (
            .O(N__88874),
            .I(N__88867));
    InMux I__20905 (
            .O(N__88873),
            .I(N__88864));
    InMux I__20904 (
            .O(N__88870),
            .I(N__88861));
    LocalMux I__20903 (
            .O(N__88867),
            .I(\quad_counter1.n3406 ));
    LocalMux I__20902 (
            .O(N__88864),
            .I(\quad_counter1.n3406 ));
    LocalMux I__20901 (
            .O(N__88861),
            .I(\quad_counter1.n3406 ));
    InMux I__20900 (
            .O(N__88854),
            .I(\quad_counter1.n30688 ));
    CascadeMux I__20899 (
            .O(N__88851),
            .I(N__88848));
    InMux I__20898 (
            .O(N__88848),
            .I(N__88845));
    LocalMux I__20897 (
            .O(N__88845),
            .I(\quad_counter1.n3504 ));
    InMux I__20896 (
            .O(N__88842),
            .I(\quad_counter1.n30689 ));
    InMux I__20895 (
            .O(N__88839),
            .I(N__88834));
    InMux I__20894 (
            .O(N__88838),
            .I(N__88831));
    InMux I__20893 (
            .O(N__88837),
            .I(N__88828));
    LocalMux I__20892 (
            .O(N__88834),
            .I(\quad_counter1.n3404 ));
    LocalMux I__20891 (
            .O(N__88831),
            .I(\quad_counter1.n3404 ));
    LocalMux I__20890 (
            .O(N__88828),
            .I(\quad_counter1.n3404 ));
    CascadeMux I__20889 (
            .O(N__88821),
            .I(N__88818));
    InMux I__20888 (
            .O(N__88818),
            .I(N__88815));
    LocalMux I__20887 (
            .O(N__88815),
            .I(N__88812));
    Odrv4 I__20886 (
            .O(N__88812),
            .I(\quad_counter1.n3503 ));
    InMux I__20885 (
            .O(N__88809),
            .I(bfn_23_14_0_));
    InMux I__20884 (
            .O(N__88806),
            .I(N__88801));
    InMux I__20883 (
            .O(N__88805),
            .I(N__88798));
    InMux I__20882 (
            .O(N__88804),
            .I(N__88795));
    LocalMux I__20881 (
            .O(N__88801),
            .I(\quad_counter1.n3403 ));
    LocalMux I__20880 (
            .O(N__88798),
            .I(\quad_counter1.n3403 ));
    LocalMux I__20879 (
            .O(N__88795),
            .I(\quad_counter1.n3403 ));
    InMux I__20878 (
            .O(N__88788),
            .I(N__88785));
    LocalMux I__20877 (
            .O(N__88785),
            .I(N__88782));
    Odrv4 I__20876 (
            .O(N__88782),
            .I(\quad_counter1.n3502 ));
    InMux I__20875 (
            .O(N__88779),
            .I(\quad_counter1.n30691 ));
    InMux I__20874 (
            .O(N__88776),
            .I(N__88771));
    InMux I__20873 (
            .O(N__88775),
            .I(N__88768));
    InMux I__20872 (
            .O(N__88774),
            .I(N__88765));
    LocalMux I__20871 (
            .O(N__88771),
            .I(N__88762));
    LocalMux I__20870 (
            .O(N__88768),
            .I(\quad_counter1.n3402 ));
    LocalMux I__20869 (
            .O(N__88765),
            .I(\quad_counter1.n3402 ));
    Odrv4 I__20868 (
            .O(N__88762),
            .I(\quad_counter1.n3402 ));
    InMux I__20867 (
            .O(N__88755),
            .I(N__88752));
    LocalMux I__20866 (
            .O(N__88752),
            .I(N__88749));
    Odrv4 I__20865 (
            .O(N__88749),
            .I(\quad_counter1.n3501 ));
    InMux I__20864 (
            .O(N__88746),
            .I(\quad_counter1.n30692 ));
    InMux I__20863 (
            .O(N__88743),
            .I(N__88738));
    InMux I__20862 (
            .O(N__88742),
            .I(N__88735));
    InMux I__20861 (
            .O(N__88741),
            .I(N__88732));
    LocalMux I__20860 (
            .O(N__88738),
            .I(\quad_counter1.n3401 ));
    LocalMux I__20859 (
            .O(N__88735),
            .I(\quad_counter1.n3401 ));
    LocalMux I__20858 (
            .O(N__88732),
            .I(\quad_counter1.n3401 ));
    InMux I__20857 (
            .O(N__88725),
            .I(N__88722));
    LocalMux I__20856 (
            .O(N__88722),
            .I(N__88719));
    Odrv4 I__20855 (
            .O(N__88719),
            .I(\quad_counter1.n3500 ));
    InMux I__20854 (
            .O(N__88716),
            .I(N__88711));
    InMux I__20853 (
            .O(N__88715),
            .I(N__88708));
    InMux I__20852 (
            .O(N__88714),
            .I(N__88705));
    LocalMux I__20851 (
            .O(N__88711),
            .I(\quad_counter1.n3417 ));
    LocalMux I__20850 (
            .O(N__88708),
            .I(\quad_counter1.n3417 ));
    LocalMux I__20849 (
            .O(N__88705),
            .I(\quad_counter1.n3417 ));
    InMux I__20848 (
            .O(N__88698),
            .I(\quad_counter1.n30677 ));
    InMux I__20847 (
            .O(N__88695),
            .I(N__88691));
    InMux I__20846 (
            .O(N__88694),
            .I(N__88688));
    LocalMux I__20845 (
            .O(N__88691),
            .I(N__88682));
    LocalMux I__20844 (
            .O(N__88688),
            .I(N__88682));
    InMux I__20843 (
            .O(N__88687),
            .I(N__88679));
    Odrv4 I__20842 (
            .O(N__88682),
            .I(\quad_counter1.n3416 ));
    LocalMux I__20841 (
            .O(N__88679),
            .I(\quad_counter1.n3416 ));
    InMux I__20840 (
            .O(N__88674),
            .I(\quad_counter1.n30678 ));
    InMux I__20839 (
            .O(N__88671),
            .I(N__88666));
    InMux I__20838 (
            .O(N__88670),
            .I(N__88663));
    InMux I__20837 (
            .O(N__88669),
            .I(N__88660));
    LocalMux I__20836 (
            .O(N__88666),
            .I(\quad_counter1.n3415 ));
    LocalMux I__20835 (
            .O(N__88663),
            .I(\quad_counter1.n3415 ));
    LocalMux I__20834 (
            .O(N__88660),
            .I(\quad_counter1.n3415 ));
    InMux I__20833 (
            .O(N__88653),
            .I(\quad_counter1.n30679 ));
    InMux I__20832 (
            .O(N__88650),
            .I(N__88645));
    InMux I__20831 (
            .O(N__88649),
            .I(N__88642));
    InMux I__20830 (
            .O(N__88648),
            .I(N__88639));
    LocalMux I__20829 (
            .O(N__88645),
            .I(\quad_counter1.n3414 ));
    LocalMux I__20828 (
            .O(N__88642),
            .I(\quad_counter1.n3414 ));
    LocalMux I__20827 (
            .O(N__88639),
            .I(\quad_counter1.n3414 ));
    InMux I__20826 (
            .O(N__88632),
            .I(N__88629));
    LocalMux I__20825 (
            .O(N__88629),
            .I(\quad_counter1.n3513 ));
    InMux I__20824 (
            .O(N__88626),
            .I(\quad_counter1.n30680 ));
    CascadeMux I__20823 (
            .O(N__88623),
            .I(N__88620));
    InMux I__20822 (
            .O(N__88620),
            .I(N__88617));
    LocalMux I__20821 (
            .O(N__88617),
            .I(\quad_counter1.n3512 ));
    InMux I__20820 (
            .O(N__88614),
            .I(\quad_counter1.n30681 ));
    CascadeMux I__20819 (
            .O(N__88611),
            .I(N__88608));
    InMux I__20818 (
            .O(N__88608),
            .I(N__88603));
    InMux I__20817 (
            .O(N__88607),
            .I(N__88600));
    InMux I__20816 (
            .O(N__88606),
            .I(N__88597));
    LocalMux I__20815 (
            .O(N__88603),
            .I(N__88594));
    LocalMux I__20814 (
            .O(N__88600),
            .I(\quad_counter1.n3412 ));
    LocalMux I__20813 (
            .O(N__88597),
            .I(\quad_counter1.n3412 ));
    Odrv4 I__20812 (
            .O(N__88594),
            .I(\quad_counter1.n3412 ));
    InMux I__20811 (
            .O(N__88587),
            .I(bfn_23_13_0_));
    InMux I__20810 (
            .O(N__88584),
            .I(N__88581));
    LocalMux I__20809 (
            .O(N__88581),
            .I(N__88578));
    Span4Mux_v I__20808 (
            .O(N__88578),
            .I(N__88575));
    Odrv4 I__20807 (
            .O(N__88575),
            .I(\quad_counter1.n3510 ));
    InMux I__20806 (
            .O(N__88572),
            .I(\quad_counter1.n30683 ));
    InMux I__20805 (
            .O(N__88569),
            .I(N__88564));
    InMux I__20804 (
            .O(N__88568),
            .I(N__88561));
    InMux I__20803 (
            .O(N__88567),
            .I(N__88558));
    LocalMux I__20802 (
            .O(N__88564),
            .I(\quad_counter1.n3410 ));
    LocalMux I__20801 (
            .O(N__88561),
            .I(\quad_counter1.n3410 ));
    LocalMux I__20800 (
            .O(N__88558),
            .I(\quad_counter1.n3410 ));
    InMux I__20799 (
            .O(N__88551),
            .I(\quad_counter1.n30684 ));
    InMux I__20798 (
            .O(N__88548),
            .I(N__88543));
    InMux I__20797 (
            .O(N__88547),
            .I(N__88540));
    InMux I__20796 (
            .O(N__88546),
            .I(N__88537));
    LocalMux I__20795 (
            .O(N__88543),
            .I(\quad_counter1.n3409 ));
    LocalMux I__20794 (
            .O(N__88540),
            .I(\quad_counter1.n3409 ));
    LocalMux I__20793 (
            .O(N__88537),
            .I(\quad_counter1.n3409 ));
    CascadeMux I__20792 (
            .O(N__88530),
            .I(N__88522));
    CascadeMux I__20791 (
            .O(N__88529),
            .I(N__88519));
    CascadeMux I__20790 (
            .O(N__88528),
            .I(N__88516));
    CascadeMux I__20789 (
            .O(N__88527),
            .I(N__88513));
    CascadeMux I__20788 (
            .O(N__88526),
            .I(N__88510));
    CascadeMux I__20787 (
            .O(N__88525),
            .I(N__88507));
    InMux I__20786 (
            .O(N__88522),
            .I(N__88502));
    InMux I__20785 (
            .O(N__88519),
            .I(N__88502));
    InMux I__20784 (
            .O(N__88516),
            .I(N__88493));
    InMux I__20783 (
            .O(N__88513),
            .I(N__88493));
    InMux I__20782 (
            .O(N__88510),
            .I(N__88493));
    InMux I__20781 (
            .O(N__88507),
            .I(N__88493));
    LocalMux I__20780 (
            .O(N__88502),
            .I(\quad_counter1.n36135 ));
    LocalMux I__20779 (
            .O(N__88493),
            .I(\quad_counter1.n36135 ));
    InMux I__20778 (
            .O(N__88488),
            .I(N__88485));
    LocalMux I__20777 (
            .O(N__88485),
            .I(\quad_counter1.n28_adj_4460 ));
    InMux I__20776 (
            .O(N__88482),
            .I(N__88479));
    LocalMux I__20775 (
            .O(N__88479),
            .I(N__88473));
    InMux I__20774 (
            .O(N__88478),
            .I(N__88470));
    InMux I__20773 (
            .O(N__88477),
            .I(N__88467));
    InMux I__20772 (
            .O(N__88476),
            .I(N__88464));
    Span4Mux_v I__20771 (
            .O(N__88473),
            .I(N__88461));
    LocalMux I__20770 (
            .O(N__88470),
            .I(\quad_counter1.millisecond_counter_20 ));
    LocalMux I__20769 (
            .O(N__88467),
            .I(\quad_counter1.millisecond_counter_20 ));
    LocalMux I__20768 (
            .O(N__88464),
            .I(\quad_counter1.millisecond_counter_20 ));
    Odrv4 I__20767 (
            .O(N__88461),
            .I(\quad_counter1.millisecond_counter_20 ));
    CascadeMux I__20766 (
            .O(N__88452),
            .I(\quad_counter1.n28277_cascade_ ));
    CascadeMux I__20765 (
            .O(N__88449),
            .I(\quad_counter1.n10_adj_4437_cascade_ ));
    CascadeMux I__20764 (
            .O(N__88446),
            .I(\quad_counter1.n7_adj_4439_cascade_ ));
    CascadeMux I__20763 (
            .O(N__88443),
            .I(N__88437));
    CascadeMux I__20762 (
            .O(N__88442),
            .I(N__88434));
    CascadeMux I__20761 (
            .O(N__88441),
            .I(N__88429));
    CascadeMux I__20760 (
            .O(N__88440),
            .I(N__88426));
    InMux I__20759 (
            .O(N__88437),
            .I(N__88421));
    InMux I__20758 (
            .O(N__88434),
            .I(N__88421));
    CascadeMux I__20757 (
            .O(N__88433),
            .I(N__88418));
    CascadeMux I__20756 (
            .O(N__88432),
            .I(N__88415));
    InMux I__20755 (
            .O(N__88429),
            .I(N__88409));
    InMux I__20754 (
            .O(N__88426),
            .I(N__88409));
    LocalMux I__20753 (
            .O(N__88421),
            .I(N__88406));
    InMux I__20752 (
            .O(N__88418),
            .I(N__88399));
    InMux I__20751 (
            .O(N__88415),
            .I(N__88399));
    InMux I__20750 (
            .O(N__88414),
            .I(N__88399));
    LocalMux I__20749 (
            .O(N__88409),
            .I(\quad_counter1.n2342 ));
    Odrv4 I__20748 (
            .O(N__88406),
            .I(\quad_counter1.n2342 ));
    LocalMux I__20747 (
            .O(N__88399),
            .I(\quad_counter1.n2342 ));
    InMux I__20746 (
            .O(N__88392),
            .I(N__88387));
    InMux I__20745 (
            .O(N__88391),
            .I(N__88384));
    InMux I__20744 (
            .O(N__88390),
            .I(N__88381));
    LocalMux I__20743 (
            .O(N__88387),
            .I(N__88375));
    LocalMux I__20742 (
            .O(N__88384),
            .I(N__88375));
    LocalMux I__20741 (
            .O(N__88381),
            .I(N__88372));
    InMux I__20740 (
            .O(N__88380),
            .I(N__88369));
    Span4Mux_v I__20739 (
            .O(N__88375),
            .I(N__88366));
    Span4Mux_v I__20738 (
            .O(N__88372),
            .I(N__88363));
    LocalMux I__20737 (
            .O(N__88369),
            .I(\quad_counter1.millisecond_counter_9 ));
    Odrv4 I__20736 (
            .O(N__88366),
            .I(\quad_counter1.millisecond_counter_9 ));
    Odrv4 I__20735 (
            .O(N__88363),
            .I(\quad_counter1.millisecond_counter_9 ));
    InMux I__20734 (
            .O(N__88356),
            .I(bfn_23_12_0_));
    CascadeMux I__20733 (
            .O(N__88353),
            .I(N__88348));
    InMux I__20732 (
            .O(N__88352),
            .I(N__88345));
    InMux I__20731 (
            .O(N__88351),
            .I(N__88342));
    InMux I__20730 (
            .O(N__88348),
            .I(N__88339));
    LocalMux I__20729 (
            .O(N__88345),
            .I(\quad_counter1.n3419 ));
    LocalMux I__20728 (
            .O(N__88342),
            .I(\quad_counter1.n3419 ));
    LocalMux I__20727 (
            .O(N__88339),
            .I(\quad_counter1.n3419 ));
    InMux I__20726 (
            .O(N__88332),
            .I(\quad_counter1.n30675 ));
    InMux I__20725 (
            .O(N__88329),
            .I(N__88324));
    InMux I__20724 (
            .O(N__88328),
            .I(N__88321));
    InMux I__20723 (
            .O(N__88327),
            .I(N__88318));
    LocalMux I__20722 (
            .O(N__88324),
            .I(\quad_counter1.n3418 ));
    LocalMux I__20721 (
            .O(N__88321),
            .I(\quad_counter1.n3418 ));
    LocalMux I__20720 (
            .O(N__88318),
            .I(\quad_counter1.n3418 ));
    InMux I__20719 (
            .O(N__88311),
            .I(\quad_counter1.n30676 ));
    InMux I__20718 (
            .O(N__88308),
            .I(N__88303));
    InMux I__20717 (
            .O(N__88307),
            .I(N__88300));
    InMux I__20716 (
            .O(N__88306),
            .I(N__88297));
    LocalMux I__20715 (
            .O(N__88303),
            .I(N__88292));
    LocalMux I__20714 (
            .O(N__88300),
            .I(N__88292));
    LocalMux I__20713 (
            .O(N__88297),
            .I(N__88289));
    Span4Mux_h I__20712 (
            .O(N__88292),
            .I(N__88286));
    Span4Mux_h I__20711 (
            .O(N__88289),
            .I(N__88283));
    Odrv4 I__20710 (
            .O(N__88286),
            .I(\quad_counter1.n2413 ));
    Odrv4 I__20709 (
            .O(N__88283),
            .I(\quad_counter1.n2413 ));
    InMux I__20708 (
            .O(N__88278),
            .I(\quad_counter1.n30504 ));
    InMux I__20707 (
            .O(N__88275),
            .I(N__88270));
    InMux I__20706 (
            .O(N__88274),
            .I(N__88267));
    InMux I__20705 (
            .O(N__88273),
            .I(N__88264));
    LocalMux I__20704 (
            .O(N__88270),
            .I(N__88259));
    LocalMux I__20703 (
            .O(N__88267),
            .I(N__88259));
    LocalMux I__20702 (
            .O(N__88264),
            .I(N__88256));
    Span4Mux_h I__20701 (
            .O(N__88259),
            .I(N__88253));
    Span4Mux_h I__20700 (
            .O(N__88256),
            .I(N__88250));
    Odrv4 I__20699 (
            .O(N__88253),
            .I(\quad_counter1.n2412 ));
    Odrv4 I__20698 (
            .O(N__88250),
            .I(\quad_counter1.n2412 ));
    InMux I__20697 (
            .O(N__88245),
            .I(\quad_counter1.n30505 ));
    InMux I__20696 (
            .O(N__88242),
            .I(N__88237));
    InMux I__20695 (
            .O(N__88241),
            .I(N__88234));
    InMux I__20694 (
            .O(N__88240),
            .I(N__88231));
    LocalMux I__20693 (
            .O(N__88237),
            .I(N__88228));
    LocalMux I__20692 (
            .O(N__88234),
            .I(N__88223));
    LocalMux I__20691 (
            .O(N__88231),
            .I(N__88223));
    Span4Mux_h I__20690 (
            .O(N__88228),
            .I(N__88220));
    Odrv4 I__20689 (
            .O(N__88223),
            .I(\quad_counter1.n2411 ));
    Odrv4 I__20688 (
            .O(N__88220),
            .I(\quad_counter1.n2411 ));
    InMux I__20687 (
            .O(N__88215),
            .I(bfn_23_10_0_));
    CascadeMux I__20686 (
            .O(N__88212),
            .I(N__88209));
    InMux I__20685 (
            .O(N__88209),
            .I(N__88204));
    InMux I__20684 (
            .O(N__88208),
            .I(N__88201));
    InMux I__20683 (
            .O(N__88207),
            .I(N__88198));
    LocalMux I__20682 (
            .O(N__88204),
            .I(N__88195));
    LocalMux I__20681 (
            .O(N__88201),
            .I(N__88190));
    LocalMux I__20680 (
            .O(N__88198),
            .I(N__88190));
    Span4Mux_h I__20679 (
            .O(N__88195),
            .I(N__88187));
    Odrv4 I__20678 (
            .O(N__88190),
            .I(\quad_counter1.n2410 ));
    Odrv4 I__20677 (
            .O(N__88187),
            .I(\quad_counter1.n2410 ));
    InMux I__20676 (
            .O(N__88182),
            .I(\quad_counter1.n30507 ));
    InMux I__20675 (
            .O(N__88179),
            .I(N__88174));
    InMux I__20674 (
            .O(N__88178),
            .I(N__88171));
    InMux I__20673 (
            .O(N__88177),
            .I(N__88168));
    LocalMux I__20672 (
            .O(N__88174),
            .I(N__88165));
    LocalMux I__20671 (
            .O(N__88171),
            .I(N__88158));
    LocalMux I__20670 (
            .O(N__88168),
            .I(N__88158));
    Span4Mux_v I__20669 (
            .O(N__88165),
            .I(N__88158));
    Odrv4 I__20668 (
            .O(N__88158),
            .I(\quad_counter1.n2409 ));
    InMux I__20667 (
            .O(N__88155),
            .I(\quad_counter1.n30508 ));
    InMux I__20666 (
            .O(N__88152),
            .I(\quad_counter1.n30509 ));
    InMux I__20665 (
            .O(N__88149),
            .I(N__88144));
    InMux I__20664 (
            .O(N__88148),
            .I(N__88141));
    InMux I__20663 (
            .O(N__88147),
            .I(N__88138));
    LocalMux I__20662 (
            .O(N__88144),
            .I(N__88135));
    LocalMux I__20661 (
            .O(N__88141),
            .I(N__88128));
    LocalMux I__20660 (
            .O(N__88138),
            .I(N__88128));
    Span4Mux_v I__20659 (
            .O(N__88135),
            .I(N__88128));
    Odrv4 I__20658 (
            .O(N__88128),
            .I(\quad_counter1.n2408 ));
    InMux I__20657 (
            .O(N__88125),
            .I(N__88119));
    InMux I__20656 (
            .O(N__88124),
            .I(N__88116));
    InMux I__20655 (
            .O(N__88123),
            .I(N__88113));
    InMux I__20654 (
            .O(N__88122),
            .I(N__88110));
    LocalMux I__20653 (
            .O(N__88119),
            .I(\quad_counter1.millisecond_counter_19 ));
    LocalMux I__20652 (
            .O(N__88116),
            .I(\quad_counter1.millisecond_counter_19 ));
    LocalMux I__20651 (
            .O(N__88113),
            .I(\quad_counter1.millisecond_counter_19 ));
    LocalMux I__20650 (
            .O(N__88110),
            .I(\quad_counter1.millisecond_counter_19 ));
    InMux I__20649 (
            .O(N__88101),
            .I(N__88097));
    InMux I__20648 (
            .O(N__88100),
            .I(N__88094));
    LocalMux I__20647 (
            .O(N__88097),
            .I(N__88088));
    LocalMux I__20646 (
            .O(N__88094),
            .I(N__88088));
    CascadeMux I__20645 (
            .O(N__88093),
            .I(N__88085));
    Span4Mux_h I__20644 (
            .O(N__88088),
            .I(N__88082));
    InMux I__20643 (
            .O(N__88085),
            .I(N__88079));
    Odrv4 I__20642 (
            .O(N__88082),
            .I(\quad_counter1.n2418 ));
    LocalMux I__20641 (
            .O(N__88079),
            .I(\quad_counter1.n2418 ));
    InMux I__20640 (
            .O(N__88074),
            .I(N__88070));
    InMux I__20639 (
            .O(N__88073),
            .I(N__88067));
    LocalMux I__20638 (
            .O(N__88070),
            .I(N__88062));
    LocalMux I__20637 (
            .O(N__88067),
            .I(N__88062));
    Span4Mux_h I__20636 (
            .O(N__88062),
            .I(N__88058));
    InMux I__20635 (
            .O(N__88061),
            .I(N__88055));
    Odrv4 I__20634 (
            .O(N__88058),
            .I(\quad_counter1.n2419 ));
    LocalMux I__20633 (
            .O(N__88055),
            .I(\quad_counter1.n2419 ));
    CascadeMux I__20632 (
            .O(N__88050),
            .I(N__88047));
    InMux I__20631 (
            .O(N__88047),
            .I(N__88044));
    LocalMux I__20630 (
            .O(N__88044),
            .I(N__88041));
    Span4Mux_h I__20629 (
            .O(N__88041),
            .I(N__88038));
    Odrv4 I__20628 (
            .O(N__88038),
            .I(\quad_counter1.n7_adj_4445 ));
    InMux I__20627 (
            .O(N__88035),
            .I(N__88031));
    InMux I__20626 (
            .O(N__88034),
            .I(N__88028));
    LocalMux I__20625 (
            .O(N__88031),
            .I(N__88022));
    LocalMux I__20624 (
            .O(N__88028),
            .I(N__88022));
    InMux I__20623 (
            .O(N__88027),
            .I(N__88019));
    Span4Mux_h I__20622 (
            .O(N__88022),
            .I(N__88016));
    LocalMux I__20621 (
            .O(N__88019),
            .I(N__88013));
    Odrv4 I__20620 (
            .O(N__88016),
            .I(\quad_counter1.n2607 ));
    Odrv4 I__20619 (
            .O(N__88013),
            .I(\quad_counter1.n2607 ));
    InMux I__20618 (
            .O(N__88008),
            .I(\quad_counter1.n30533 ));
    InMux I__20617 (
            .O(N__88005),
            .I(N__88001));
    InMux I__20616 (
            .O(N__88004),
            .I(N__87998));
    LocalMux I__20615 (
            .O(N__88001),
            .I(N__87992));
    LocalMux I__20614 (
            .O(N__87998),
            .I(N__87992));
    InMux I__20613 (
            .O(N__87997),
            .I(N__87989));
    Span4Mux_h I__20612 (
            .O(N__87992),
            .I(N__87986));
    LocalMux I__20611 (
            .O(N__87989),
            .I(N__87983));
    Odrv4 I__20610 (
            .O(N__87986),
            .I(\quad_counter1.n2507 ));
    Odrv4 I__20609 (
            .O(N__87983),
            .I(\quad_counter1.n2507 ));
    InMux I__20608 (
            .O(N__87978),
            .I(\quad_counter1.n30534 ));
    InMux I__20607 (
            .O(N__87975),
            .I(N__87971));
    InMux I__20606 (
            .O(N__87974),
            .I(N__87968));
    LocalMux I__20605 (
            .O(N__87971),
            .I(N__87962));
    LocalMux I__20604 (
            .O(N__87968),
            .I(N__87962));
    InMux I__20603 (
            .O(N__87967),
            .I(N__87959));
    Span4Mux_v I__20602 (
            .O(N__87962),
            .I(N__87956));
    LocalMux I__20601 (
            .O(N__87959),
            .I(N__87953));
    Odrv4 I__20600 (
            .O(N__87956),
            .I(\quad_counter1.n2606 ));
    Odrv4 I__20599 (
            .O(N__87953),
            .I(\quad_counter1.n2606 ));
    CascadeMux I__20598 (
            .O(N__87948),
            .I(N__87941));
    CascadeMux I__20597 (
            .O(N__87947),
            .I(N__87938));
    CascadeMux I__20596 (
            .O(N__87946),
            .I(N__87932));
    CascadeMux I__20595 (
            .O(N__87945),
            .I(N__87929));
    CascadeMux I__20594 (
            .O(N__87944),
            .I(N__87926));
    InMux I__20593 (
            .O(N__87941),
            .I(N__87921));
    InMux I__20592 (
            .O(N__87938),
            .I(N__87921));
    CascadeMux I__20591 (
            .O(N__87937),
            .I(N__87918));
    CascadeMux I__20590 (
            .O(N__87936),
            .I(N__87915));
    CascadeMux I__20589 (
            .O(N__87935),
            .I(N__87912));
    InMux I__20588 (
            .O(N__87932),
            .I(N__87904));
    InMux I__20587 (
            .O(N__87929),
            .I(N__87904));
    InMux I__20586 (
            .O(N__87926),
            .I(N__87904));
    LocalMux I__20585 (
            .O(N__87921),
            .I(N__87901));
    InMux I__20584 (
            .O(N__87918),
            .I(N__87892));
    InMux I__20583 (
            .O(N__87915),
            .I(N__87892));
    InMux I__20582 (
            .O(N__87912),
            .I(N__87892));
    InMux I__20581 (
            .O(N__87911),
            .I(N__87892));
    LocalMux I__20580 (
            .O(N__87904),
            .I(N__87885));
    Span4Mux_v I__20579 (
            .O(N__87901),
            .I(N__87885));
    LocalMux I__20578 (
            .O(N__87892),
            .I(N__87885));
    Odrv4 I__20577 (
            .O(N__87885),
            .I(\quad_counter1.n2540 ));
    CascadeMux I__20576 (
            .O(N__87882),
            .I(N__87874));
    CascadeMux I__20575 (
            .O(N__87881),
            .I(N__87871));
    CascadeMux I__20574 (
            .O(N__87880),
            .I(N__87868));
    CascadeMux I__20573 (
            .O(N__87879),
            .I(N__87865));
    CascadeMux I__20572 (
            .O(N__87878),
            .I(N__87862));
    CascadeMux I__20571 (
            .O(N__87877),
            .I(N__87859));
    InMux I__20570 (
            .O(N__87874),
            .I(N__87854));
    InMux I__20569 (
            .O(N__87871),
            .I(N__87854));
    InMux I__20568 (
            .O(N__87868),
            .I(N__87845));
    InMux I__20567 (
            .O(N__87865),
            .I(N__87845));
    InMux I__20566 (
            .O(N__87862),
            .I(N__87845));
    InMux I__20565 (
            .O(N__87859),
            .I(N__87845));
    LocalMux I__20564 (
            .O(N__87854),
            .I(\quad_counter1.n36133 ));
    LocalMux I__20563 (
            .O(N__87845),
            .I(\quad_counter1.n36133 ));
    InMux I__20562 (
            .O(N__87840),
            .I(bfn_23_9_0_));
    InMux I__20561 (
            .O(N__87837),
            .I(\quad_counter1.n30499 ));
    InMux I__20560 (
            .O(N__87834),
            .I(N__87829));
    InMux I__20559 (
            .O(N__87833),
            .I(N__87826));
    InMux I__20558 (
            .O(N__87832),
            .I(N__87823));
    LocalMux I__20557 (
            .O(N__87829),
            .I(N__87820));
    LocalMux I__20556 (
            .O(N__87826),
            .I(N__87813));
    LocalMux I__20555 (
            .O(N__87823),
            .I(N__87813));
    Span4Mux_v I__20554 (
            .O(N__87820),
            .I(N__87813));
    Odrv4 I__20553 (
            .O(N__87813),
            .I(\quad_counter1.n2417 ));
    InMux I__20552 (
            .O(N__87810),
            .I(\quad_counter1.n30500 ));
    InMux I__20551 (
            .O(N__87807),
            .I(N__87802));
    InMux I__20550 (
            .O(N__87806),
            .I(N__87799));
    InMux I__20549 (
            .O(N__87805),
            .I(N__87796));
    LocalMux I__20548 (
            .O(N__87802),
            .I(N__87793));
    LocalMux I__20547 (
            .O(N__87799),
            .I(N__87788));
    LocalMux I__20546 (
            .O(N__87796),
            .I(N__87788));
    Span4Mux_h I__20545 (
            .O(N__87793),
            .I(N__87785));
    Odrv4 I__20544 (
            .O(N__87788),
            .I(\quad_counter1.n2416 ));
    Odrv4 I__20543 (
            .O(N__87785),
            .I(\quad_counter1.n2416 ));
    InMux I__20542 (
            .O(N__87780),
            .I(\quad_counter1.n30501 ));
    InMux I__20541 (
            .O(N__87777),
            .I(N__87772));
    InMux I__20540 (
            .O(N__87776),
            .I(N__87769));
    InMux I__20539 (
            .O(N__87775),
            .I(N__87766));
    LocalMux I__20538 (
            .O(N__87772),
            .I(N__87763));
    LocalMux I__20537 (
            .O(N__87769),
            .I(N__87758));
    LocalMux I__20536 (
            .O(N__87766),
            .I(N__87758));
    Span4Mux_h I__20535 (
            .O(N__87763),
            .I(N__87755));
    Odrv4 I__20534 (
            .O(N__87758),
            .I(\quad_counter1.n2415 ));
    Odrv4 I__20533 (
            .O(N__87755),
            .I(\quad_counter1.n2415 ));
    InMux I__20532 (
            .O(N__87750),
            .I(\quad_counter1.n30502 ));
    InMux I__20531 (
            .O(N__87747),
            .I(N__87742));
    InMux I__20530 (
            .O(N__87746),
            .I(N__87739));
    InMux I__20529 (
            .O(N__87745),
            .I(N__87736));
    LocalMux I__20528 (
            .O(N__87742),
            .I(N__87733));
    LocalMux I__20527 (
            .O(N__87739),
            .I(N__87728));
    LocalMux I__20526 (
            .O(N__87736),
            .I(N__87728));
    Span4Mux_h I__20525 (
            .O(N__87733),
            .I(N__87725));
    Odrv4 I__20524 (
            .O(N__87728),
            .I(\quad_counter1.n2414 ));
    Odrv4 I__20523 (
            .O(N__87725),
            .I(\quad_counter1.n2414 ));
    InMux I__20522 (
            .O(N__87720),
            .I(\quad_counter1.n30503 ));
    InMux I__20521 (
            .O(N__87717),
            .I(N__87713));
    InMux I__20520 (
            .O(N__87716),
            .I(N__87710));
    LocalMux I__20519 (
            .O(N__87713),
            .I(N__87705));
    LocalMux I__20518 (
            .O(N__87710),
            .I(N__87705));
    Span4Mux_h I__20517 (
            .O(N__87705),
            .I(N__87701));
    InMux I__20516 (
            .O(N__87704),
            .I(N__87698));
    Odrv4 I__20515 (
            .O(N__87701),
            .I(\quad_counter1.n2515 ));
    LocalMux I__20514 (
            .O(N__87698),
            .I(\quad_counter1.n2515 ));
    InMux I__20513 (
            .O(N__87693),
            .I(N__87689));
    InMux I__20512 (
            .O(N__87692),
            .I(N__87686));
    LocalMux I__20511 (
            .O(N__87689),
            .I(N__87681));
    LocalMux I__20510 (
            .O(N__87686),
            .I(N__87681));
    Span4Mux_h I__20509 (
            .O(N__87681),
            .I(N__87677));
    InMux I__20508 (
            .O(N__87680),
            .I(N__87674));
    Odrv4 I__20507 (
            .O(N__87677),
            .I(\quad_counter1.n2614 ));
    LocalMux I__20506 (
            .O(N__87674),
            .I(\quad_counter1.n2614 ));
    InMux I__20505 (
            .O(N__87669),
            .I(\quad_counter1.n30526 ));
    InMux I__20504 (
            .O(N__87666),
            .I(N__87662));
    InMux I__20503 (
            .O(N__87665),
            .I(N__87659));
    LocalMux I__20502 (
            .O(N__87662),
            .I(N__87654));
    LocalMux I__20501 (
            .O(N__87659),
            .I(N__87654));
    Span4Mux_h I__20500 (
            .O(N__87654),
            .I(N__87650));
    InMux I__20499 (
            .O(N__87653),
            .I(N__87647));
    Odrv4 I__20498 (
            .O(N__87650),
            .I(\quad_counter1.n2514 ));
    LocalMux I__20497 (
            .O(N__87647),
            .I(\quad_counter1.n2514 ));
    InMux I__20496 (
            .O(N__87642),
            .I(N__87638));
    InMux I__20495 (
            .O(N__87641),
            .I(N__87635));
    LocalMux I__20494 (
            .O(N__87638),
            .I(N__87630));
    LocalMux I__20493 (
            .O(N__87635),
            .I(N__87630));
    Span4Mux_v I__20492 (
            .O(N__87630),
            .I(N__87626));
    InMux I__20491 (
            .O(N__87629),
            .I(N__87623));
    Odrv4 I__20490 (
            .O(N__87626),
            .I(\quad_counter1.n2613 ));
    LocalMux I__20489 (
            .O(N__87623),
            .I(\quad_counter1.n2613 ));
    InMux I__20488 (
            .O(N__87618),
            .I(\quad_counter1.n30527 ));
    InMux I__20487 (
            .O(N__87615),
            .I(N__87611));
    InMux I__20486 (
            .O(N__87614),
            .I(N__87608));
    LocalMux I__20485 (
            .O(N__87611),
            .I(N__87603));
    LocalMux I__20484 (
            .O(N__87608),
            .I(N__87603));
    Span4Mux_h I__20483 (
            .O(N__87603),
            .I(N__87599));
    InMux I__20482 (
            .O(N__87602),
            .I(N__87596));
    Odrv4 I__20481 (
            .O(N__87599),
            .I(\quad_counter1.n2513 ));
    LocalMux I__20480 (
            .O(N__87596),
            .I(\quad_counter1.n2513 ));
    InMux I__20479 (
            .O(N__87591),
            .I(N__87587));
    InMux I__20478 (
            .O(N__87590),
            .I(N__87584));
    LocalMux I__20477 (
            .O(N__87587),
            .I(N__87579));
    LocalMux I__20476 (
            .O(N__87584),
            .I(N__87579));
    Span4Mux_h I__20475 (
            .O(N__87579),
            .I(N__87575));
    InMux I__20474 (
            .O(N__87578),
            .I(N__87572));
    Odrv4 I__20473 (
            .O(N__87575),
            .I(\quad_counter1.n2612 ));
    LocalMux I__20472 (
            .O(N__87572),
            .I(\quad_counter1.n2612 ));
    InMux I__20471 (
            .O(N__87567),
            .I(\quad_counter1.n30528 ));
    InMux I__20470 (
            .O(N__87564),
            .I(N__87560));
    InMux I__20469 (
            .O(N__87563),
            .I(N__87557));
    LocalMux I__20468 (
            .O(N__87560),
            .I(N__87552));
    LocalMux I__20467 (
            .O(N__87557),
            .I(N__87552));
    Span4Mux_h I__20466 (
            .O(N__87552),
            .I(N__87548));
    InMux I__20465 (
            .O(N__87551),
            .I(N__87545));
    Odrv4 I__20464 (
            .O(N__87548),
            .I(\quad_counter1.n2512 ));
    LocalMux I__20463 (
            .O(N__87545),
            .I(\quad_counter1.n2512 ));
    InMux I__20462 (
            .O(N__87540),
            .I(N__87536));
    InMux I__20461 (
            .O(N__87539),
            .I(N__87533));
    LocalMux I__20460 (
            .O(N__87536),
            .I(N__87527));
    LocalMux I__20459 (
            .O(N__87533),
            .I(N__87527));
    InMux I__20458 (
            .O(N__87532),
            .I(N__87524));
    Span4Mux_h I__20457 (
            .O(N__87527),
            .I(N__87521));
    LocalMux I__20456 (
            .O(N__87524),
            .I(N__87518));
    Odrv4 I__20455 (
            .O(N__87521),
            .I(\quad_counter1.n2611 ));
    Odrv4 I__20454 (
            .O(N__87518),
            .I(\quad_counter1.n2611 ));
    InMux I__20453 (
            .O(N__87513),
            .I(bfn_23_8_0_));
    InMux I__20452 (
            .O(N__87510),
            .I(N__87505));
    InMux I__20451 (
            .O(N__87509),
            .I(N__87502));
    CascadeMux I__20450 (
            .O(N__87508),
            .I(N__87499));
    LocalMux I__20449 (
            .O(N__87505),
            .I(N__87494));
    LocalMux I__20448 (
            .O(N__87502),
            .I(N__87494));
    InMux I__20447 (
            .O(N__87499),
            .I(N__87491));
    Span4Mux_h I__20446 (
            .O(N__87494),
            .I(N__87488));
    LocalMux I__20445 (
            .O(N__87491),
            .I(N__87485));
    Odrv4 I__20444 (
            .O(N__87488),
            .I(\quad_counter1.n2511 ));
    Odrv4 I__20443 (
            .O(N__87485),
            .I(\quad_counter1.n2511 ));
    InMux I__20442 (
            .O(N__87480),
            .I(N__87476));
    InMux I__20441 (
            .O(N__87479),
            .I(N__87473));
    LocalMux I__20440 (
            .O(N__87476),
            .I(N__87467));
    LocalMux I__20439 (
            .O(N__87473),
            .I(N__87467));
    InMux I__20438 (
            .O(N__87472),
            .I(N__87464));
    Span4Mux_h I__20437 (
            .O(N__87467),
            .I(N__87461));
    LocalMux I__20436 (
            .O(N__87464),
            .I(N__87458));
    Odrv4 I__20435 (
            .O(N__87461),
            .I(\quad_counter1.n2610 ));
    Odrv4 I__20434 (
            .O(N__87458),
            .I(\quad_counter1.n2610 ));
    InMux I__20433 (
            .O(N__87453),
            .I(\quad_counter1.n30530 ));
    InMux I__20432 (
            .O(N__87450),
            .I(N__87446));
    InMux I__20431 (
            .O(N__87449),
            .I(N__87443));
    LocalMux I__20430 (
            .O(N__87446),
            .I(N__87437));
    LocalMux I__20429 (
            .O(N__87443),
            .I(N__87437));
    InMux I__20428 (
            .O(N__87442),
            .I(N__87434));
    Span4Mux_h I__20427 (
            .O(N__87437),
            .I(N__87431));
    LocalMux I__20426 (
            .O(N__87434),
            .I(N__87428));
    Odrv4 I__20425 (
            .O(N__87431),
            .I(\quad_counter1.n2510 ));
    Odrv4 I__20424 (
            .O(N__87428),
            .I(\quad_counter1.n2510 ));
    InMux I__20423 (
            .O(N__87423),
            .I(N__87419));
    InMux I__20422 (
            .O(N__87422),
            .I(N__87416));
    LocalMux I__20421 (
            .O(N__87419),
            .I(N__87410));
    LocalMux I__20420 (
            .O(N__87416),
            .I(N__87410));
    InMux I__20419 (
            .O(N__87415),
            .I(N__87407));
    Span4Mux_v I__20418 (
            .O(N__87410),
            .I(N__87404));
    LocalMux I__20417 (
            .O(N__87407),
            .I(N__87401));
    Odrv4 I__20416 (
            .O(N__87404),
            .I(\quad_counter1.n2609 ));
    Odrv4 I__20415 (
            .O(N__87401),
            .I(\quad_counter1.n2609 ));
    InMux I__20414 (
            .O(N__87396),
            .I(\quad_counter1.n30531 ));
    InMux I__20413 (
            .O(N__87393),
            .I(N__87389));
    InMux I__20412 (
            .O(N__87392),
            .I(N__87386));
    LocalMux I__20411 (
            .O(N__87389),
            .I(N__87382));
    LocalMux I__20410 (
            .O(N__87386),
            .I(N__87379));
    InMux I__20409 (
            .O(N__87385),
            .I(N__87376));
    Span4Mux_v I__20408 (
            .O(N__87382),
            .I(N__87371));
    Span4Mux_v I__20407 (
            .O(N__87379),
            .I(N__87371));
    LocalMux I__20406 (
            .O(N__87376),
            .I(N__87368));
    Odrv4 I__20405 (
            .O(N__87371),
            .I(\quad_counter1.n2509 ));
    Odrv4 I__20404 (
            .O(N__87368),
            .I(\quad_counter1.n2509 ));
    InMux I__20403 (
            .O(N__87363),
            .I(N__87359));
    InMux I__20402 (
            .O(N__87362),
            .I(N__87356));
    LocalMux I__20401 (
            .O(N__87359),
            .I(N__87350));
    LocalMux I__20400 (
            .O(N__87356),
            .I(N__87350));
    InMux I__20399 (
            .O(N__87355),
            .I(N__87347));
    Span4Mux_v I__20398 (
            .O(N__87350),
            .I(N__87344));
    LocalMux I__20397 (
            .O(N__87347),
            .I(N__87341));
    Odrv4 I__20396 (
            .O(N__87344),
            .I(\quad_counter1.n2608 ));
    Odrv4 I__20395 (
            .O(N__87341),
            .I(\quad_counter1.n2608 ));
    InMux I__20394 (
            .O(N__87336),
            .I(\quad_counter1.n30532 ));
    InMux I__20393 (
            .O(N__87333),
            .I(N__87329));
    InMux I__20392 (
            .O(N__87332),
            .I(N__87326));
    LocalMux I__20391 (
            .O(N__87329),
            .I(N__87320));
    LocalMux I__20390 (
            .O(N__87326),
            .I(N__87320));
    InMux I__20389 (
            .O(N__87325),
            .I(N__87317));
    Span4Mux_v I__20388 (
            .O(N__87320),
            .I(N__87314));
    LocalMux I__20387 (
            .O(N__87317),
            .I(N__87311));
    Odrv4 I__20386 (
            .O(N__87314),
            .I(\quad_counter1.n2508 ));
    Odrv4 I__20385 (
            .O(N__87311),
            .I(\quad_counter1.n2508 ));
    CascadeMux I__20384 (
            .O(N__87306),
            .I(N__87291));
    InMux I__20383 (
            .O(N__87305),
            .I(N__87287));
    CascadeMux I__20382 (
            .O(N__87304),
            .I(N__87284));
    CascadeMux I__20381 (
            .O(N__87303),
            .I(N__87281));
    InMux I__20380 (
            .O(N__87302),
            .I(N__87278));
    CascadeMux I__20379 (
            .O(N__87301),
            .I(N__87275));
    CascadeMux I__20378 (
            .O(N__87300),
            .I(N__87271));
    CascadeMux I__20377 (
            .O(N__87299),
            .I(N__87267));
    InMux I__20376 (
            .O(N__87298),
            .I(N__87264));
    InMux I__20375 (
            .O(N__87297),
            .I(N__87260));
    InMux I__20374 (
            .O(N__87296),
            .I(N__87256));
    InMux I__20373 (
            .O(N__87295),
            .I(N__87253));
    InMux I__20372 (
            .O(N__87294),
            .I(N__87248));
    InMux I__20371 (
            .O(N__87291),
            .I(N__87248));
    InMux I__20370 (
            .O(N__87290),
            .I(N__87245));
    LocalMux I__20369 (
            .O(N__87287),
            .I(N__87242));
    InMux I__20368 (
            .O(N__87284),
            .I(N__87234));
    InMux I__20367 (
            .O(N__87281),
            .I(N__87234));
    LocalMux I__20366 (
            .O(N__87278),
            .I(N__87231));
    InMux I__20365 (
            .O(N__87275),
            .I(N__87228));
    InMux I__20364 (
            .O(N__87274),
            .I(N__87225));
    InMux I__20363 (
            .O(N__87271),
            .I(N__87222));
    InMux I__20362 (
            .O(N__87270),
            .I(N__87215));
    InMux I__20361 (
            .O(N__87267),
            .I(N__87215));
    LocalMux I__20360 (
            .O(N__87264),
            .I(N__87212));
    InMux I__20359 (
            .O(N__87263),
            .I(N__87209));
    LocalMux I__20358 (
            .O(N__87260),
            .I(N__87206));
    InMux I__20357 (
            .O(N__87259),
            .I(N__87203));
    LocalMux I__20356 (
            .O(N__87256),
            .I(N__87200));
    LocalMux I__20355 (
            .O(N__87253),
            .I(N__87193));
    LocalMux I__20354 (
            .O(N__87248),
            .I(N__87193));
    LocalMux I__20353 (
            .O(N__87245),
            .I(N__87188));
    Span4Mux_v I__20352 (
            .O(N__87242),
            .I(N__87188));
    InMux I__20351 (
            .O(N__87241),
            .I(N__87184));
    InMux I__20350 (
            .O(N__87240),
            .I(N__87179));
    InMux I__20349 (
            .O(N__87239),
            .I(N__87179));
    LocalMux I__20348 (
            .O(N__87234),
            .I(N__87176));
    Span4Mux_v I__20347 (
            .O(N__87231),
            .I(N__87173));
    LocalMux I__20346 (
            .O(N__87228),
            .I(N__87170));
    LocalMux I__20345 (
            .O(N__87225),
            .I(N__87163));
    LocalMux I__20344 (
            .O(N__87222),
            .I(N__87163));
    InMux I__20343 (
            .O(N__87221),
            .I(N__87160));
    InMux I__20342 (
            .O(N__87220),
            .I(N__87157));
    LocalMux I__20341 (
            .O(N__87215),
            .I(N__87154));
    Span4Mux_h I__20340 (
            .O(N__87212),
            .I(N__87149));
    LocalMux I__20339 (
            .O(N__87209),
            .I(N__87149));
    Span4Mux_h I__20338 (
            .O(N__87206),
            .I(N__87143));
    LocalMux I__20337 (
            .O(N__87203),
            .I(N__87143));
    Span4Mux_v I__20336 (
            .O(N__87200),
            .I(N__87140));
    CascadeMux I__20335 (
            .O(N__87199),
            .I(N__87136));
    InMux I__20334 (
            .O(N__87198),
            .I(N__87133));
    Span4Mux_v I__20333 (
            .O(N__87193),
            .I(N__87130));
    Span4Mux_v I__20332 (
            .O(N__87188),
            .I(N__87127));
    InMux I__20331 (
            .O(N__87187),
            .I(N__87123));
    LocalMux I__20330 (
            .O(N__87184),
            .I(N__87118));
    LocalMux I__20329 (
            .O(N__87179),
            .I(N__87118));
    Span4Mux_v I__20328 (
            .O(N__87176),
            .I(N__87115));
    Span4Mux_h I__20327 (
            .O(N__87173),
            .I(N__87112));
    Span4Mux_v I__20326 (
            .O(N__87170),
            .I(N__87109));
    CascadeMux I__20325 (
            .O(N__87169),
            .I(N__87106));
    CascadeMux I__20324 (
            .O(N__87168),
            .I(N__87102));
    Span4Mux_v I__20323 (
            .O(N__87163),
            .I(N__87099));
    LocalMux I__20322 (
            .O(N__87160),
            .I(N__87094));
    LocalMux I__20321 (
            .O(N__87157),
            .I(N__87094));
    Span4Mux_h I__20320 (
            .O(N__87154),
            .I(N__87091));
    Span4Mux_h I__20319 (
            .O(N__87149),
            .I(N__87088));
    InMux I__20318 (
            .O(N__87148),
            .I(N__87085));
    Span4Mux_v I__20317 (
            .O(N__87143),
            .I(N__87080));
    Span4Mux_v I__20316 (
            .O(N__87140),
            .I(N__87080));
    InMux I__20315 (
            .O(N__87139),
            .I(N__87077));
    InMux I__20314 (
            .O(N__87136),
            .I(N__87074));
    LocalMux I__20313 (
            .O(N__87133),
            .I(N__87071));
    Span4Mux_h I__20312 (
            .O(N__87130),
            .I(N__87066));
    Span4Mux_h I__20311 (
            .O(N__87127),
            .I(N__87066));
    InMux I__20310 (
            .O(N__87126),
            .I(N__87063));
    LocalMux I__20309 (
            .O(N__87123),
            .I(N__87060));
    Span4Mux_v I__20308 (
            .O(N__87118),
            .I(N__87057));
    Span4Mux_h I__20307 (
            .O(N__87115),
            .I(N__87054));
    Span4Mux_h I__20306 (
            .O(N__87112),
            .I(N__87051));
    Span4Mux_h I__20305 (
            .O(N__87109),
            .I(N__87048));
    InMux I__20304 (
            .O(N__87106),
            .I(N__87041));
    InMux I__20303 (
            .O(N__87105),
            .I(N__87041));
    InMux I__20302 (
            .O(N__87102),
            .I(N__87041));
    Sp12to4 I__20301 (
            .O(N__87099),
            .I(N__87036));
    Span12Mux_v I__20300 (
            .O(N__87094),
            .I(N__87036));
    Span4Mux_h I__20299 (
            .O(N__87091),
            .I(N__87033));
    Sp12to4 I__20298 (
            .O(N__87088),
            .I(N__87028));
    LocalMux I__20297 (
            .O(N__87085),
            .I(N__87028));
    Span4Mux_v I__20296 (
            .O(N__87080),
            .I(N__87025));
    LocalMux I__20295 (
            .O(N__87077),
            .I(N__87018));
    LocalMux I__20294 (
            .O(N__87074),
            .I(N__87018));
    Sp12to4 I__20293 (
            .O(N__87071),
            .I(N__87018));
    Span4Mux_v I__20292 (
            .O(N__87066),
            .I(N__87015));
    LocalMux I__20291 (
            .O(N__87063),
            .I(N__87012));
    Span4Mux_h I__20290 (
            .O(N__87060),
            .I(N__87007));
    Span4Mux_h I__20289 (
            .O(N__87057),
            .I(N__87007));
    Sp12to4 I__20288 (
            .O(N__87054),
            .I(N__87004));
    Span4Mux_h I__20287 (
            .O(N__87051),
            .I(N__86999));
    Span4Mux_h I__20286 (
            .O(N__87048),
            .I(N__86999));
    LocalMux I__20285 (
            .O(N__87041),
            .I(N__86996));
    Span12Mux_v I__20284 (
            .O(N__87036),
            .I(N__86993));
    Sp12to4 I__20283 (
            .O(N__87033),
            .I(N__86988));
    Span12Mux_v I__20282 (
            .O(N__87028),
            .I(N__86988));
    Sp12to4 I__20281 (
            .O(N__87025),
            .I(N__86981));
    Span12Mux_v I__20280 (
            .O(N__87018),
            .I(N__86981));
    Sp12to4 I__20279 (
            .O(N__87015),
            .I(N__86981));
    Sp12to4 I__20278 (
            .O(N__87012),
            .I(N__86970));
    Sp12to4 I__20277 (
            .O(N__87007),
            .I(N__86970));
    Span12Mux_s9_h I__20276 (
            .O(N__87004),
            .I(N__86970));
    Sp12to4 I__20275 (
            .O(N__86999),
            .I(N__86970));
    Span12Mux_h I__20274 (
            .O(N__86996),
            .I(N__86970));
    Span12Mux_h I__20273 (
            .O(N__86993),
            .I(N__86965));
    Span12Mux_v I__20272 (
            .O(N__86988),
            .I(N__86965));
    Span12Mux_h I__20271 (
            .O(N__86981),
            .I(N__86960));
    Span12Mux_v I__20270 (
            .O(N__86970),
            .I(N__86960));
    Odrv12 I__20269 (
            .O(N__86965),
            .I(\c0.n9_adj_4493 ));
    Odrv12 I__20268 (
            .O(N__86960),
            .I(\c0.n9_adj_4493 ));
    InMux I__20267 (
            .O(N__86955),
            .I(N__86951));
    InMux I__20266 (
            .O(N__86954),
            .I(N__86948));
    LocalMux I__20265 (
            .O(N__86951),
            .I(N__86941));
    LocalMux I__20264 (
            .O(N__86948),
            .I(N__86941));
    InMux I__20263 (
            .O(N__86947),
            .I(N__86938));
    InMux I__20262 (
            .O(N__86946),
            .I(N__86935));
    Span4Mux_h I__20261 (
            .O(N__86941),
            .I(N__86930));
    LocalMux I__20260 (
            .O(N__86938),
            .I(N__86930));
    LocalMux I__20259 (
            .O(N__86935),
            .I(\quad_counter1.millisecond_counter_17 ));
    Odrv4 I__20258 (
            .O(N__86930),
            .I(\quad_counter1.millisecond_counter_17 ));
    CascadeMux I__20257 (
            .O(N__86925),
            .I(\quad_counter1.n28271_cascade_ ));
    CascadeMux I__20256 (
            .O(N__86922),
            .I(\quad_counter1.n10_adj_4423_cascade_ ));
    InMux I__20255 (
            .O(N__86919),
            .I(N__86916));
    LocalMux I__20254 (
            .O(N__86916),
            .I(\quad_counter1.n11 ));
    InMux I__20253 (
            .O(N__86913),
            .I(N__86909));
    InMux I__20252 (
            .O(N__86912),
            .I(N__86906));
    LocalMux I__20251 (
            .O(N__86909),
            .I(N__86900));
    LocalMux I__20250 (
            .O(N__86906),
            .I(N__86900));
    InMux I__20249 (
            .O(N__86905),
            .I(N__86896));
    Span4Mux_v I__20248 (
            .O(N__86900),
            .I(N__86893));
    InMux I__20247 (
            .O(N__86899),
            .I(N__86890));
    LocalMux I__20246 (
            .O(N__86896),
            .I(\quad_counter1.millisecond_counter_18 ));
    Odrv4 I__20245 (
            .O(N__86893),
            .I(\quad_counter1.millisecond_counter_18 ));
    LocalMux I__20244 (
            .O(N__86890),
            .I(\quad_counter1.millisecond_counter_18 ));
    InMux I__20243 (
            .O(N__86883),
            .I(N__86879));
    InMux I__20242 (
            .O(N__86882),
            .I(N__86876));
    LocalMux I__20241 (
            .O(N__86879),
            .I(N__86873));
    LocalMux I__20240 (
            .O(N__86876),
            .I(N__86870));
    Span4Mux_h I__20239 (
            .O(N__86873),
            .I(N__86866));
    Span4Mux_h I__20238 (
            .O(N__86870),
            .I(N__86863));
    InMux I__20237 (
            .O(N__86869),
            .I(N__86860));
    Odrv4 I__20236 (
            .O(N__86866),
            .I(\quad_counter1.n2619 ));
    Odrv4 I__20235 (
            .O(N__86863),
            .I(\quad_counter1.n2619 ));
    LocalMux I__20234 (
            .O(N__86860),
            .I(\quad_counter1.n2619 ));
    InMux I__20233 (
            .O(N__86853),
            .I(bfn_23_7_0_));
    InMux I__20232 (
            .O(N__86850),
            .I(N__86846));
    InMux I__20231 (
            .O(N__86849),
            .I(N__86843));
    LocalMux I__20230 (
            .O(N__86846),
            .I(N__86838));
    LocalMux I__20229 (
            .O(N__86843),
            .I(N__86838));
    Span4Mux_h I__20228 (
            .O(N__86838),
            .I(N__86834));
    InMux I__20227 (
            .O(N__86837),
            .I(N__86831));
    Odrv4 I__20226 (
            .O(N__86834),
            .I(\quad_counter1.n2519 ));
    LocalMux I__20225 (
            .O(N__86831),
            .I(\quad_counter1.n2519 ));
    InMux I__20224 (
            .O(N__86826),
            .I(N__86822));
    InMux I__20223 (
            .O(N__86825),
            .I(N__86819));
    LocalMux I__20222 (
            .O(N__86822),
            .I(N__86814));
    LocalMux I__20221 (
            .O(N__86819),
            .I(N__86814));
    Span4Mux_h I__20220 (
            .O(N__86814),
            .I(N__86810));
    InMux I__20219 (
            .O(N__86813),
            .I(N__86807));
    Odrv4 I__20218 (
            .O(N__86810),
            .I(\quad_counter1.n2618 ));
    LocalMux I__20217 (
            .O(N__86807),
            .I(\quad_counter1.n2618 ));
    InMux I__20216 (
            .O(N__86802),
            .I(\quad_counter1.n30522 ));
    InMux I__20215 (
            .O(N__86799),
            .I(N__86795));
    InMux I__20214 (
            .O(N__86798),
            .I(N__86792));
    LocalMux I__20213 (
            .O(N__86795),
            .I(N__86787));
    LocalMux I__20212 (
            .O(N__86792),
            .I(N__86787));
    Span4Mux_h I__20211 (
            .O(N__86787),
            .I(N__86783));
    InMux I__20210 (
            .O(N__86786),
            .I(N__86780));
    Odrv4 I__20209 (
            .O(N__86783),
            .I(\quad_counter1.n2518 ));
    LocalMux I__20208 (
            .O(N__86780),
            .I(\quad_counter1.n2518 ));
    InMux I__20207 (
            .O(N__86775),
            .I(N__86771));
    InMux I__20206 (
            .O(N__86774),
            .I(N__86768));
    LocalMux I__20205 (
            .O(N__86771),
            .I(N__86763));
    LocalMux I__20204 (
            .O(N__86768),
            .I(N__86763));
    Span4Mux_v I__20203 (
            .O(N__86763),
            .I(N__86759));
    InMux I__20202 (
            .O(N__86762),
            .I(N__86756));
    Odrv4 I__20201 (
            .O(N__86759),
            .I(\quad_counter1.n2617 ));
    LocalMux I__20200 (
            .O(N__86756),
            .I(\quad_counter1.n2617 ));
    InMux I__20199 (
            .O(N__86751),
            .I(\quad_counter1.n30523 ));
    InMux I__20198 (
            .O(N__86748),
            .I(N__86744));
    InMux I__20197 (
            .O(N__86747),
            .I(N__86741));
    LocalMux I__20196 (
            .O(N__86744),
            .I(N__86736));
    LocalMux I__20195 (
            .O(N__86741),
            .I(N__86736));
    Span4Mux_v I__20194 (
            .O(N__86736),
            .I(N__86732));
    InMux I__20193 (
            .O(N__86735),
            .I(N__86729));
    Odrv4 I__20192 (
            .O(N__86732),
            .I(\quad_counter1.n2517 ));
    LocalMux I__20191 (
            .O(N__86729),
            .I(\quad_counter1.n2517 ));
    InMux I__20190 (
            .O(N__86724),
            .I(N__86720));
    InMux I__20189 (
            .O(N__86723),
            .I(N__86717));
    LocalMux I__20188 (
            .O(N__86720),
            .I(N__86712));
    LocalMux I__20187 (
            .O(N__86717),
            .I(N__86712));
    Span4Mux_v I__20186 (
            .O(N__86712),
            .I(N__86708));
    InMux I__20185 (
            .O(N__86711),
            .I(N__86705));
    Odrv4 I__20184 (
            .O(N__86708),
            .I(\quad_counter1.n2616 ));
    LocalMux I__20183 (
            .O(N__86705),
            .I(\quad_counter1.n2616 ));
    InMux I__20182 (
            .O(N__86700),
            .I(\quad_counter1.n30524 ));
    InMux I__20181 (
            .O(N__86697),
            .I(N__86693));
    InMux I__20180 (
            .O(N__86696),
            .I(N__86690));
    LocalMux I__20179 (
            .O(N__86693),
            .I(N__86685));
    LocalMux I__20178 (
            .O(N__86690),
            .I(N__86685));
    Span4Mux_v I__20177 (
            .O(N__86685),
            .I(N__86681));
    InMux I__20176 (
            .O(N__86684),
            .I(N__86678));
    Odrv4 I__20175 (
            .O(N__86681),
            .I(\quad_counter1.n2516 ));
    LocalMux I__20174 (
            .O(N__86678),
            .I(\quad_counter1.n2516 ));
    InMux I__20173 (
            .O(N__86673),
            .I(N__86669));
    InMux I__20172 (
            .O(N__86672),
            .I(N__86666));
    LocalMux I__20171 (
            .O(N__86669),
            .I(N__86661));
    LocalMux I__20170 (
            .O(N__86666),
            .I(N__86661));
    Span4Mux_h I__20169 (
            .O(N__86661),
            .I(N__86657));
    InMux I__20168 (
            .O(N__86660),
            .I(N__86654));
    Odrv4 I__20167 (
            .O(N__86657),
            .I(\quad_counter1.n2615 ));
    LocalMux I__20166 (
            .O(N__86654),
            .I(\quad_counter1.n2615 ));
    InMux I__20165 (
            .O(N__86649),
            .I(\quad_counter1.n30525 ));
    InMux I__20164 (
            .O(N__86646),
            .I(N__86642));
    InMux I__20163 (
            .O(N__86645),
            .I(N__86639));
    LocalMux I__20162 (
            .O(N__86642),
            .I(N__86631));
    LocalMux I__20161 (
            .O(N__86639),
            .I(N__86631));
    InMux I__20160 (
            .O(N__86638),
            .I(N__86628));
    InMux I__20159 (
            .O(N__86637),
            .I(N__86623));
    InMux I__20158 (
            .O(N__86636),
            .I(N__86623));
    Span4Mux_v I__20157 (
            .O(N__86631),
            .I(N__86620));
    LocalMux I__20156 (
            .O(N__86628),
            .I(N__86617));
    LocalMux I__20155 (
            .O(N__86623),
            .I(\c0.n31429 ));
    Odrv4 I__20154 (
            .O(N__86620),
            .I(\c0.n31429 ));
    Odrv12 I__20153 (
            .O(N__86617),
            .I(\c0.n31429 ));
    InMux I__20152 (
            .O(N__86610),
            .I(N__86601));
    InMux I__20151 (
            .O(N__86609),
            .I(N__86601));
    CascadeMux I__20150 (
            .O(N__86608),
            .I(N__86596));
    InMux I__20149 (
            .O(N__86607),
            .I(N__86593));
    InMux I__20148 (
            .O(N__86606),
            .I(N__86590));
    LocalMux I__20147 (
            .O(N__86601),
            .I(N__86587));
    CascadeMux I__20146 (
            .O(N__86600),
            .I(N__86584));
    CascadeMux I__20145 (
            .O(N__86599),
            .I(N__86580));
    InMux I__20144 (
            .O(N__86596),
            .I(N__86577));
    LocalMux I__20143 (
            .O(N__86593),
            .I(N__86570));
    LocalMux I__20142 (
            .O(N__86590),
            .I(N__86570));
    Span4Mux_v I__20141 (
            .O(N__86587),
            .I(N__86570));
    InMux I__20140 (
            .O(N__86584),
            .I(N__86567));
    InMux I__20139 (
            .O(N__86583),
            .I(N__86564));
    InMux I__20138 (
            .O(N__86580),
            .I(N__86561));
    LocalMux I__20137 (
            .O(N__86577),
            .I(N__86558));
    Span4Mux_v I__20136 (
            .O(N__86570),
            .I(N__86553));
    LocalMux I__20135 (
            .O(N__86567),
            .I(N__86553));
    LocalMux I__20134 (
            .O(N__86564),
            .I(encoder1_position_2));
    LocalMux I__20133 (
            .O(N__86561),
            .I(encoder1_position_2));
    Odrv12 I__20132 (
            .O(N__86558),
            .I(encoder1_position_2));
    Odrv4 I__20131 (
            .O(N__86553),
            .I(encoder1_position_2));
    CascadeMux I__20130 (
            .O(N__86544),
            .I(\c0.n33897_cascade_ ));
    InMux I__20129 (
            .O(N__86541),
            .I(N__86535));
    InMux I__20128 (
            .O(N__86540),
            .I(N__86535));
    LocalMux I__20127 (
            .O(N__86535),
            .I(N__86532));
    Odrv4 I__20126 (
            .O(N__86532),
            .I(\c0.n33732 ));
    CascadeMux I__20125 (
            .O(N__86529),
            .I(N__86526));
    InMux I__20124 (
            .O(N__86526),
            .I(N__86522));
    InMux I__20123 (
            .O(N__86525),
            .I(N__86519));
    LocalMux I__20122 (
            .O(N__86522),
            .I(N__86516));
    LocalMux I__20121 (
            .O(N__86519),
            .I(N__86512));
    Span4Mux_v I__20120 (
            .O(N__86516),
            .I(N__86509));
    InMux I__20119 (
            .O(N__86515),
            .I(N__86506));
    Odrv12 I__20118 (
            .O(N__86512),
            .I(\c0.n33892 ));
    Odrv4 I__20117 (
            .O(N__86509),
            .I(\c0.n33892 ));
    LocalMux I__20116 (
            .O(N__86506),
            .I(\c0.n33892 ));
    CascadeMux I__20115 (
            .O(N__86499),
            .I(N__86496));
    InMux I__20114 (
            .O(N__86496),
            .I(N__86492));
    InMux I__20113 (
            .O(N__86495),
            .I(N__86486));
    LocalMux I__20112 (
            .O(N__86492),
            .I(N__86483));
    InMux I__20111 (
            .O(N__86491),
            .I(N__86480));
    InMux I__20110 (
            .O(N__86490),
            .I(N__86477));
    InMux I__20109 (
            .O(N__86489),
            .I(N__86474));
    LocalMux I__20108 (
            .O(N__86486),
            .I(N__86470));
    Span4Mux_h I__20107 (
            .O(N__86483),
            .I(N__86461));
    LocalMux I__20106 (
            .O(N__86480),
            .I(N__86461));
    LocalMux I__20105 (
            .O(N__86477),
            .I(N__86461));
    LocalMux I__20104 (
            .O(N__86474),
            .I(N__86461));
    InMux I__20103 (
            .O(N__86473),
            .I(N__86458));
    Span4Mux_h I__20102 (
            .O(N__86470),
            .I(N__86453));
    Span4Mux_v I__20101 (
            .O(N__86461),
            .I(N__86453));
    LocalMux I__20100 (
            .O(N__86458),
            .I(encoder0_position_15));
    Odrv4 I__20099 (
            .O(N__86453),
            .I(encoder0_position_15));
    InMux I__20098 (
            .O(N__86448),
            .I(N__86445));
    LocalMux I__20097 (
            .O(N__86445),
            .I(N__86440));
    InMux I__20096 (
            .O(N__86444),
            .I(N__86435));
    InMux I__20095 (
            .O(N__86443),
            .I(N__86435));
    Odrv4 I__20094 (
            .O(N__86440),
            .I(\c0.n18895 ));
    LocalMux I__20093 (
            .O(N__86435),
            .I(\c0.n18895 ));
    CascadeMux I__20092 (
            .O(N__86430),
            .I(N__86427));
    InMux I__20091 (
            .O(N__86427),
            .I(N__86423));
    CascadeMux I__20090 (
            .O(N__86426),
            .I(N__86420));
    LocalMux I__20089 (
            .O(N__86423),
            .I(N__86416));
    InMux I__20088 (
            .O(N__86420),
            .I(N__86413));
    InMux I__20087 (
            .O(N__86419),
            .I(N__86408));
    Sp12to4 I__20086 (
            .O(N__86416),
            .I(N__86404));
    LocalMux I__20085 (
            .O(N__86413),
            .I(N__86401));
    InMux I__20084 (
            .O(N__86412),
            .I(N__86398));
    InMux I__20083 (
            .O(N__86411),
            .I(N__86395));
    LocalMux I__20082 (
            .O(N__86408),
            .I(N__86392));
    InMux I__20081 (
            .O(N__86407),
            .I(N__86389));
    Span12Mux_v I__20080 (
            .O(N__86404),
            .I(N__86386));
    Span4Mux_h I__20079 (
            .O(N__86401),
            .I(N__86379));
    LocalMux I__20078 (
            .O(N__86398),
            .I(N__86379));
    LocalMux I__20077 (
            .O(N__86395),
            .I(N__86379));
    Span4Mux_h I__20076 (
            .O(N__86392),
            .I(N__86376));
    LocalMux I__20075 (
            .O(N__86389),
            .I(encoder0_position_16));
    Odrv12 I__20074 (
            .O(N__86386),
            .I(encoder0_position_16));
    Odrv4 I__20073 (
            .O(N__86379),
            .I(encoder0_position_16));
    Odrv4 I__20072 (
            .O(N__86376),
            .I(encoder0_position_16));
    CascadeMux I__20071 (
            .O(N__86367),
            .I(N__86364));
    InMux I__20070 (
            .O(N__86364),
            .I(N__86360));
    CascadeMux I__20069 (
            .O(N__86363),
            .I(N__86357));
    LocalMux I__20068 (
            .O(N__86360),
            .I(N__86354));
    InMux I__20067 (
            .O(N__86357),
            .I(N__86349));
    Span4Mux_v I__20066 (
            .O(N__86354),
            .I(N__86345));
    InMux I__20065 (
            .O(N__86353),
            .I(N__86342));
    InMux I__20064 (
            .O(N__86352),
            .I(N__86339));
    LocalMux I__20063 (
            .O(N__86349),
            .I(N__86336));
    InMux I__20062 (
            .O(N__86348),
            .I(N__86333));
    Span4Mux_h I__20061 (
            .O(N__86345),
            .I(N__86330));
    LocalMux I__20060 (
            .O(N__86342),
            .I(N__86327));
    LocalMux I__20059 (
            .O(N__86339),
            .I(N__86324));
    Span12Mux_v I__20058 (
            .O(N__86336),
            .I(N__86321));
    LocalMux I__20057 (
            .O(N__86333),
            .I(encoder1_position_18));
    Odrv4 I__20056 (
            .O(N__86330),
            .I(encoder1_position_18));
    Odrv4 I__20055 (
            .O(N__86327),
            .I(encoder1_position_18));
    Odrv4 I__20054 (
            .O(N__86324),
            .I(encoder1_position_18));
    Odrv12 I__20053 (
            .O(N__86321),
            .I(encoder1_position_18));
    InMux I__20052 (
            .O(N__86310),
            .I(N__86305));
    InMux I__20051 (
            .O(N__86309),
            .I(N__86300));
    InMux I__20050 (
            .O(N__86308),
            .I(N__86300));
    LocalMux I__20049 (
            .O(N__86305),
            .I(N__86295));
    LocalMux I__20048 (
            .O(N__86300),
            .I(N__86295));
    Odrv12 I__20047 (
            .O(N__86295),
            .I(\c0.n33353 ));
    InMux I__20046 (
            .O(N__86292),
            .I(N__86289));
    LocalMux I__20045 (
            .O(N__86289),
            .I(N__86286));
    Span4Mux_h I__20044 (
            .O(N__86286),
            .I(N__86283));
    Odrv4 I__20043 (
            .O(N__86283),
            .I(\c0.n33318 ));
    CascadeMux I__20042 (
            .O(N__86280),
            .I(N__86277));
    InMux I__20041 (
            .O(N__86277),
            .I(N__86274));
    LocalMux I__20040 (
            .O(N__86274),
            .I(N__86268));
    InMux I__20039 (
            .O(N__86273),
            .I(N__86265));
    InMux I__20038 (
            .O(N__86272),
            .I(N__86262));
    InMux I__20037 (
            .O(N__86271),
            .I(N__86259));
    Span4Mux_v I__20036 (
            .O(N__86268),
            .I(N__86255));
    LocalMux I__20035 (
            .O(N__86265),
            .I(N__86252));
    LocalMux I__20034 (
            .O(N__86262),
            .I(N__86247));
    LocalMux I__20033 (
            .O(N__86259),
            .I(N__86247));
    InMux I__20032 (
            .O(N__86258),
            .I(N__86244));
    Span4Mux_v I__20031 (
            .O(N__86255),
            .I(N__86241));
    Span4Mux_v I__20030 (
            .O(N__86252),
            .I(N__86238));
    Span4Mux_h I__20029 (
            .O(N__86247),
            .I(N__86235));
    LocalMux I__20028 (
            .O(N__86244),
            .I(encoder1_position_30));
    Odrv4 I__20027 (
            .O(N__86241),
            .I(encoder1_position_30));
    Odrv4 I__20026 (
            .O(N__86238),
            .I(encoder1_position_30));
    Odrv4 I__20025 (
            .O(N__86235),
            .I(encoder1_position_30));
    InMux I__20024 (
            .O(N__86226),
            .I(N__86222));
    InMux I__20023 (
            .O(N__86225),
            .I(N__86219));
    LocalMux I__20022 (
            .O(N__86222),
            .I(\c0.n33487 ));
    LocalMux I__20021 (
            .O(N__86219),
            .I(\c0.n33487 ));
    InMux I__20020 (
            .O(N__86214),
            .I(N__86211));
    LocalMux I__20019 (
            .O(N__86211),
            .I(N__86208));
    Odrv12 I__20018 (
            .O(N__86208),
            .I(n2317));
    CascadeMux I__20017 (
            .O(N__86205),
            .I(N__86202));
    InMux I__20016 (
            .O(N__86202),
            .I(N__86199));
    LocalMux I__20015 (
            .O(N__86199),
            .I(N__86195));
    InMux I__20014 (
            .O(N__86198),
            .I(N__86192));
    Span4Mux_v I__20013 (
            .O(N__86195),
            .I(N__86187));
    LocalMux I__20012 (
            .O(N__86192),
            .I(N__86187));
    Span4Mux_h I__20011 (
            .O(N__86187),
            .I(N__86178));
    InMux I__20010 (
            .O(N__86186),
            .I(N__86175));
    InMux I__20009 (
            .O(N__86185),
            .I(N__86170));
    InMux I__20008 (
            .O(N__86184),
            .I(N__86170));
    InMux I__20007 (
            .O(N__86183),
            .I(N__86165));
    InMux I__20006 (
            .O(N__86182),
            .I(N__86165));
    InMux I__20005 (
            .O(N__86181),
            .I(N__86162));
    Span4Mux_h I__20004 (
            .O(N__86178),
            .I(N__86159));
    LocalMux I__20003 (
            .O(N__86175),
            .I(N__86156));
    LocalMux I__20002 (
            .O(N__86170),
            .I(N__86151));
    LocalMux I__20001 (
            .O(N__86165),
            .I(N__86151));
    LocalMux I__20000 (
            .O(N__86162),
            .I(encoder0_position_28));
    Odrv4 I__19999 (
            .O(N__86159),
            .I(encoder0_position_28));
    Odrv4 I__19998 (
            .O(N__86156),
            .I(encoder0_position_28));
    Odrv4 I__19997 (
            .O(N__86151),
            .I(encoder0_position_28));
    InMux I__19996 (
            .O(N__86142),
            .I(N__86132));
    InMux I__19995 (
            .O(N__86141),
            .I(N__86132));
    InMux I__19994 (
            .O(N__86140),
            .I(N__86129));
    InMux I__19993 (
            .O(N__86139),
            .I(N__86126));
    InMux I__19992 (
            .O(N__86138),
            .I(N__86121));
    InMux I__19991 (
            .O(N__86137),
            .I(N__86121));
    LocalMux I__19990 (
            .O(N__86132),
            .I(N__86094));
    LocalMux I__19989 (
            .O(N__86129),
            .I(N__86094));
    LocalMux I__19988 (
            .O(N__86126),
            .I(N__86094));
    LocalMux I__19987 (
            .O(N__86121),
            .I(N__86094));
    InMux I__19986 (
            .O(N__86120),
            .I(N__86087));
    InMux I__19985 (
            .O(N__86119),
            .I(N__86087));
    InMux I__19984 (
            .O(N__86118),
            .I(N__86087));
    InMux I__19983 (
            .O(N__86117),
            .I(N__86082));
    InMux I__19982 (
            .O(N__86116),
            .I(N__86082));
    InMux I__19981 (
            .O(N__86115),
            .I(N__86077));
    InMux I__19980 (
            .O(N__86114),
            .I(N__86074));
    InMux I__19979 (
            .O(N__86113),
            .I(N__86071));
    InMux I__19978 (
            .O(N__86112),
            .I(N__86064));
    InMux I__19977 (
            .O(N__86111),
            .I(N__86064));
    InMux I__19976 (
            .O(N__86110),
            .I(N__86064));
    InMux I__19975 (
            .O(N__86109),
            .I(N__86061));
    InMux I__19974 (
            .O(N__86108),
            .I(N__86056));
    InMux I__19973 (
            .O(N__86107),
            .I(N__86056));
    InMux I__19972 (
            .O(N__86106),
            .I(N__86047));
    InMux I__19971 (
            .O(N__86105),
            .I(N__86047));
    InMux I__19970 (
            .O(N__86104),
            .I(N__86047));
    InMux I__19969 (
            .O(N__86103),
            .I(N__86047));
    Span4Mux_v I__19968 (
            .O(N__86094),
            .I(N__86038));
    LocalMux I__19967 (
            .O(N__86087),
            .I(N__86033));
    LocalMux I__19966 (
            .O(N__86082),
            .I(N__86033));
    InMux I__19965 (
            .O(N__86081),
            .I(N__86030));
    InMux I__19964 (
            .O(N__86080),
            .I(N__86027));
    LocalMux I__19963 (
            .O(N__86077),
            .I(N__86022));
    LocalMux I__19962 (
            .O(N__86074),
            .I(N__86022));
    LocalMux I__19961 (
            .O(N__86071),
            .I(N__86013));
    LocalMux I__19960 (
            .O(N__86064),
            .I(N__86013));
    LocalMux I__19959 (
            .O(N__86061),
            .I(N__86013));
    LocalMux I__19958 (
            .O(N__86056),
            .I(N__86013));
    LocalMux I__19957 (
            .O(N__86047),
            .I(N__86010));
    InMux I__19956 (
            .O(N__86046),
            .I(N__86007));
    InMux I__19955 (
            .O(N__86045),
            .I(N__86002));
    InMux I__19954 (
            .O(N__86044),
            .I(N__86002));
    InMux I__19953 (
            .O(N__86043),
            .I(N__85997));
    InMux I__19952 (
            .O(N__86042),
            .I(N__85997));
    InMux I__19951 (
            .O(N__86041),
            .I(N__85994));
    Span4Mux_h I__19950 (
            .O(N__86038),
            .I(N__85989));
    Span4Mux_v I__19949 (
            .O(N__86033),
            .I(N__85989));
    LocalMux I__19948 (
            .O(N__86030),
            .I(N__85986));
    LocalMux I__19947 (
            .O(N__86027),
            .I(N__85983));
    Span4Mux_v I__19946 (
            .O(N__86022),
            .I(N__85972));
    Span4Mux_v I__19945 (
            .O(N__86013),
            .I(N__85972));
    Span4Mux_h I__19944 (
            .O(N__86010),
            .I(N__85972));
    LocalMux I__19943 (
            .O(N__86007),
            .I(N__85972));
    LocalMux I__19942 (
            .O(N__86002),
            .I(N__85972));
    LocalMux I__19941 (
            .O(N__85997),
            .I(N__85967));
    LocalMux I__19940 (
            .O(N__85994),
            .I(N__85967));
    Span4Mux_h I__19939 (
            .O(N__85989),
            .I(N__85964));
    Span4Mux_v I__19938 (
            .O(N__85986),
            .I(N__85959));
    Span4Mux_v I__19937 (
            .O(N__85983),
            .I(N__85959));
    Span4Mux_h I__19936 (
            .O(N__85972),
            .I(N__85954));
    Span4Mux_v I__19935 (
            .O(N__85967),
            .I(N__85954));
    Span4Mux_h I__19934 (
            .O(N__85964),
            .I(N__85951));
    Span4Mux_h I__19933 (
            .O(N__85959),
            .I(N__85946));
    Span4Mux_h I__19932 (
            .O(N__85954),
            .I(N__85946));
    Odrv4 I__19931 (
            .O(N__85951),
            .I(count_enable));
    Odrv4 I__19930 (
            .O(N__85946),
            .I(count_enable));
    InMux I__19929 (
            .O(N__85941),
            .I(N__85938));
    LocalMux I__19928 (
            .O(N__85938),
            .I(N__85935));
    Span4Mux_h I__19927 (
            .O(N__85935),
            .I(N__85932));
    Odrv4 I__19926 (
            .O(N__85932),
            .I(n2319));
    InMux I__19925 (
            .O(N__85929),
            .I(N__85926));
    LocalMux I__19924 (
            .O(N__85926),
            .I(N__85923));
    Span4Mux_h I__19923 (
            .O(N__85923),
            .I(N__85917));
    CascadeMux I__19922 (
            .O(N__85922),
            .I(N__85914));
    InMux I__19921 (
            .O(N__85921),
            .I(N__85911));
    InMux I__19920 (
            .O(N__85920),
            .I(N__85908));
    Span4Mux_h I__19919 (
            .O(N__85917),
            .I(N__85905));
    InMux I__19918 (
            .O(N__85914),
            .I(N__85902));
    LocalMux I__19917 (
            .O(N__85911),
            .I(N__85897));
    LocalMux I__19916 (
            .O(N__85908),
            .I(N__85893));
    Span4Mux_v I__19915 (
            .O(N__85905),
            .I(N__85888));
    LocalMux I__19914 (
            .O(N__85902),
            .I(N__85888));
    CascadeMux I__19913 (
            .O(N__85901),
            .I(N__85885));
    InMux I__19912 (
            .O(N__85900),
            .I(N__85882));
    Span4Mux_v I__19911 (
            .O(N__85897),
            .I(N__85879));
    InMux I__19910 (
            .O(N__85896),
            .I(N__85876));
    Span4Mux_h I__19909 (
            .O(N__85893),
            .I(N__85871));
    Span4Mux_v I__19908 (
            .O(N__85888),
            .I(N__85871));
    InMux I__19907 (
            .O(N__85885),
            .I(N__85868));
    LocalMux I__19906 (
            .O(N__85882),
            .I(encoder0_position_26));
    Odrv4 I__19905 (
            .O(N__85879),
            .I(encoder0_position_26));
    LocalMux I__19904 (
            .O(N__85876),
            .I(encoder0_position_26));
    Odrv4 I__19903 (
            .O(N__85871),
            .I(encoder0_position_26));
    LocalMux I__19902 (
            .O(N__85868),
            .I(encoder0_position_26));
    CascadeMux I__19901 (
            .O(N__85857),
            .I(N__85854));
    InMux I__19900 (
            .O(N__85854),
            .I(N__85851));
    LocalMux I__19899 (
            .O(N__85851),
            .I(N__85848));
    Odrv4 I__19898 (
            .O(N__85848),
            .I(\c0.n33579 ));
    CascadeMux I__19897 (
            .O(N__85845),
            .I(N__85841));
    CascadeMux I__19896 (
            .O(N__85844),
            .I(N__85837));
    InMux I__19895 (
            .O(N__85841),
            .I(N__85834));
    CascadeMux I__19894 (
            .O(N__85840),
            .I(N__85831));
    InMux I__19893 (
            .O(N__85837),
            .I(N__85827));
    LocalMux I__19892 (
            .O(N__85834),
            .I(N__85824));
    InMux I__19891 (
            .O(N__85831),
            .I(N__85821));
    InMux I__19890 (
            .O(N__85830),
            .I(N__85818));
    LocalMux I__19889 (
            .O(N__85827),
            .I(N__85814));
    Span4Mux_h I__19888 (
            .O(N__85824),
            .I(N__85807));
    LocalMux I__19887 (
            .O(N__85821),
            .I(N__85807));
    LocalMux I__19886 (
            .O(N__85818),
            .I(N__85807));
    InMux I__19885 (
            .O(N__85817),
            .I(N__85804));
    Span4Mux_h I__19884 (
            .O(N__85814),
            .I(N__85801));
    Span4Mux_v I__19883 (
            .O(N__85807),
            .I(N__85798));
    LocalMux I__19882 (
            .O(N__85804),
            .I(encoder1_position_4));
    Odrv4 I__19881 (
            .O(N__85801),
            .I(encoder1_position_4));
    Odrv4 I__19880 (
            .O(N__85798),
            .I(encoder1_position_4));
    CascadeMux I__19879 (
            .O(N__85791),
            .I(\c0.n6_adj_4558_cascade_ ));
    InMux I__19878 (
            .O(N__85788),
            .I(N__85784));
    InMux I__19877 (
            .O(N__85787),
            .I(N__85778));
    LocalMux I__19876 (
            .O(N__85784),
            .I(N__85774));
    InMux I__19875 (
            .O(N__85783),
            .I(N__85769));
    InMux I__19874 (
            .O(N__85782),
            .I(N__85769));
    InMux I__19873 (
            .O(N__85781),
            .I(N__85766));
    LocalMux I__19872 (
            .O(N__85778),
            .I(N__85763));
    InMux I__19871 (
            .O(N__85777),
            .I(N__85760));
    Span4Mux_h I__19870 (
            .O(N__85774),
            .I(N__85757));
    LocalMux I__19869 (
            .O(N__85769),
            .I(N__85754));
    LocalMux I__19868 (
            .O(N__85766),
            .I(encoder0_position_14));
    Odrv4 I__19867 (
            .O(N__85763),
            .I(encoder0_position_14));
    LocalMux I__19866 (
            .O(N__85760),
            .I(encoder0_position_14));
    Odrv4 I__19865 (
            .O(N__85757),
            .I(encoder0_position_14));
    Odrv4 I__19864 (
            .O(N__85754),
            .I(encoder0_position_14));
    CascadeMux I__19863 (
            .O(N__85743),
            .I(N__85740));
    InMux I__19862 (
            .O(N__85740),
            .I(N__85736));
    CascadeMux I__19861 (
            .O(N__85739),
            .I(N__85732));
    LocalMux I__19860 (
            .O(N__85736),
            .I(N__85729));
    InMux I__19859 (
            .O(N__85735),
            .I(N__85726));
    InMux I__19858 (
            .O(N__85732),
            .I(N__85723));
    Span4Mux_v I__19857 (
            .O(N__85729),
            .I(N__85720));
    LocalMux I__19856 (
            .O(N__85726),
            .I(N__85717));
    LocalMux I__19855 (
            .O(N__85723),
            .I(N__85713));
    Span4Mux_h I__19854 (
            .O(N__85720),
            .I(N__85708));
    Span4Mux_v I__19853 (
            .O(N__85717),
            .I(N__85708));
    InMux I__19852 (
            .O(N__85716),
            .I(N__85705));
    Span4Mux_h I__19851 (
            .O(N__85713),
            .I(N__85700));
    Span4Mux_v I__19850 (
            .O(N__85708),
            .I(N__85700));
    LocalMux I__19849 (
            .O(N__85705),
            .I(encoder1_position_5));
    Odrv4 I__19848 (
            .O(N__85700),
            .I(encoder1_position_5));
    CascadeMux I__19847 (
            .O(N__85695),
            .I(\c0.n18499_cascade_ ));
    CascadeMux I__19846 (
            .O(N__85692),
            .I(\c0.n33569_cascade_ ));
    InMux I__19845 (
            .O(N__85689),
            .I(N__85685));
    InMux I__19844 (
            .O(N__85688),
            .I(N__85680));
    LocalMux I__19843 (
            .O(N__85685),
            .I(N__85677));
    InMux I__19842 (
            .O(N__85684),
            .I(N__85671));
    InMux I__19841 (
            .O(N__85683),
            .I(N__85668));
    LocalMux I__19840 (
            .O(N__85680),
            .I(N__85665));
    Span4Mux_h I__19839 (
            .O(N__85677),
            .I(N__85662));
    InMux I__19838 (
            .O(N__85676),
            .I(N__85657));
    InMux I__19837 (
            .O(N__85675),
            .I(N__85657));
    InMux I__19836 (
            .O(N__85674),
            .I(N__85654));
    LocalMux I__19835 (
            .O(N__85671),
            .I(N__85649));
    LocalMux I__19834 (
            .O(N__85668),
            .I(N__85649));
    Span4Mux_h I__19833 (
            .O(N__85665),
            .I(N__85646));
    Span4Mux_h I__19832 (
            .O(N__85662),
            .I(N__85641));
    LocalMux I__19831 (
            .O(N__85657),
            .I(N__85641));
    LocalMux I__19830 (
            .O(N__85654),
            .I(encoder1_position_31));
    Odrv4 I__19829 (
            .O(N__85649),
            .I(encoder1_position_31));
    Odrv4 I__19828 (
            .O(N__85646),
            .I(encoder1_position_31));
    Odrv4 I__19827 (
            .O(N__85641),
            .I(encoder1_position_31));
    CascadeMux I__19826 (
            .O(N__85632),
            .I(N__85627));
    CascadeMux I__19825 (
            .O(N__85631),
            .I(N__85622));
    InMux I__19824 (
            .O(N__85630),
            .I(N__85619));
    InMux I__19823 (
            .O(N__85627),
            .I(N__85616));
    InMux I__19822 (
            .O(N__85626),
            .I(N__85613));
    CascadeMux I__19821 (
            .O(N__85625),
            .I(N__85610));
    InMux I__19820 (
            .O(N__85622),
            .I(N__85607));
    LocalMux I__19819 (
            .O(N__85619),
            .I(N__85604));
    LocalMux I__19818 (
            .O(N__85616),
            .I(N__85600));
    LocalMux I__19817 (
            .O(N__85613),
            .I(N__85597));
    InMux I__19816 (
            .O(N__85610),
            .I(N__85594));
    LocalMux I__19815 (
            .O(N__85607),
            .I(N__85590));
    Span4Mux_h I__19814 (
            .O(N__85604),
            .I(N__85587));
    CascadeMux I__19813 (
            .O(N__85603),
            .I(N__85584));
    Span4Mux_v I__19812 (
            .O(N__85600),
            .I(N__85581));
    Span4Mux_v I__19811 (
            .O(N__85597),
            .I(N__85576));
    LocalMux I__19810 (
            .O(N__85594),
            .I(N__85576));
    InMux I__19809 (
            .O(N__85593),
            .I(N__85573));
    Span4Mux_h I__19808 (
            .O(N__85590),
            .I(N__85570));
    Sp12to4 I__19807 (
            .O(N__85587),
            .I(N__85567));
    InMux I__19806 (
            .O(N__85584),
            .I(N__85564));
    Span4Mux_h I__19805 (
            .O(N__85581),
            .I(N__85559));
    Span4Mux_h I__19804 (
            .O(N__85576),
            .I(N__85559));
    LocalMux I__19803 (
            .O(N__85573),
            .I(encoder0_position_0));
    Odrv4 I__19802 (
            .O(N__85570),
            .I(encoder0_position_0));
    Odrv12 I__19801 (
            .O(N__85567),
            .I(encoder0_position_0));
    LocalMux I__19800 (
            .O(N__85564),
            .I(encoder0_position_0));
    Odrv4 I__19799 (
            .O(N__85559),
            .I(encoder0_position_0));
    InMux I__19798 (
            .O(N__85548),
            .I(N__85545));
    LocalMux I__19797 (
            .O(N__85545),
            .I(\c0.n6_adj_4565 ));
    InMux I__19796 (
            .O(N__85542),
            .I(N__85538));
    InMux I__19795 (
            .O(N__85541),
            .I(N__85534));
    LocalMux I__19794 (
            .O(N__85538),
            .I(N__85531));
    InMux I__19793 (
            .O(N__85537),
            .I(N__85528));
    LocalMux I__19792 (
            .O(N__85534),
            .I(N__85525));
    Span4Mux_h I__19791 (
            .O(N__85531),
            .I(N__85522));
    LocalMux I__19790 (
            .O(N__85528),
            .I(\c0.n33897 ));
    Odrv12 I__19789 (
            .O(N__85525),
            .I(\c0.n33897 ));
    Odrv4 I__19788 (
            .O(N__85522),
            .I(\c0.n33897 ));
    CascadeMux I__19787 (
            .O(N__85515),
            .I(N__85512));
    InMux I__19786 (
            .O(N__85512),
            .I(N__85507));
    InMux I__19785 (
            .O(N__85511),
            .I(N__85501));
    InMux I__19784 (
            .O(N__85510),
            .I(N__85501));
    LocalMux I__19783 (
            .O(N__85507),
            .I(N__85497));
    CascadeMux I__19782 (
            .O(N__85506),
            .I(N__85494));
    LocalMux I__19781 (
            .O(N__85501),
            .I(N__85491));
    InMux I__19780 (
            .O(N__85500),
            .I(N__85487));
    Span4Mux_h I__19779 (
            .O(N__85497),
            .I(N__85484));
    InMux I__19778 (
            .O(N__85494),
            .I(N__85481));
    Span4Mux_h I__19777 (
            .O(N__85491),
            .I(N__85478));
    InMux I__19776 (
            .O(N__85490),
            .I(N__85475));
    LocalMux I__19775 (
            .O(N__85487),
            .I(encoder1_position_21));
    Odrv4 I__19774 (
            .O(N__85484),
            .I(encoder1_position_21));
    LocalMux I__19773 (
            .O(N__85481),
            .I(encoder1_position_21));
    Odrv4 I__19772 (
            .O(N__85478),
            .I(encoder1_position_21));
    LocalMux I__19771 (
            .O(N__85475),
            .I(encoder1_position_21));
    CascadeMux I__19770 (
            .O(N__85464),
            .I(N__85460));
    InMux I__19769 (
            .O(N__85463),
            .I(N__85456));
    InMux I__19768 (
            .O(N__85460),
            .I(N__85452));
    InMux I__19767 (
            .O(N__85459),
            .I(N__85448));
    LocalMux I__19766 (
            .O(N__85456),
            .I(N__85445));
    InMux I__19765 (
            .O(N__85455),
            .I(N__85442));
    LocalMux I__19764 (
            .O(N__85452),
            .I(N__85438));
    CascadeMux I__19763 (
            .O(N__85451),
            .I(N__85435));
    LocalMux I__19762 (
            .O(N__85448),
            .I(N__85432));
    Span4Mux_v I__19761 (
            .O(N__85445),
            .I(N__85427));
    LocalMux I__19760 (
            .O(N__85442),
            .I(N__85427));
    InMux I__19759 (
            .O(N__85441),
            .I(N__85424));
    Sp12to4 I__19758 (
            .O(N__85438),
            .I(N__85421));
    InMux I__19757 (
            .O(N__85435),
            .I(N__85418));
    Span4Mux_v I__19756 (
            .O(N__85432),
            .I(N__85415));
    Span4Mux_h I__19755 (
            .O(N__85427),
            .I(N__85412));
    LocalMux I__19754 (
            .O(N__85424),
            .I(encoder0_position_3));
    Odrv12 I__19753 (
            .O(N__85421),
            .I(encoder0_position_3));
    LocalMux I__19752 (
            .O(N__85418),
            .I(encoder0_position_3));
    Odrv4 I__19751 (
            .O(N__85415),
            .I(encoder0_position_3));
    Odrv4 I__19750 (
            .O(N__85412),
            .I(encoder0_position_3));
    CascadeMux I__19749 (
            .O(N__85401),
            .I(N__85398));
    InMux I__19748 (
            .O(N__85398),
            .I(N__85395));
    LocalMux I__19747 (
            .O(N__85395),
            .I(N__85392));
    Span4Mux_h I__19746 (
            .O(N__85392),
            .I(N__85388));
    InMux I__19745 (
            .O(N__85391),
            .I(N__85385));
    Odrv4 I__19744 (
            .O(N__85388),
            .I(\c0.n18218 ));
    LocalMux I__19743 (
            .O(N__85385),
            .I(\c0.n18218 ));
    InMux I__19742 (
            .O(N__85380),
            .I(N__85375));
    CascadeMux I__19741 (
            .O(N__85379),
            .I(N__85371));
    InMux I__19740 (
            .O(N__85378),
            .I(N__85368));
    LocalMux I__19739 (
            .O(N__85375),
            .I(N__85365));
    InMux I__19738 (
            .O(N__85374),
            .I(N__85362));
    InMux I__19737 (
            .O(N__85371),
            .I(N__85358));
    LocalMux I__19736 (
            .O(N__85368),
            .I(N__85355));
    Span4Mux_h I__19735 (
            .O(N__85365),
            .I(N__85352));
    LocalMux I__19734 (
            .O(N__85362),
            .I(N__85349));
    InMux I__19733 (
            .O(N__85361),
            .I(N__85346));
    LocalMux I__19732 (
            .O(N__85358),
            .I(N__85341));
    Span4Mux_h I__19731 (
            .O(N__85355),
            .I(N__85341));
    Span4Mux_v I__19730 (
            .O(N__85352),
            .I(N__85338));
    Span4Mux_h I__19729 (
            .O(N__85349),
            .I(N__85335));
    LocalMux I__19728 (
            .O(N__85346),
            .I(encoder0_position_4));
    Odrv4 I__19727 (
            .O(N__85341),
            .I(encoder0_position_4));
    Odrv4 I__19726 (
            .O(N__85338),
            .I(encoder0_position_4));
    Odrv4 I__19725 (
            .O(N__85335),
            .I(encoder0_position_4));
    CascadeMux I__19724 (
            .O(N__85326),
            .I(\c0.n18469_cascade_ ));
    InMux I__19723 (
            .O(N__85323),
            .I(N__85318));
    InMux I__19722 (
            .O(N__85322),
            .I(N__85315));
    InMux I__19721 (
            .O(N__85321),
            .I(N__85312));
    LocalMux I__19720 (
            .O(N__85318),
            .I(N__85305));
    LocalMux I__19719 (
            .O(N__85315),
            .I(N__85305));
    LocalMux I__19718 (
            .O(N__85312),
            .I(N__85305));
    Span4Mux_v I__19717 (
            .O(N__85305),
            .I(N__85302));
    Odrv4 I__19716 (
            .O(N__85302),
            .I(\c0.n33681 ));
    CascadeMux I__19715 (
            .O(N__85299),
            .I(\c0.n18241_cascade_ ));
    InMux I__19714 (
            .O(N__85296),
            .I(N__85293));
    LocalMux I__19713 (
            .O(N__85293),
            .I(\c0.n10_adj_4528 ));
    CascadeMux I__19712 (
            .O(N__85290),
            .I(\c0.n14_adj_4527_cascade_ ));
    CascadeMux I__19711 (
            .O(N__85287),
            .I(\c0.n31511_cascade_ ));
    InMux I__19710 (
            .O(N__85284),
            .I(N__85270));
    InMux I__19709 (
            .O(N__85283),
            .I(N__85263));
    InMux I__19708 (
            .O(N__85282),
            .I(N__85263));
    InMux I__19707 (
            .O(N__85281),
            .I(N__85263));
    InMux I__19706 (
            .O(N__85280),
            .I(N__85256));
    InMux I__19705 (
            .O(N__85279),
            .I(N__85256));
    InMux I__19704 (
            .O(N__85278),
            .I(N__85256));
    InMux I__19703 (
            .O(N__85277),
            .I(N__85253));
    CascadeMux I__19702 (
            .O(N__85276),
            .I(N__85247));
    CascadeMux I__19701 (
            .O(N__85275),
            .I(N__85242));
    InMux I__19700 (
            .O(N__85274),
            .I(N__85239));
    InMux I__19699 (
            .O(N__85273),
            .I(N__85236));
    LocalMux I__19698 (
            .O(N__85270),
            .I(N__85220));
    LocalMux I__19697 (
            .O(N__85263),
            .I(N__85220));
    LocalMux I__19696 (
            .O(N__85256),
            .I(N__85220));
    LocalMux I__19695 (
            .O(N__85253),
            .I(N__85217));
    CascadeMux I__19694 (
            .O(N__85252),
            .I(N__85206));
    InMux I__19693 (
            .O(N__85251),
            .I(N__85200));
    CascadeMux I__19692 (
            .O(N__85250),
            .I(N__85194));
    InMux I__19691 (
            .O(N__85247),
            .I(N__85191));
    InMux I__19690 (
            .O(N__85246),
            .I(N__85184));
    InMux I__19689 (
            .O(N__85245),
            .I(N__85184));
    InMux I__19688 (
            .O(N__85242),
            .I(N__85184));
    LocalMux I__19687 (
            .O(N__85239),
            .I(N__85179));
    LocalMux I__19686 (
            .O(N__85236),
            .I(N__85179));
    InMux I__19685 (
            .O(N__85235),
            .I(N__85166));
    InMux I__19684 (
            .O(N__85234),
            .I(N__85166));
    CascadeMux I__19683 (
            .O(N__85233),
            .I(N__85155));
    CascadeMux I__19682 (
            .O(N__85232),
            .I(N__85152));
    CascadeMux I__19681 (
            .O(N__85231),
            .I(N__85147));
    InMux I__19680 (
            .O(N__85230),
            .I(N__85143));
    InMux I__19679 (
            .O(N__85229),
            .I(N__85136));
    InMux I__19678 (
            .O(N__85228),
            .I(N__85136));
    InMux I__19677 (
            .O(N__85227),
            .I(N__85133));
    Span4Mux_v I__19676 (
            .O(N__85220),
            .I(N__85128));
    Span4Mux_v I__19675 (
            .O(N__85217),
            .I(N__85128));
    InMux I__19674 (
            .O(N__85216),
            .I(N__85117));
    InMux I__19673 (
            .O(N__85215),
            .I(N__85117));
    InMux I__19672 (
            .O(N__85214),
            .I(N__85117));
    InMux I__19671 (
            .O(N__85213),
            .I(N__85117));
    InMux I__19670 (
            .O(N__85212),
            .I(N__85117));
    InMux I__19669 (
            .O(N__85211),
            .I(N__85108));
    InMux I__19668 (
            .O(N__85210),
            .I(N__85108));
    InMux I__19667 (
            .O(N__85209),
            .I(N__85108));
    InMux I__19666 (
            .O(N__85206),
            .I(N__85108));
    InMux I__19665 (
            .O(N__85205),
            .I(N__85101));
    InMux I__19664 (
            .O(N__85204),
            .I(N__85101));
    InMux I__19663 (
            .O(N__85203),
            .I(N__85101));
    LocalMux I__19662 (
            .O(N__85200),
            .I(N__85097));
    InMux I__19661 (
            .O(N__85199),
            .I(N__85093));
    InMux I__19660 (
            .O(N__85198),
            .I(N__85088));
    InMux I__19659 (
            .O(N__85197),
            .I(N__85088));
    InMux I__19658 (
            .O(N__85194),
            .I(N__85085));
    LocalMux I__19657 (
            .O(N__85191),
            .I(N__85082));
    LocalMux I__19656 (
            .O(N__85184),
            .I(N__85077));
    Span4Mux_h I__19655 (
            .O(N__85179),
            .I(N__85077));
    CascadeMux I__19654 (
            .O(N__85178),
            .I(N__85073));
    CascadeMux I__19653 (
            .O(N__85177),
            .I(N__85063));
    InMux I__19652 (
            .O(N__85176),
            .I(N__85060));
    CascadeMux I__19651 (
            .O(N__85175),
            .I(N__85057));
    CascadeMux I__19650 (
            .O(N__85174),
            .I(N__85053));
    InMux I__19649 (
            .O(N__85173),
            .I(N__85045));
    InMux I__19648 (
            .O(N__85172),
            .I(N__85045));
    InMux I__19647 (
            .O(N__85171),
            .I(N__85045));
    LocalMux I__19646 (
            .O(N__85166),
            .I(N__85042));
    CascadeMux I__19645 (
            .O(N__85165),
            .I(N__85037));
    InMux I__19644 (
            .O(N__85164),
            .I(N__85034));
    CascadeMux I__19643 (
            .O(N__85163),
            .I(N__85030));
    InMux I__19642 (
            .O(N__85162),
            .I(N__85021));
    InMux I__19641 (
            .O(N__85161),
            .I(N__85021));
    InMux I__19640 (
            .O(N__85160),
            .I(N__85021));
    InMux I__19639 (
            .O(N__85159),
            .I(N__85012));
    InMux I__19638 (
            .O(N__85158),
            .I(N__85012));
    InMux I__19637 (
            .O(N__85155),
            .I(N__85012));
    InMux I__19636 (
            .O(N__85152),
            .I(N__85012));
    InMux I__19635 (
            .O(N__85151),
            .I(N__85007));
    InMux I__19634 (
            .O(N__85150),
            .I(N__85007));
    InMux I__19633 (
            .O(N__85147),
            .I(N__85004));
    InMux I__19632 (
            .O(N__85146),
            .I(N__85001));
    LocalMux I__19631 (
            .O(N__85143),
            .I(N__84998));
    InMux I__19630 (
            .O(N__85142),
            .I(N__84993));
    InMux I__19629 (
            .O(N__85141),
            .I(N__84993));
    LocalMux I__19628 (
            .O(N__85136),
            .I(N__84990));
    LocalMux I__19627 (
            .O(N__85133),
            .I(N__84985));
    Span4Mux_h I__19626 (
            .O(N__85128),
            .I(N__84985));
    LocalMux I__19625 (
            .O(N__85117),
            .I(N__84980));
    LocalMux I__19624 (
            .O(N__85108),
            .I(N__84980));
    LocalMux I__19623 (
            .O(N__85101),
            .I(N__84977));
    InMux I__19622 (
            .O(N__85100),
            .I(N__84974));
    Span12Mux_h I__19621 (
            .O(N__85097),
            .I(N__84971));
    InMux I__19620 (
            .O(N__85096),
            .I(N__84968));
    LocalMux I__19619 (
            .O(N__85093),
            .I(N__84965));
    LocalMux I__19618 (
            .O(N__85088),
            .I(N__84958));
    LocalMux I__19617 (
            .O(N__85085),
            .I(N__84958));
    Span4Mux_h I__19616 (
            .O(N__85082),
            .I(N__84958));
    Span4Mux_h I__19615 (
            .O(N__85077),
            .I(N__84955));
    InMux I__19614 (
            .O(N__85076),
            .I(N__84950));
    InMux I__19613 (
            .O(N__85073),
            .I(N__84950));
    InMux I__19612 (
            .O(N__85072),
            .I(N__84945));
    InMux I__19611 (
            .O(N__85071),
            .I(N__84945));
    InMux I__19610 (
            .O(N__85070),
            .I(N__84940));
    InMux I__19609 (
            .O(N__85069),
            .I(N__84940));
    InMux I__19608 (
            .O(N__85068),
            .I(N__84931));
    InMux I__19607 (
            .O(N__85067),
            .I(N__84931));
    InMux I__19606 (
            .O(N__85066),
            .I(N__84931));
    InMux I__19605 (
            .O(N__85063),
            .I(N__84931));
    LocalMux I__19604 (
            .O(N__85060),
            .I(N__84928));
    InMux I__19603 (
            .O(N__85057),
            .I(N__84921));
    InMux I__19602 (
            .O(N__85056),
            .I(N__84921));
    InMux I__19601 (
            .O(N__85053),
            .I(N__84921));
    InMux I__19600 (
            .O(N__85052),
            .I(N__84918));
    LocalMux I__19599 (
            .O(N__85045),
            .I(N__84913));
    Span4Mux_v I__19598 (
            .O(N__85042),
            .I(N__84913));
    InMux I__19597 (
            .O(N__85041),
            .I(N__84906));
    InMux I__19596 (
            .O(N__85040),
            .I(N__84906));
    InMux I__19595 (
            .O(N__85037),
            .I(N__84906));
    LocalMux I__19594 (
            .O(N__85034),
            .I(N__84903));
    InMux I__19593 (
            .O(N__85033),
            .I(N__84898));
    InMux I__19592 (
            .O(N__85030),
            .I(N__84898));
    InMux I__19591 (
            .O(N__85029),
            .I(N__84893));
    InMux I__19590 (
            .O(N__85028),
            .I(N__84893));
    LocalMux I__19589 (
            .O(N__85021),
            .I(N__84890));
    LocalMux I__19588 (
            .O(N__85012),
            .I(N__84881));
    LocalMux I__19587 (
            .O(N__85007),
            .I(N__84881));
    LocalMux I__19586 (
            .O(N__85004),
            .I(N__84881));
    LocalMux I__19585 (
            .O(N__85001),
            .I(N__84881));
    Span4Mux_v I__19584 (
            .O(N__84998),
            .I(N__84878));
    LocalMux I__19583 (
            .O(N__84993),
            .I(N__84869));
    Span4Mux_h I__19582 (
            .O(N__84990),
            .I(N__84869));
    Span4Mux_v I__19581 (
            .O(N__84985),
            .I(N__84869));
    Span4Mux_v I__19580 (
            .O(N__84980),
            .I(N__84869));
    Sp12to4 I__19579 (
            .O(N__84977),
            .I(N__84864));
    LocalMux I__19578 (
            .O(N__84974),
            .I(N__84864));
    Span12Mux_h I__19577 (
            .O(N__84971),
            .I(N__84861));
    LocalMux I__19576 (
            .O(N__84968),
            .I(N__84850));
    Span4Mux_v I__19575 (
            .O(N__84965),
            .I(N__84850));
    Span4Mux_h I__19574 (
            .O(N__84958),
            .I(N__84850));
    Span4Mux_v I__19573 (
            .O(N__84955),
            .I(N__84850));
    LocalMux I__19572 (
            .O(N__84950),
            .I(N__84850));
    LocalMux I__19571 (
            .O(N__84945),
            .I(N__84845));
    LocalMux I__19570 (
            .O(N__84940),
            .I(N__84845));
    LocalMux I__19569 (
            .O(N__84931),
            .I(N__84838));
    Span4Mux_v I__19568 (
            .O(N__84928),
            .I(N__84838));
    LocalMux I__19567 (
            .O(N__84921),
            .I(N__84838));
    LocalMux I__19566 (
            .O(N__84918),
            .I(N__84833));
    Span4Mux_h I__19565 (
            .O(N__84913),
            .I(N__84833));
    LocalMux I__19564 (
            .O(N__84906),
            .I(N__84824));
    Span4Mux_v I__19563 (
            .O(N__84903),
            .I(N__84824));
    LocalMux I__19562 (
            .O(N__84898),
            .I(N__84824));
    LocalMux I__19561 (
            .O(N__84893),
            .I(N__84824));
    Span4Mux_h I__19560 (
            .O(N__84890),
            .I(N__84819));
    Span12Mux_h I__19559 (
            .O(N__84881),
            .I(N__84816));
    Span4Mux_v I__19558 (
            .O(N__84878),
            .I(N__84811));
    Span4Mux_h I__19557 (
            .O(N__84869),
            .I(N__84811));
    Span12Mux_v I__19556 (
            .O(N__84864),
            .I(N__84806));
    Span12Mux_v I__19555 (
            .O(N__84861),
            .I(N__84806));
    Span4Mux_h I__19554 (
            .O(N__84850),
            .I(N__84803));
    Span4Mux_v I__19553 (
            .O(N__84845),
            .I(N__84794));
    Span4Mux_h I__19552 (
            .O(N__84838),
            .I(N__84794));
    Span4Mux_v I__19551 (
            .O(N__84833),
            .I(N__84794));
    Span4Mux_v I__19550 (
            .O(N__84824),
            .I(N__84794));
    InMux I__19549 (
            .O(N__84823),
            .I(N__84789));
    InMux I__19548 (
            .O(N__84822),
            .I(N__84789));
    Odrv4 I__19547 (
            .O(N__84819),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv12 I__19546 (
            .O(N__84816),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv4 I__19545 (
            .O(N__84811),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv12 I__19544 (
            .O(N__84806),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv4 I__19543 (
            .O(N__84803),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    Odrv4 I__19542 (
            .O(N__84794),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    LocalMux I__19541 (
            .O(N__84789),
            .I(FRAME_MATCHER_state_31_N_2976_2));
    CascadeMux I__19540 (
            .O(N__84774),
            .I(N__84770));
    CascadeMux I__19539 (
            .O(N__84773),
            .I(N__84766));
    InMux I__19538 (
            .O(N__84770),
            .I(N__84761));
    InMux I__19537 (
            .O(N__84769),
            .I(N__84761));
    InMux I__19536 (
            .O(N__84766),
            .I(N__84756));
    LocalMux I__19535 (
            .O(N__84761),
            .I(N__84753));
    InMux I__19534 (
            .O(N__84760),
            .I(N__84750));
    InMux I__19533 (
            .O(N__84759),
            .I(N__84747));
    LocalMux I__19532 (
            .O(N__84756),
            .I(N__84743));
    Span4Mux_v I__19531 (
            .O(N__84753),
            .I(N__84738));
    LocalMux I__19530 (
            .O(N__84750),
            .I(N__84738));
    LocalMux I__19529 (
            .O(N__84747),
            .I(N__84735));
    InMux I__19528 (
            .O(N__84746),
            .I(N__84732));
    Span4Mux_v I__19527 (
            .O(N__84743),
            .I(N__84727));
    Span4Mux_v I__19526 (
            .O(N__84738),
            .I(N__84727));
    Span4Mux_h I__19525 (
            .O(N__84735),
            .I(N__84724));
    LocalMux I__19524 (
            .O(N__84732),
            .I(encoder1_position_1));
    Odrv4 I__19523 (
            .O(N__84727),
            .I(encoder1_position_1));
    Odrv4 I__19522 (
            .O(N__84724),
            .I(encoder1_position_1));
    CascadeMux I__19521 (
            .O(N__84717),
            .I(N__84674));
    CascadeMux I__19520 (
            .O(N__84716),
            .I(N__84671));
    InMux I__19519 (
            .O(N__84715),
            .I(N__84662));
    InMux I__19518 (
            .O(N__84714),
            .I(N__84662));
    InMux I__19517 (
            .O(N__84713),
            .I(N__84662));
    InMux I__19516 (
            .O(N__84712),
            .I(N__84655));
    InMux I__19515 (
            .O(N__84711),
            .I(N__84655));
    InMux I__19514 (
            .O(N__84710),
            .I(N__84655));
    InMux I__19513 (
            .O(N__84709),
            .I(N__84652));
    InMux I__19512 (
            .O(N__84708),
            .I(N__84647));
    InMux I__19511 (
            .O(N__84707),
            .I(N__84647));
    InMux I__19510 (
            .O(N__84706),
            .I(N__84640));
    InMux I__19509 (
            .O(N__84705),
            .I(N__84640));
    InMux I__19508 (
            .O(N__84704),
            .I(N__84640));
    InMux I__19507 (
            .O(N__84703),
            .I(N__84634));
    InMux I__19506 (
            .O(N__84702),
            .I(N__84629));
    InMux I__19505 (
            .O(N__84701),
            .I(N__84629));
    CascadeMux I__19504 (
            .O(N__84700),
            .I(N__84620));
    InMux I__19503 (
            .O(N__84699),
            .I(N__84611));
    InMux I__19502 (
            .O(N__84698),
            .I(N__84606));
    InMux I__19501 (
            .O(N__84697),
            .I(N__84606));
    InMux I__19500 (
            .O(N__84696),
            .I(N__84597));
    InMux I__19499 (
            .O(N__84695),
            .I(N__84597));
    InMux I__19498 (
            .O(N__84694),
            .I(N__84597));
    InMux I__19497 (
            .O(N__84693),
            .I(N__84590));
    InMux I__19496 (
            .O(N__84692),
            .I(N__84590));
    InMux I__19495 (
            .O(N__84691),
            .I(N__84590));
    InMux I__19494 (
            .O(N__84690),
            .I(N__84581));
    InMux I__19493 (
            .O(N__84689),
            .I(N__84581));
    InMux I__19492 (
            .O(N__84688),
            .I(N__84581));
    InMux I__19491 (
            .O(N__84687),
            .I(N__84581));
    InMux I__19490 (
            .O(N__84686),
            .I(N__84574));
    InMux I__19489 (
            .O(N__84685),
            .I(N__84574));
    InMux I__19488 (
            .O(N__84684),
            .I(N__84574));
    InMux I__19487 (
            .O(N__84683),
            .I(N__84571));
    InMux I__19486 (
            .O(N__84682),
            .I(N__84562));
    InMux I__19485 (
            .O(N__84681),
            .I(N__84562));
    InMux I__19484 (
            .O(N__84680),
            .I(N__84562));
    InMux I__19483 (
            .O(N__84679),
            .I(N__84562));
    InMux I__19482 (
            .O(N__84678),
            .I(N__84555));
    InMux I__19481 (
            .O(N__84677),
            .I(N__84543));
    InMux I__19480 (
            .O(N__84674),
            .I(N__84543));
    InMux I__19479 (
            .O(N__84671),
            .I(N__84543));
    InMux I__19478 (
            .O(N__84670),
            .I(N__84543));
    InMux I__19477 (
            .O(N__84669),
            .I(N__84543));
    LocalMux I__19476 (
            .O(N__84662),
            .I(N__84538));
    LocalMux I__19475 (
            .O(N__84655),
            .I(N__84538));
    LocalMux I__19474 (
            .O(N__84652),
            .I(N__84535));
    LocalMux I__19473 (
            .O(N__84647),
            .I(N__84530));
    LocalMux I__19472 (
            .O(N__84640),
            .I(N__84530));
    InMux I__19471 (
            .O(N__84639),
            .I(N__84525));
    InMux I__19470 (
            .O(N__84638),
            .I(N__84525));
    InMux I__19469 (
            .O(N__84637),
            .I(N__84522));
    LocalMux I__19468 (
            .O(N__84634),
            .I(N__84519));
    LocalMux I__19467 (
            .O(N__84629),
            .I(N__84516));
    InMux I__19466 (
            .O(N__84628),
            .I(N__84509));
    InMux I__19465 (
            .O(N__84627),
            .I(N__84509));
    InMux I__19464 (
            .O(N__84626),
            .I(N__84509));
    InMux I__19463 (
            .O(N__84625),
            .I(N__84506));
    InMux I__19462 (
            .O(N__84624),
            .I(N__84501));
    InMux I__19461 (
            .O(N__84623),
            .I(N__84501));
    InMux I__19460 (
            .O(N__84620),
            .I(N__84498));
    InMux I__19459 (
            .O(N__84619),
            .I(N__84488));
    InMux I__19458 (
            .O(N__84618),
            .I(N__84488));
    InMux I__19457 (
            .O(N__84617),
            .I(N__84488));
    InMux I__19456 (
            .O(N__84616),
            .I(N__84488));
    InMux I__19455 (
            .O(N__84615),
            .I(N__84483));
    InMux I__19454 (
            .O(N__84614),
            .I(N__84483));
    LocalMux I__19453 (
            .O(N__84611),
            .I(N__84480));
    LocalMux I__19452 (
            .O(N__84606),
            .I(N__84477));
    InMux I__19451 (
            .O(N__84605),
            .I(N__84470));
    InMux I__19450 (
            .O(N__84604),
            .I(N__84470));
    LocalMux I__19449 (
            .O(N__84597),
            .I(N__84465));
    LocalMux I__19448 (
            .O(N__84590),
            .I(N__84465));
    LocalMux I__19447 (
            .O(N__84581),
            .I(N__84462));
    LocalMux I__19446 (
            .O(N__84574),
            .I(N__84455));
    LocalMux I__19445 (
            .O(N__84571),
            .I(N__84455));
    LocalMux I__19444 (
            .O(N__84562),
            .I(N__84455));
    CascadeMux I__19443 (
            .O(N__84561),
            .I(N__84451));
    InMux I__19442 (
            .O(N__84560),
            .I(N__84448));
    InMux I__19441 (
            .O(N__84559),
            .I(N__84445));
    InMux I__19440 (
            .O(N__84558),
            .I(N__84442));
    LocalMux I__19439 (
            .O(N__84555),
            .I(N__84439));
    InMux I__19438 (
            .O(N__84554),
            .I(N__84436));
    LocalMux I__19437 (
            .O(N__84543),
            .I(N__84427));
    Span4Mux_v I__19436 (
            .O(N__84538),
            .I(N__84427));
    Span4Mux_h I__19435 (
            .O(N__84535),
            .I(N__84427));
    Span4Mux_v I__19434 (
            .O(N__84530),
            .I(N__84427));
    LocalMux I__19433 (
            .O(N__84525),
            .I(N__84417));
    LocalMux I__19432 (
            .O(N__84522),
            .I(N__84417));
    Span4Mux_h I__19431 (
            .O(N__84519),
            .I(N__84414));
    Span4Mux_v I__19430 (
            .O(N__84516),
            .I(N__84411));
    LocalMux I__19429 (
            .O(N__84509),
            .I(N__84402));
    LocalMux I__19428 (
            .O(N__84506),
            .I(N__84402));
    LocalMux I__19427 (
            .O(N__84501),
            .I(N__84402));
    LocalMux I__19426 (
            .O(N__84498),
            .I(N__84402));
    InMux I__19425 (
            .O(N__84497),
            .I(N__84399));
    LocalMux I__19424 (
            .O(N__84488),
            .I(N__84390));
    LocalMux I__19423 (
            .O(N__84483),
            .I(N__84390));
    Span4Mux_v I__19422 (
            .O(N__84480),
            .I(N__84390));
    Span4Mux_h I__19421 (
            .O(N__84477),
            .I(N__84390));
    InMux I__19420 (
            .O(N__84476),
            .I(N__84385));
    InMux I__19419 (
            .O(N__84475),
            .I(N__84385));
    LocalMux I__19418 (
            .O(N__84470),
            .I(N__84380));
    Span4Mux_h I__19417 (
            .O(N__84465),
            .I(N__84380));
    Span4Mux_v I__19416 (
            .O(N__84462),
            .I(N__84375));
    Span4Mux_v I__19415 (
            .O(N__84455),
            .I(N__84375));
    InMux I__19414 (
            .O(N__84454),
            .I(N__84372));
    InMux I__19413 (
            .O(N__84451),
            .I(N__84369));
    LocalMux I__19412 (
            .O(N__84448),
            .I(N__84364));
    LocalMux I__19411 (
            .O(N__84445),
            .I(N__84364));
    LocalMux I__19410 (
            .O(N__84442),
            .I(N__84359));
    Sp12to4 I__19409 (
            .O(N__84439),
            .I(N__84359));
    LocalMux I__19408 (
            .O(N__84436),
            .I(N__84354));
    Span4Mux_h I__19407 (
            .O(N__84427),
            .I(N__84354));
    InMux I__19406 (
            .O(N__84426),
            .I(N__84347));
    InMux I__19405 (
            .O(N__84425),
            .I(N__84342));
    InMux I__19404 (
            .O(N__84424),
            .I(N__84342));
    InMux I__19403 (
            .O(N__84423),
            .I(N__84337));
    InMux I__19402 (
            .O(N__84422),
            .I(N__84337));
    Span4Mux_h I__19401 (
            .O(N__84417),
            .I(N__84328));
    Span4Mux_v I__19400 (
            .O(N__84414),
            .I(N__84328));
    Span4Mux_h I__19399 (
            .O(N__84411),
            .I(N__84328));
    Span4Mux_v I__19398 (
            .O(N__84402),
            .I(N__84328));
    LocalMux I__19397 (
            .O(N__84399),
            .I(N__84323));
    Span4Mux_h I__19396 (
            .O(N__84390),
            .I(N__84323));
    LocalMux I__19395 (
            .O(N__84385),
            .I(N__84316));
    Span4Mux_h I__19394 (
            .O(N__84380),
            .I(N__84316));
    Span4Mux_h I__19393 (
            .O(N__84375),
            .I(N__84316));
    LocalMux I__19392 (
            .O(N__84372),
            .I(N__84307));
    LocalMux I__19391 (
            .O(N__84369),
            .I(N__84307));
    Span12Mux_v I__19390 (
            .O(N__84364),
            .I(N__84307));
    Span12Mux_v I__19389 (
            .O(N__84359),
            .I(N__84307));
    Span4Mux_v I__19388 (
            .O(N__84354),
            .I(N__84304));
    InMux I__19387 (
            .O(N__84353),
            .I(N__84299));
    InMux I__19386 (
            .O(N__84352),
            .I(N__84299));
    InMux I__19385 (
            .O(N__84351),
            .I(N__84294));
    InMux I__19384 (
            .O(N__84350),
            .I(N__84294));
    LocalMux I__19383 (
            .O(N__84347),
            .I(data_out_frame_29__7__N_1482));
    LocalMux I__19382 (
            .O(N__84342),
            .I(data_out_frame_29__7__N_1482));
    LocalMux I__19381 (
            .O(N__84337),
            .I(data_out_frame_29__7__N_1482));
    Odrv4 I__19380 (
            .O(N__84328),
            .I(data_out_frame_29__7__N_1482));
    Odrv4 I__19379 (
            .O(N__84323),
            .I(data_out_frame_29__7__N_1482));
    Odrv4 I__19378 (
            .O(N__84316),
            .I(data_out_frame_29__7__N_1482));
    Odrv12 I__19377 (
            .O(N__84307),
            .I(data_out_frame_29__7__N_1482));
    Odrv4 I__19376 (
            .O(N__84304),
            .I(data_out_frame_29__7__N_1482));
    LocalMux I__19375 (
            .O(N__84299),
            .I(data_out_frame_29__7__N_1482));
    LocalMux I__19374 (
            .O(N__84294),
            .I(data_out_frame_29__7__N_1482));
    InMux I__19373 (
            .O(N__84273),
            .I(N__84270));
    LocalMux I__19372 (
            .O(N__84270),
            .I(N__84266));
    InMux I__19371 (
            .O(N__84269),
            .I(N__84263));
    Span12Mux_v I__19370 (
            .O(N__84266),
            .I(N__84260));
    LocalMux I__19369 (
            .O(N__84263),
            .I(data_out_frame_13_1));
    Odrv12 I__19368 (
            .O(N__84260),
            .I(data_out_frame_13_1));
    CascadeMux I__19367 (
            .O(N__84255),
            .I(N__84251));
    InMux I__19366 (
            .O(N__84254),
            .I(N__84248));
    InMux I__19365 (
            .O(N__84251),
            .I(N__84237));
    LocalMux I__19364 (
            .O(N__84248),
            .I(N__84227));
    InMux I__19363 (
            .O(N__84247),
            .I(N__84222));
    InMux I__19362 (
            .O(N__84246),
            .I(N__84222));
    InMux I__19361 (
            .O(N__84245),
            .I(N__84218));
    InMux I__19360 (
            .O(N__84244),
            .I(N__84214));
    InMux I__19359 (
            .O(N__84243),
            .I(N__84207));
    InMux I__19358 (
            .O(N__84242),
            .I(N__84207));
    InMux I__19357 (
            .O(N__84241),
            .I(N__84207));
    InMux I__19356 (
            .O(N__84240),
            .I(N__84204));
    LocalMux I__19355 (
            .O(N__84237),
            .I(N__84200));
    InMux I__19354 (
            .O(N__84236),
            .I(N__84197));
    InMux I__19353 (
            .O(N__84235),
            .I(N__84190));
    InMux I__19352 (
            .O(N__84234),
            .I(N__84190));
    InMux I__19351 (
            .O(N__84233),
            .I(N__84190));
    InMux I__19350 (
            .O(N__84232),
            .I(N__84187));
    InMux I__19349 (
            .O(N__84231),
            .I(N__84184));
    InMux I__19348 (
            .O(N__84230),
            .I(N__84181));
    Span4Mux_v I__19347 (
            .O(N__84227),
            .I(N__84175));
    LocalMux I__19346 (
            .O(N__84222),
            .I(N__84175));
    InMux I__19345 (
            .O(N__84221),
            .I(N__84172));
    LocalMux I__19344 (
            .O(N__84218),
            .I(N__84168));
    CascadeMux I__19343 (
            .O(N__84217),
            .I(N__84165));
    LocalMux I__19342 (
            .O(N__84214),
            .I(N__84162));
    LocalMux I__19341 (
            .O(N__84207),
            .I(N__84157));
    LocalMux I__19340 (
            .O(N__84204),
            .I(N__84157));
    InMux I__19339 (
            .O(N__84203),
            .I(N__84154));
    Span4Mux_v I__19338 (
            .O(N__84200),
            .I(N__84147));
    LocalMux I__19337 (
            .O(N__84197),
            .I(N__84147));
    LocalMux I__19336 (
            .O(N__84190),
            .I(N__84147));
    LocalMux I__19335 (
            .O(N__84187),
            .I(N__84143));
    LocalMux I__19334 (
            .O(N__84184),
            .I(N__84139));
    LocalMux I__19333 (
            .O(N__84181),
            .I(N__84136));
    InMux I__19332 (
            .O(N__84180),
            .I(N__84133));
    Span4Mux_h I__19331 (
            .O(N__84175),
            .I(N__84128));
    LocalMux I__19330 (
            .O(N__84172),
            .I(N__84128));
    InMux I__19329 (
            .O(N__84171),
            .I(N__84125));
    Span4Mux_v I__19328 (
            .O(N__84168),
            .I(N__84122));
    InMux I__19327 (
            .O(N__84165),
            .I(N__84118));
    Span4Mux_h I__19326 (
            .O(N__84162),
            .I(N__84111));
    Span4Mux_v I__19325 (
            .O(N__84157),
            .I(N__84111));
    LocalMux I__19324 (
            .O(N__84154),
            .I(N__84106));
    Span4Mux_v I__19323 (
            .O(N__84147),
            .I(N__84106));
    InMux I__19322 (
            .O(N__84146),
            .I(N__84103));
    Span4Mux_v I__19321 (
            .O(N__84143),
            .I(N__84100));
    InMux I__19320 (
            .O(N__84142),
            .I(N__84097));
    Span4Mux_h I__19319 (
            .O(N__84139),
            .I(N__84092));
    Span4Mux_v I__19318 (
            .O(N__84136),
            .I(N__84092));
    LocalMux I__19317 (
            .O(N__84133),
            .I(N__84089));
    Span4Mux_v I__19316 (
            .O(N__84128),
            .I(N__84084));
    LocalMux I__19315 (
            .O(N__84125),
            .I(N__84084));
    Span4Mux_h I__19314 (
            .O(N__84122),
            .I(N__84081));
    InMux I__19313 (
            .O(N__84121),
            .I(N__84078));
    LocalMux I__19312 (
            .O(N__84118),
            .I(N__84075));
    InMux I__19311 (
            .O(N__84117),
            .I(N__84072));
    InMux I__19310 (
            .O(N__84116),
            .I(N__84068));
    Sp12to4 I__19309 (
            .O(N__84111),
            .I(N__84057));
    Sp12to4 I__19308 (
            .O(N__84106),
            .I(N__84057));
    LocalMux I__19307 (
            .O(N__84103),
            .I(N__84057));
    Sp12to4 I__19306 (
            .O(N__84100),
            .I(N__84057));
    LocalMux I__19305 (
            .O(N__84097),
            .I(N__84057));
    Span4Mux_h I__19304 (
            .O(N__84092),
            .I(N__84050));
    Span4Mux_v I__19303 (
            .O(N__84089),
            .I(N__84050));
    Span4Mux_v I__19302 (
            .O(N__84084),
            .I(N__84050));
    Span4Mux_h I__19301 (
            .O(N__84081),
            .I(N__84047));
    LocalMux I__19300 (
            .O(N__84078),
            .I(N__84044));
    Span4Mux_h I__19299 (
            .O(N__84075),
            .I(N__84039));
    LocalMux I__19298 (
            .O(N__84072),
            .I(N__84039));
    InMux I__19297 (
            .O(N__84071),
            .I(N__84036));
    LocalMux I__19296 (
            .O(N__84068),
            .I(N__84033));
    Span12Mux_h I__19295 (
            .O(N__84057),
            .I(N__84026));
    Span4Mux_h I__19294 (
            .O(N__84050),
            .I(N__84023));
    Span4Mux_h I__19293 (
            .O(N__84047),
            .I(N__84018));
    Span4Mux_v I__19292 (
            .O(N__84044),
            .I(N__84018));
    Span4Mux_v I__19291 (
            .O(N__84039),
            .I(N__84013));
    LocalMux I__19290 (
            .O(N__84036),
            .I(N__84013));
    Span12Mux_v I__19289 (
            .O(N__84033),
            .I(N__84010));
    InMux I__19288 (
            .O(N__84032),
            .I(N__84007));
    InMux I__19287 (
            .O(N__84031),
            .I(N__84004));
    InMux I__19286 (
            .O(N__84030),
            .I(N__84001));
    InMux I__19285 (
            .O(N__84029),
            .I(N__83998));
    Odrv12 I__19284 (
            .O(N__84026),
            .I(rx_data_4));
    Odrv4 I__19283 (
            .O(N__84023),
            .I(rx_data_4));
    Odrv4 I__19282 (
            .O(N__84018),
            .I(rx_data_4));
    Odrv4 I__19281 (
            .O(N__84013),
            .I(rx_data_4));
    Odrv12 I__19280 (
            .O(N__84010),
            .I(rx_data_4));
    LocalMux I__19279 (
            .O(N__84007),
            .I(rx_data_4));
    LocalMux I__19278 (
            .O(N__84004),
            .I(rx_data_4));
    LocalMux I__19277 (
            .O(N__84001),
            .I(rx_data_4));
    LocalMux I__19276 (
            .O(N__83998),
            .I(rx_data_4));
    InMux I__19275 (
            .O(N__83979),
            .I(N__83944));
    InMux I__19274 (
            .O(N__83978),
            .I(N__83944));
    InMux I__19273 (
            .O(N__83977),
            .I(N__83944));
    InMux I__19272 (
            .O(N__83976),
            .I(N__83944));
    CascadeMux I__19271 (
            .O(N__83975),
            .I(N__83938));
    InMux I__19270 (
            .O(N__83974),
            .I(N__83933));
    InMux I__19269 (
            .O(N__83973),
            .I(N__83928));
    InMux I__19268 (
            .O(N__83972),
            .I(N__83928));
    InMux I__19267 (
            .O(N__83971),
            .I(N__83921));
    InMux I__19266 (
            .O(N__83970),
            .I(N__83921));
    InMux I__19265 (
            .O(N__83969),
            .I(N__83921));
    InMux I__19264 (
            .O(N__83968),
            .I(N__83915));
    InMux I__19263 (
            .O(N__83967),
            .I(N__83906));
    InMux I__19262 (
            .O(N__83966),
            .I(N__83899));
    InMux I__19261 (
            .O(N__83965),
            .I(N__83899));
    InMux I__19260 (
            .O(N__83964),
            .I(N__83899));
    InMux I__19259 (
            .O(N__83963),
            .I(N__83894));
    InMux I__19258 (
            .O(N__83962),
            .I(N__83894));
    InMux I__19257 (
            .O(N__83961),
            .I(N__83888));
    InMux I__19256 (
            .O(N__83960),
            .I(N__83885));
    InMux I__19255 (
            .O(N__83959),
            .I(N__83882));
    InMux I__19254 (
            .O(N__83958),
            .I(N__83877));
    InMux I__19253 (
            .O(N__83957),
            .I(N__83877));
    InMux I__19252 (
            .O(N__83956),
            .I(N__83872));
    InMux I__19251 (
            .O(N__83955),
            .I(N__83872));
    CascadeMux I__19250 (
            .O(N__83954),
            .I(N__83869));
    InMux I__19249 (
            .O(N__83953),
            .I(N__83864));
    LocalMux I__19248 (
            .O(N__83944),
            .I(N__83860));
    InMux I__19247 (
            .O(N__83943),
            .I(N__83855));
    InMux I__19246 (
            .O(N__83942),
            .I(N__83855));
    InMux I__19245 (
            .O(N__83941),
            .I(N__83852));
    InMux I__19244 (
            .O(N__83938),
            .I(N__83849));
    InMux I__19243 (
            .O(N__83937),
            .I(N__83844));
    InMux I__19242 (
            .O(N__83936),
            .I(N__83844));
    LocalMux I__19241 (
            .O(N__83933),
            .I(N__83841));
    LocalMux I__19240 (
            .O(N__83928),
            .I(N__83836));
    LocalMux I__19239 (
            .O(N__83921),
            .I(N__83836));
    InMux I__19238 (
            .O(N__83920),
            .I(N__83829));
    InMux I__19237 (
            .O(N__83919),
            .I(N__83829));
    InMux I__19236 (
            .O(N__83918),
            .I(N__83829));
    LocalMux I__19235 (
            .O(N__83915),
            .I(N__83826));
    InMux I__19234 (
            .O(N__83914),
            .I(N__83823));
    InMux I__19233 (
            .O(N__83913),
            .I(N__83820));
    InMux I__19232 (
            .O(N__83912),
            .I(N__83813));
    InMux I__19231 (
            .O(N__83911),
            .I(N__83813));
    InMux I__19230 (
            .O(N__83910),
            .I(N__83813));
    InMux I__19229 (
            .O(N__83909),
            .I(N__83804));
    LocalMux I__19228 (
            .O(N__83906),
            .I(N__83797));
    LocalMux I__19227 (
            .O(N__83899),
            .I(N__83797));
    LocalMux I__19226 (
            .O(N__83894),
            .I(N__83797));
    InMux I__19225 (
            .O(N__83893),
            .I(N__83794));
    InMux I__19224 (
            .O(N__83892),
            .I(N__83789));
    InMux I__19223 (
            .O(N__83891),
            .I(N__83789));
    LocalMux I__19222 (
            .O(N__83888),
            .I(N__83786));
    LocalMux I__19221 (
            .O(N__83885),
            .I(N__83781));
    LocalMux I__19220 (
            .O(N__83882),
            .I(N__83781));
    LocalMux I__19219 (
            .O(N__83877),
            .I(N__83776));
    LocalMux I__19218 (
            .O(N__83872),
            .I(N__83776));
    InMux I__19217 (
            .O(N__83869),
            .I(N__83773));
    InMux I__19216 (
            .O(N__83868),
            .I(N__83770));
    InMux I__19215 (
            .O(N__83867),
            .I(N__83767));
    LocalMux I__19214 (
            .O(N__83864),
            .I(N__83764));
    InMux I__19213 (
            .O(N__83863),
            .I(N__83761));
    Span4Mux_v I__19212 (
            .O(N__83860),
            .I(N__83756));
    LocalMux I__19211 (
            .O(N__83855),
            .I(N__83756));
    LocalMux I__19210 (
            .O(N__83852),
            .I(N__83751));
    LocalMux I__19209 (
            .O(N__83849),
            .I(N__83751));
    LocalMux I__19208 (
            .O(N__83844),
            .I(N__83744));
    Span4Mux_h I__19207 (
            .O(N__83841),
            .I(N__83744));
    Span4Mux_v I__19206 (
            .O(N__83836),
            .I(N__83744));
    LocalMux I__19205 (
            .O(N__83829),
            .I(N__83733));
    Span4Mux_h I__19204 (
            .O(N__83826),
            .I(N__83733));
    LocalMux I__19203 (
            .O(N__83823),
            .I(N__83733));
    LocalMux I__19202 (
            .O(N__83820),
            .I(N__83733));
    LocalMux I__19201 (
            .O(N__83813),
            .I(N__83733));
    InMux I__19200 (
            .O(N__83812),
            .I(N__83729));
    InMux I__19199 (
            .O(N__83811),
            .I(N__83724));
    InMux I__19198 (
            .O(N__83810),
            .I(N__83724));
    InMux I__19197 (
            .O(N__83809),
            .I(N__83717));
    InMux I__19196 (
            .O(N__83808),
            .I(N__83717));
    InMux I__19195 (
            .O(N__83807),
            .I(N__83717));
    LocalMux I__19194 (
            .O(N__83804),
            .I(N__83712));
    Span4Mux_v I__19193 (
            .O(N__83797),
            .I(N__83712));
    LocalMux I__19192 (
            .O(N__83794),
            .I(N__83707));
    LocalMux I__19191 (
            .O(N__83789),
            .I(N__83707));
    Span4Mux_v I__19190 (
            .O(N__83786),
            .I(N__83700));
    Span4Mux_v I__19189 (
            .O(N__83781),
            .I(N__83700));
    Span4Mux_v I__19188 (
            .O(N__83776),
            .I(N__83700));
    LocalMux I__19187 (
            .O(N__83773),
            .I(N__83695));
    LocalMux I__19186 (
            .O(N__83770),
            .I(N__83692));
    LocalMux I__19185 (
            .O(N__83767),
            .I(N__83689));
    Span4Mux_h I__19184 (
            .O(N__83764),
            .I(N__83676));
    LocalMux I__19183 (
            .O(N__83761),
            .I(N__83676));
    Span4Mux_v I__19182 (
            .O(N__83756),
            .I(N__83676));
    Span4Mux_v I__19181 (
            .O(N__83751),
            .I(N__83676));
    Span4Mux_h I__19180 (
            .O(N__83744),
            .I(N__83676));
    Span4Mux_v I__19179 (
            .O(N__83733),
            .I(N__83676));
    InMux I__19178 (
            .O(N__83732),
            .I(N__83673));
    LocalMux I__19177 (
            .O(N__83729),
            .I(N__83670));
    LocalMux I__19176 (
            .O(N__83724),
            .I(N__83665));
    LocalMux I__19175 (
            .O(N__83717),
            .I(N__83665));
    Span4Mux_h I__19174 (
            .O(N__83712),
            .I(N__83662));
    Span4Mux_v I__19173 (
            .O(N__83707),
            .I(N__83657));
    Span4Mux_h I__19172 (
            .O(N__83700),
            .I(N__83657));
    InMux I__19171 (
            .O(N__83699),
            .I(N__83654));
    InMux I__19170 (
            .O(N__83698),
            .I(N__83651));
    Span4Mux_v I__19169 (
            .O(N__83695),
            .I(N__83646));
    Span4Mux_v I__19168 (
            .O(N__83692),
            .I(N__83646));
    Span12Mux_s11_v I__19167 (
            .O(N__83689),
            .I(N__83641));
    Sp12to4 I__19166 (
            .O(N__83676),
            .I(N__83641));
    LocalMux I__19165 (
            .O(N__83673),
            .I(N__83630));
    Span4Mux_v I__19164 (
            .O(N__83670),
            .I(N__83630));
    Span4Mux_v I__19163 (
            .O(N__83665),
            .I(N__83630));
    Span4Mux_h I__19162 (
            .O(N__83662),
            .I(N__83630));
    Span4Mux_h I__19161 (
            .O(N__83657),
            .I(N__83630));
    LocalMux I__19160 (
            .O(N__83654),
            .I(\c0.n33249 ));
    LocalMux I__19159 (
            .O(N__83651),
            .I(\c0.n33249 ));
    Odrv4 I__19158 (
            .O(N__83646),
            .I(\c0.n33249 ));
    Odrv12 I__19157 (
            .O(N__83641),
            .I(\c0.n33249 ));
    Odrv4 I__19156 (
            .O(N__83630),
            .I(\c0.n33249 ));
    InMux I__19155 (
            .O(N__83619),
            .I(N__83613));
    InMux I__19154 (
            .O(N__83618),
            .I(N__83610));
    InMux I__19153 (
            .O(N__83617),
            .I(N__83605));
    InMux I__19152 (
            .O(N__83616),
            .I(N__83605));
    LocalMux I__19151 (
            .O(N__83613),
            .I(N__83602));
    LocalMux I__19150 (
            .O(N__83610),
            .I(N__83599));
    LocalMux I__19149 (
            .O(N__83605),
            .I(N__83596));
    Span4Mux_v I__19148 (
            .O(N__83602),
            .I(N__83591));
    Span4Mux_h I__19147 (
            .O(N__83599),
            .I(N__83586));
    Span4Mux_v I__19146 (
            .O(N__83596),
            .I(N__83586));
    CascadeMux I__19145 (
            .O(N__83595),
            .I(N__83583));
    InMux I__19144 (
            .O(N__83594),
            .I(N__83580));
    Span4Mux_h I__19143 (
            .O(N__83591),
            .I(N__83577));
    Span4Mux_h I__19142 (
            .O(N__83586),
            .I(N__83574));
    InMux I__19141 (
            .O(N__83583),
            .I(N__83571));
    LocalMux I__19140 (
            .O(N__83580),
            .I(N__83568));
    Span4Mux_h I__19139 (
            .O(N__83577),
            .I(N__83565));
    Span4Mux_h I__19138 (
            .O(N__83574),
            .I(N__83562));
    LocalMux I__19137 (
            .O(N__83571),
            .I(data_in_frame_1_4));
    Odrv4 I__19136 (
            .O(N__83568),
            .I(data_in_frame_1_4));
    Odrv4 I__19135 (
            .O(N__83565),
            .I(data_in_frame_1_4));
    Odrv4 I__19134 (
            .O(N__83562),
            .I(data_in_frame_1_4));
    InMux I__19133 (
            .O(N__83553),
            .I(N__83550));
    LocalMux I__19132 (
            .O(N__83550),
            .I(N__83547));
    Span4Mux_v I__19131 (
            .O(N__83547),
            .I(N__83544));
    Odrv4 I__19130 (
            .O(N__83544),
            .I(\c0.n26_adj_4654 ));
    CascadeMux I__19129 (
            .O(N__83541),
            .I(N__83538));
    InMux I__19128 (
            .O(N__83538),
            .I(N__83535));
    LocalMux I__19127 (
            .O(N__83535),
            .I(N__83530));
    InMux I__19126 (
            .O(N__83534),
            .I(N__83526));
    InMux I__19125 (
            .O(N__83533),
            .I(N__83523));
    Span4Mux_v I__19124 (
            .O(N__83530),
            .I(N__83519));
    CascadeMux I__19123 (
            .O(N__83529),
            .I(N__83516));
    LocalMux I__19122 (
            .O(N__83526),
            .I(N__83513));
    LocalMux I__19121 (
            .O(N__83523),
            .I(N__83510));
    InMux I__19120 (
            .O(N__83522),
            .I(N__83507));
    Span4Mux_h I__19119 (
            .O(N__83519),
            .I(N__83504));
    InMux I__19118 (
            .O(N__83516),
            .I(N__83501));
    Span4Mux_v I__19117 (
            .O(N__83513),
            .I(N__83498));
    Span4Mux_v I__19116 (
            .O(N__83510),
            .I(N__83495));
    LocalMux I__19115 (
            .O(N__83507),
            .I(encoder1_position_3));
    Odrv4 I__19114 (
            .O(N__83504),
            .I(encoder1_position_3));
    LocalMux I__19113 (
            .O(N__83501),
            .I(encoder1_position_3));
    Odrv4 I__19112 (
            .O(N__83498),
            .I(encoder1_position_3));
    Odrv4 I__19111 (
            .O(N__83495),
            .I(encoder1_position_3));
    CascadeMux I__19110 (
            .O(N__83484),
            .I(N__83478));
    InMux I__19109 (
            .O(N__83483),
            .I(N__83474));
    InMux I__19108 (
            .O(N__83482),
            .I(N__83471));
    InMux I__19107 (
            .O(N__83481),
            .I(N__83468));
    InMux I__19106 (
            .O(N__83478),
            .I(N__83463));
    InMux I__19105 (
            .O(N__83477),
            .I(N__83460));
    LocalMux I__19104 (
            .O(N__83474),
            .I(N__83455));
    LocalMux I__19103 (
            .O(N__83471),
            .I(N__83455));
    LocalMux I__19102 (
            .O(N__83468),
            .I(N__83452));
    InMux I__19101 (
            .O(N__83467),
            .I(N__83449));
    InMux I__19100 (
            .O(N__83466),
            .I(N__83446));
    LocalMux I__19099 (
            .O(N__83463),
            .I(N__83443));
    LocalMux I__19098 (
            .O(N__83460),
            .I(N__83438));
    Span4Mux_h I__19097 (
            .O(N__83455),
            .I(N__83438));
    Span4Mux_h I__19096 (
            .O(N__83452),
            .I(N__83433));
    LocalMux I__19095 (
            .O(N__83449),
            .I(N__83433));
    LocalMux I__19094 (
            .O(N__83446),
            .I(encoder1_position_11));
    Odrv12 I__19093 (
            .O(N__83443),
            .I(encoder1_position_11));
    Odrv4 I__19092 (
            .O(N__83438),
            .I(encoder1_position_11));
    Odrv4 I__19091 (
            .O(N__83433),
            .I(encoder1_position_11));
    InMux I__19090 (
            .O(N__83424),
            .I(N__83418));
    InMux I__19089 (
            .O(N__83423),
            .I(N__83415));
    InMux I__19088 (
            .O(N__83422),
            .I(N__83412));
    InMux I__19087 (
            .O(N__83421),
            .I(N__83409));
    LocalMux I__19086 (
            .O(N__83418),
            .I(N__83404));
    LocalMux I__19085 (
            .O(N__83415),
            .I(N__83404));
    LocalMux I__19084 (
            .O(N__83412),
            .I(N__83401));
    LocalMux I__19083 (
            .O(N__83409),
            .I(N__83398));
    Span4Mux_h I__19082 (
            .O(N__83404),
            .I(N__83395));
    Span4Mux_h I__19081 (
            .O(N__83401),
            .I(N__83392));
    Odrv12 I__19080 (
            .O(N__83398),
            .I(\c0.n31673 ));
    Odrv4 I__19079 (
            .O(N__83395),
            .I(\c0.n31673 ));
    Odrv4 I__19078 (
            .O(N__83392),
            .I(\c0.n31673 ));
    InMux I__19077 (
            .O(N__83385),
            .I(N__83382));
    LocalMux I__19076 (
            .O(N__83382),
            .I(\c0.n33425 ));
    CascadeMux I__19075 (
            .O(N__83379),
            .I(\c0.data_out_frame_29__7__N_658_cascade_ ));
    InMux I__19074 (
            .O(N__83376),
            .I(N__83373));
    LocalMux I__19073 (
            .O(N__83373),
            .I(N__83370));
    Odrv12 I__19072 (
            .O(N__83370),
            .I(\quad_counter1.n33_adj_4466 ));
    InMux I__19071 (
            .O(N__83367),
            .I(N__83364));
    LocalMux I__19070 (
            .O(N__83364),
            .I(N__83361));
    Span4Mux_v I__19069 (
            .O(N__83361),
            .I(N__83358));
    Span4Mux_h I__19068 (
            .O(N__83358),
            .I(N__83355));
    Odrv4 I__19067 (
            .O(N__83355),
            .I(\c0.n35821 ));
    InMux I__19066 (
            .O(N__83352),
            .I(N__83349));
    LocalMux I__19065 (
            .O(N__83349),
            .I(N__83346));
    Odrv12 I__19064 (
            .O(N__83346),
            .I(n35823));
    InMux I__19063 (
            .O(N__83343),
            .I(N__83339));
    InMux I__19062 (
            .O(N__83342),
            .I(N__83336));
    LocalMux I__19061 (
            .O(N__83339),
            .I(data_out_frame_28_3));
    LocalMux I__19060 (
            .O(N__83336),
            .I(data_out_frame_28_3));
    InMux I__19059 (
            .O(N__83331),
            .I(N__83327));
    InMux I__19058 (
            .O(N__83330),
            .I(N__83324));
    LocalMux I__19057 (
            .O(N__83327),
            .I(N__83321));
    LocalMux I__19056 (
            .O(N__83324),
            .I(N__83317));
    Sp12to4 I__19055 (
            .O(N__83321),
            .I(N__83313));
    InMux I__19054 (
            .O(N__83320),
            .I(N__83310));
    Span4Mux_h I__19053 (
            .O(N__83317),
            .I(N__83306));
    InMux I__19052 (
            .O(N__83316),
            .I(N__83303));
    Span12Mux_h I__19051 (
            .O(N__83313),
            .I(N__83300));
    LocalMux I__19050 (
            .O(N__83310),
            .I(N__83297));
    InMux I__19049 (
            .O(N__83309),
            .I(N__83294));
    Span4Mux_v I__19048 (
            .O(N__83306),
            .I(N__83291));
    LocalMux I__19047 (
            .O(N__83303),
            .I(encoder0_position_2));
    Odrv12 I__19046 (
            .O(N__83300),
            .I(encoder0_position_2));
    Odrv12 I__19045 (
            .O(N__83297),
            .I(encoder0_position_2));
    LocalMux I__19044 (
            .O(N__83294),
            .I(encoder0_position_2));
    Odrv4 I__19043 (
            .O(N__83291),
            .I(encoder0_position_2));
    InMux I__19042 (
            .O(N__83280),
            .I(N__83276));
    InMux I__19041 (
            .O(N__83279),
            .I(N__83273));
    LocalMux I__19040 (
            .O(N__83276),
            .I(N__83268));
    LocalMux I__19039 (
            .O(N__83273),
            .I(N__83264));
    InMux I__19038 (
            .O(N__83272),
            .I(N__83261));
    InMux I__19037 (
            .O(N__83271),
            .I(N__83258));
    Span4Mux_v I__19036 (
            .O(N__83268),
            .I(N__83255));
    InMux I__19035 (
            .O(N__83267),
            .I(N__83252));
    Span4Mux_h I__19034 (
            .O(N__83264),
            .I(N__83249));
    LocalMux I__19033 (
            .O(N__83261),
            .I(N__83244));
    LocalMux I__19032 (
            .O(N__83258),
            .I(N__83244));
    Span4Mux_v I__19031 (
            .O(N__83255),
            .I(N__83241));
    LocalMux I__19030 (
            .O(N__83252),
            .I(encoder0_position_17));
    Odrv4 I__19029 (
            .O(N__83249),
            .I(encoder0_position_17));
    Odrv12 I__19028 (
            .O(N__83244),
            .I(encoder0_position_17));
    Odrv4 I__19027 (
            .O(N__83241),
            .I(encoder0_position_17));
    CascadeMux I__19026 (
            .O(N__83232),
            .I(N__83229));
    InMux I__19025 (
            .O(N__83229),
            .I(N__83225));
    CascadeMux I__19024 (
            .O(N__83228),
            .I(N__83221));
    LocalMux I__19023 (
            .O(N__83225),
            .I(N__83217));
    CascadeMux I__19022 (
            .O(N__83224),
            .I(N__83214));
    InMux I__19021 (
            .O(N__83221),
            .I(N__83211));
    InMux I__19020 (
            .O(N__83220),
            .I(N__83208));
    Span12Mux_h I__19019 (
            .O(N__83217),
            .I(N__83205));
    InMux I__19018 (
            .O(N__83214),
            .I(N__83202));
    LocalMux I__19017 (
            .O(N__83211),
            .I(N__83199));
    LocalMux I__19016 (
            .O(N__83208),
            .I(encoder1_position_19));
    Odrv12 I__19015 (
            .O(N__83205),
            .I(encoder1_position_19));
    LocalMux I__19014 (
            .O(N__83202),
            .I(encoder1_position_19));
    Odrv12 I__19013 (
            .O(N__83199),
            .I(encoder1_position_19));
    CascadeMux I__19012 (
            .O(N__83190),
            .I(N__83187));
    InMux I__19011 (
            .O(N__83187),
            .I(N__83183));
    CascadeMux I__19010 (
            .O(N__83186),
            .I(N__83180));
    LocalMux I__19009 (
            .O(N__83183),
            .I(N__83175));
    InMux I__19008 (
            .O(N__83180),
            .I(N__83170));
    InMux I__19007 (
            .O(N__83179),
            .I(N__83170));
    InMux I__19006 (
            .O(N__83178),
            .I(N__83166));
    Span4Mux_v I__19005 (
            .O(N__83175),
            .I(N__83161));
    LocalMux I__19004 (
            .O(N__83170),
            .I(N__83161));
    InMux I__19003 (
            .O(N__83169),
            .I(N__83158));
    LocalMux I__19002 (
            .O(N__83166),
            .I(control_mode_0));
    Odrv4 I__19001 (
            .O(N__83161),
            .I(control_mode_0));
    LocalMux I__19000 (
            .O(N__83158),
            .I(control_mode_0));
    CascadeMux I__18999 (
            .O(N__83151),
            .I(N__83148));
    InMux I__18998 (
            .O(N__83148),
            .I(N__83142));
    InMux I__18997 (
            .O(N__83147),
            .I(N__83142));
    LocalMux I__18996 (
            .O(N__83142),
            .I(\c0.n35113 ));
    InMux I__18995 (
            .O(N__83139),
            .I(N__83132));
    InMux I__18994 (
            .O(N__83138),
            .I(N__83132));
    CascadeMux I__18993 (
            .O(N__83137),
            .I(N__83129));
    LocalMux I__18992 (
            .O(N__83132),
            .I(N__83124));
    InMux I__18991 (
            .O(N__83129),
            .I(N__83121));
    InMux I__18990 (
            .O(N__83128),
            .I(N__83118));
    InMux I__18989 (
            .O(N__83127),
            .I(N__83114));
    Span4Mux_v I__18988 (
            .O(N__83124),
            .I(N__83111));
    LocalMux I__18987 (
            .O(N__83121),
            .I(N__83106));
    LocalMux I__18986 (
            .O(N__83118),
            .I(N__83106));
    InMux I__18985 (
            .O(N__83117),
            .I(N__83103));
    LocalMux I__18984 (
            .O(N__83114),
            .I(N__83100));
    Span4Mux_h I__18983 (
            .O(N__83111),
            .I(N__83097));
    Span4Mux_v I__18982 (
            .O(N__83106),
            .I(N__83094));
    LocalMux I__18981 (
            .O(N__83103),
            .I(encoder1_position_10));
    Odrv4 I__18980 (
            .O(N__83100),
            .I(encoder1_position_10));
    Odrv4 I__18979 (
            .O(N__83097),
            .I(encoder1_position_10));
    Odrv4 I__18978 (
            .O(N__83094),
            .I(encoder1_position_10));
    InMux I__18977 (
            .O(N__83085),
            .I(N__83082));
    LocalMux I__18976 (
            .O(N__83082),
            .I(N__83078));
    InMux I__18975 (
            .O(N__83081),
            .I(N__83075));
    Span4Mux_v I__18974 (
            .O(N__83078),
            .I(N__83070));
    LocalMux I__18973 (
            .O(N__83075),
            .I(N__83070));
    Odrv4 I__18972 (
            .O(N__83070),
            .I(\c0.n33755 ));
    CascadeMux I__18971 (
            .O(N__83067),
            .I(\c0.n31446_cascade_ ));
    InMux I__18970 (
            .O(N__83064),
            .I(N__83061));
    LocalMux I__18969 (
            .O(N__83061),
            .I(N__83055));
    CascadeMux I__18968 (
            .O(N__83060),
            .I(N__83051));
    InMux I__18967 (
            .O(N__83059),
            .I(N__83048));
    InMux I__18966 (
            .O(N__83058),
            .I(N__83045));
    Span4Mux_v I__18965 (
            .O(N__83055),
            .I(N__83042));
    InMux I__18964 (
            .O(N__83054),
            .I(N__83038));
    InMux I__18963 (
            .O(N__83051),
            .I(N__83035));
    LocalMux I__18962 (
            .O(N__83048),
            .I(N__83032));
    LocalMux I__18961 (
            .O(N__83045),
            .I(N__83027));
    Span4Mux_h I__18960 (
            .O(N__83042),
            .I(N__83027));
    InMux I__18959 (
            .O(N__83041),
            .I(N__83024));
    LocalMux I__18958 (
            .O(N__83038),
            .I(encoder1_position_9));
    LocalMux I__18957 (
            .O(N__83035),
            .I(encoder1_position_9));
    Odrv12 I__18956 (
            .O(N__83032),
            .I(encoder1_position_9));
    Odrv4 I__18955 (
            .O(N__83027),
            .I(encoder1_position_9));
    LocalMux I__18954 (
            .O(N__83024),
            .I(encoder1_position_9));
    InMux I__18953 (
            .O(N__83013),
            .I(N__83009));
    InMux I__18952 (
            .O(N__83012),
            .I(N__83006));
    LocalMux I__18951 (
            .O(N__83009),
            .I(N__83001));
    LocalMux I__18950 (
            .O(N__83006),
            .I(N__83001));
    Span4Mux_v I__18949 (
            .O(N__83001),
            .I(N__82997));
    InMux I__18948 (
            .O(N__83000),
            .I(N__82994));
    Odrv4 I__18947 (
            .O(N__82997),
            .I(\quad_counter1.n3304 ));
    LocalMux I__18946 (
            .O(N__82994),
            .I(\quad_counter1.n3304 ));
    InMux I__18945 (
            .O(N__82989),
            .I(bfn_22_15_0_));
    InMux I__18944 (
            .O(N__82986),
            .I(N__82982));
    InMux I__18943 (
            .O(N__82985),
            .I(N__82979));
    LocalMux I__18942 (
            .O(N__82982),
            .I(N__82973));
    LocalMux I__18941 (
            .O(N__82979),
            .I(N__82973));
    CascadeMux I__18940 (
            .O(N__82978),
            .I(N__82970));
    Span4Mux_h I__18939 (
            .O(N__82973),
            .I(N__82967));
    InMux I__18938 (
            .O(N__82970),
            .I(N__82964));
    Odrv4 I__18937 (
            .O(N__82967),
            .I(\quad_counter1.n3303 ));
    LocalMux I__18936 (
            .O(N__82964),
            .I(\quad_counter1.n3303 ));
    InMux I__18935 (
            .O(N__82959),
            .I(\quad_counter1.n30670 ));
    InMux I__18934 (
            .O(N__82956),
            .I(N__82952));
    InMux I__18933 (
            .O(N__82955),
            .I(N__82949));
    LocalMux I__18932 (
            .O(N__82952),
            .I(N__82944));
    LocalMux I__18931 (
            .O(N__82949),
            .I(N__82944));
    Span4Mux_h I__18930 (
            .O(N__82944),
            .I(N__82940));
    InMux I__18929 (
            .O(N__82943),
            .I(N__82937));
    Odrv4 I__18928 (
            .O(N__82940),
            .I(\quad_counter1.n3302 ));
    LocalMux I__18927 (
            .O(N__82937),
            .I(\quad_counter1.n3302 ));
    InMux I__18926 (
            .O(N__82932),
            .I(\quad_counter1.n30671 ));
    InMux I__18925 (
            .O(N__82929),
            .I(N__82925));
    InMux I__18924 (
            .O(N__82928),
            .I(N__82922));
    LocalMux I__18923 (
            .O(N__82925),
            .I(N__82917));
    LocalMux I__18922 (
            .O(N__82922),
            .I(N__82917));
    Span4Mux_v I__18921 (
            .O(N__82917),
            .I(N__82913));
    InMux I__18920 (
            .O(N__82916),
            .I(N__82910));
    Odrv4 I__18919 (
            .O(N__82913),
            .I(\quad_counter1.n3301 ));
    LocalMux I__18918 (
            .O(N__82910),
            .I(\quad_counter1.n3301 ));
    InMux I__18917 (
            .O(N__82905),
            .I(\quad_counter1.n30672 ));
    InMux I__18916 (
            .O(N__82902),
            .I(N__82898));
    InMux I__18915 (
            .O(N__82901),
            .I(N__82895));
    LocalMux I__18914 (
            .O(N__82898),
            .I(N__82890));
    LocalMux I__18913 (
            .O(N__82895),
            .I(N__82890));
    Span4Mux_v I__18912 (
            .O(N__82890),
            .I(N__82886));
    InMux I__18911 (
            .O(N__82889),
            .I(N__82883));
    Odrv4 I__18910 (
            .O(N__82886),
            .I(\quad_counter1.n3300 ));
    LocalMux I__18909 (
            .O(N__82883),
            .I(\quad_counter1.n3300 ));
    InMux I__18908 (
            .O(N__82878),
            .I(\quad_counter1.n30673 ));
    InMux I__18907 (
            .O(N__82875),
            .I(N__82871));
    InMux I__18906 (
            .O(N__82874),
            .I(N__82868));
    LocalMux I__18905 (
            .O(N__82871),
            .I(N__82863));
    LocalMux I__18904 (
            .O(N__82868),
            .I(N__82863));
    Span4Mux_h I__18903 (
            .O(N__82863),
            .I(N__82859));
    InMux I__18902 (
            .O(N__82862),
            .I(N__82856));
    Odrv4 I__18901 (
            .O(N__82859),
            .I(\quad_counter1.n3299 ));
    LocalMux I__18900 (
            .O(N__82856),
            .I(\quad_counter1.n3299 ));
    CascadeMux I__18899 (
            .O(N__82851),
            .I(N__82833));
    CascadeMux I__18898 (
            .O(N__82850),
            .I(N__82830));
    CascadeMux I__18897 (
            .O(N__82849),
            .I(N__82827));
    CascadeMux I__18896 (
            .O(N__82848),
            .I(N__82824));
    CascadeMux I__18895 (
            .O(N__82847),
            .I(N__82821));
    CascadeMux I__18894 (
            .O(N__82846),
            .I(N__82818));
    CascadeMux I__18893 (
            .O(N__82845),
            .I(N__82815));
    CascadeMux I__18892 (
            .O(N__82844),
            .I(N__82812));
    CascadeMux I__18891 (
            .O(N__82843),
            .I(N__82809));
    CascadeMux I__18890 (
            .O(N__82842),
            .I(N__82806));
    CascadeMux I__18889 (
            .O(N__82841),
            .I(N__82803));
    CascadeMux I__18888 (
            .O(N__82840),
            .I(N__82800));
    CascadeMux I__18887 (
            .O(N__82839),
            .I(N__82797));
    CascadeMux I__18886 (
            .O(N__82838),
            .I(N__82794));
    CascadeMux I__18885 (
            .O(N__82837),
            .I(N__82791));
    CascadeMux I__18884 (
            .O(N__82836),
            .I(N__82788));
    InMux I__18883 (
            .O(N__82833),
            .I(N__82781));
    InMux I__18882 (
            .O(N__82830),
            .I(N__82781));
    InMux I__18881 (
            .O(N__82827),
            .I(N__82781));
    InMux I__18880 (
            .O(N__82824),
            .I(N__82774));
    InMux I__18879 (
            .O(N__82821),
            .I(N__82774));
    InMux I__18878 (
            .O(N__82818),
            .I(N__82774));
    InMux I__18877 (
            .O(N__82815),
            .I(N__82765));
    InMux I__18876 (
            .O(N__82812),
            .I(N__82765));
    InMux I__18875 (
            .O(N__82809),
            .I(N__82765));
    InMux I__18874 (
            .O(N__82806),
            .I(N__82765));
    InMux I__18873 (
            .O(N__82803),
            .I(N__82756));
    InMux I__18872 (
            .O(N__82800),
            .I(N__82756));
    InMux I__18871 (
            .O(N__82797),
            .I(N__82756));
    InMux I__18870 (
            .O(N__82794),
            .I(N__82756));
    InMux I__18869 (
            .O(N__82791),
            .I(N__82751));
    InMux I__18868 (
            .O(N__82788),
            .I(N__82751));
    LocalMux I__18867 (
            .O(N__82781),
            .I(\quad_counter1.n3332 ));
    LocalMux I__18866 (
            .O(N__82774),
            .I(\quad_counter1.n3332 ));
    LocalMux I__18865 (
            .O(N__82765),
            .I(\quad_counter1.n3332 ));
    LocalMux I__18864 (
            .O(N__82756),
            .I(\quad_counter1.n3332 ));
    LocalMux I__18863 (
            .O(N__82751),
            .I(\quad_counter1.n3332 ));
    InMux I__18862 (
            .O(N__82740),
            .I(\quad_counter1.n30674 ));
    InMux I__18861 (
            .O(N__82737),
            .I(N__82734));
    LocalMux I__18860 (
            .O(N__82734),
            .I(N__82731));
    Odrv4 I__18859 (
            .O(N__82731),
            .I(\quad_counter1.n35050 ));
    InMux I__18858 (
            .O(N__82728),
            .I(N__82724));
    InMux I__18857 (
            .O(N__82727),
            .I(N__82721));
    LocalMux I__18856 (
            .O(N__82724),
            .I(N__82715));
    LocalMux I__18855 (
            .O(N__82721),
            .I(N__82715));
    InMux I__18854 (
            .O(N__82720),
            .I(N__82712));
    Span4Mux_h I__18853 (
            .O(N__82715),
            .I(N__82707));
    LocalMux I__18852 (
            .O(N__82712),
            .I(N__82707));
    Odrv4 I__18851 (
            .O(N__82707),
            .I(\quad_counter1.n3313 ));
    InMux I__18850 (
            .O(N__82704),
            .I(\quad_counter1.n30660 ));
    InMux I__18849 (
            .O(N__82701),
            .I(N__82697));
    InMux I__18848 (
            .O(N__82700),
            .I(N__82694));
    LocalMux I__18847 (
            .O(N__82697),
            .I(N__82688));
    LocalMux I__18846 (
            .O(N__82694),
            .I(N__82688));
    InMux I__18845 (
            .O(N__82693),
            .I(N__82685));
    Span4Mux_h I__18844 (
            .O(N__82688),
            .I(N__82680));
    LocalMux I__18843 (
            .O(N__82685),
            .I(N__82680));
    Odrv4 I__18842 (
            .O(N__82680),
            .I(\quad_counter1.n3312 ));
    InMux I__18841 (
            .O(N__82677),
            .I(bfn_22_14_0_));
    InMux I__18840 (
            .O(N__82674),
            .I(N__82670));
    InMux I__18839 (
            .O(N__82673),
            .I(N__82667));
    LocalMux I__18838 (
            .O(N__82670),
            .I(N__82661));
    LocalMux I__18837 (
            .O(N__82667),
            .I(N__82661));
    CascadeMux I__18836 (
            .O(N__82666),
            .I(N__82658));
    Span4Mux_v I__18835 (
            .O(N__82661),
            .I(N__82655));
    InMux I__18834 (
            .O(N__82658),
            .I(N__82652));
    Odrv4 I__18833 (
            .O(N__82655),
            .I(\quad_counter1.n3311 ));
    LocalMux I__18832 (
            .O(N__82652),
            .I(\quad_counter1.n3311 ));
    InMux I__18831 (
            .O(N__82647),
            .I(\quad_counter1.n30662 ));
    InMux I__18830 (
            .O(N__82644),
            .I(N__82640));
    InMux I__18829 (
            .O(N__82643),
            .I(N__82637));
    LocalMux I__18828 (
            .O(N__82640),
            .I(N__82632));
    LocalMux I__18827 (
            .O(N__82637),
            .I(N__82632));
    Span4Mux_v I__18826 (
            .O(N__82632),
            .I(N__82628));
    InMux I__18825 (
            .O(N__82631),
            .I(N__82625));
    Odrv4 I__18824 (
            .O(N__82628),
            .I(\quad_counter1.n3310 ));
    LocalMux I__18823 (
            .O(N__82625),
            .I(\quad_counter1.n3310 ));
    InMux I__18822 (
            .O(N__82620),
            .I(\quad_counter1.n30663 ));
    InMux I__18821 (
            .O(N__82617),
            .I(N__82613));
    InMux I__18820 (
            .O(N__82616),
            .I(N__82610));
    LocalMux I__18819 (
            .O(N__82613),
            .I(N__82604));
    LocalMux I__18818 (
            .O(N__82610),
            .I(N__82604));
    CascadeMux I__18817 (
            .O(N__82609),
            .I(N__82601));
    Span4Mux_v I__18816 (
            .O(N__82604),
            .I(N__82598));
    InMux I__18815 (
            .O(N__82601),
            .I(N__82595));
    Odrv4 I__18814 (
            .O(N__82598),
            .I(\quad_counter1.n3309 ));
    LocalMux I__18813 (
            .O(N__82595),
            .I(\quad_counter1.n3309 ));
    InMux I__18812 (
            .O(N__82590),
            .I(\quad_counter1.n30664 ));
    InMux I__18811 (
            .O(N__82587),
            .I(N__82583));
    InMux I__18810 (
            .O(N__82586),
            .I(N__82580));
    LocalMux I__18809 (
            .O(N__82583),
            .I(N__82575));
    LocalMux I__18808 (
            .O(N__82580),
            .I(N__82575));
    Span4Mux_v I__18807 (
            .O(N__82575),
            .I(N__82571));
    InMux I__18806 (
            .O(N__82574),
            .I(N__82568));
    Odrv4 I__18805 (
            .O(N__82571),
            .I(\quad_counter1.n3308 ));
    LocalMux I__18804 (
            .O(N__82568),
            .I(\quad_counter1.n3308 ));
    InMux I__18803 (
            .O(N__82563),
            .I(\quad_counter1.n30665 ));
    InMux I__18802 (
            .O(N__82560),
            .I(N__82556));
    InMux I__18801 (
            .O(N__82559),
            .I(N__82553));
    LocalMux I__18800 (
            .O(N__82556),
            .I(N__82547));
    LocalMux I__18799 (
            .O(N__82553),
            .I(N__82547));
    CascadeMux I__18798 (
            .O(N__82552),
            .I(N__82544));
    Span4Mux_h I__18797 (
            .O(N__82547),
            .I(N__82541));
    InMux I__18796 (
            .O(N__82544),
            .I(N__82538));
    Odrv4 I__18795 (
            .O(N__82541),
            .I(\quad_counter1.n3307 ));
    LocalMux I__18794 (
            .O(N__82538),
            .I(\quad_counter1.n3307 ));
    InMux I__18793 (
            .O(N__82533),
            .I(\quad_counter1.n30666 ));
    InMux I__18792 (
            .O(N__82530),
            .I(N__82526));
    InMux I__18791 (
            .O(N__82529),
            .I(N__82523));
    LocalMux I__18790 (
            .O(N__82526),
            .I(N__82517));
    LocalMux I__18789 (
            .O(N__82523),
            .I(N__82517));
    InMux I__18788 (
            .O(N__82522),
            .I(N__82514));
    Span4Mux_h I__18787 (
            .O(N__82517),
            .I(N__82511));
    LocalMux I__18786 (
            .O(N__82514),
            .I(N__82508));
    Odrv4 I__18785 (
            .O(N__82511),
            .I(\quad_counter1.n3306 ));
    Odrv4 I__18784 (
            .O(N__82508),
            .I(\quad_counter1.n3306 ));
    InMux I__18783 (
            .O(N__82503),
            .I(\quad_counter1.n30667 ));
    InMux I__18782 (
            .O(N__82500),
            .I(N__82496));
    InMux I__18781 (
            .O(N__82499),
            .I(N__82493));
    LocalMux I__18780 (
            .O(N__82496),
            .I(N__82488));
    LocalMux I__18779 (
            .O(N__82493),
            .I(N__82488));
    Span4Mux_h I__18778 (
            .O(N__82488),
            .I(N__82484));
    InMux I__18777 (
            .O(N__82487),
            .I(N__82481));
    Odrv4 I__18776 (
            .O(N__82484),
            .I(\quad_counter1.n3305 ));
    LocalMux I__18775 (
            .O(N__82481),
            .I(\quad_counter1.n3305 ));
    InMux I__18774 (
            .O(N__82476),
            .I(\quad_counter1.n30668 ));
    InMux I__18773 (
            .O(N__82473),
            .I(N__82469));
    InMux I__18772 (
            .O(N__82472),
            .I(N__82466));
    LocalMux I__18771 (
            .O(N__82469),
            .I(N__82463));
    LocalMux I__18770 (
            .O(N__82466),
            .I(\quad_counter1.millisecond_counter_1 ));
    Odrv12 I__18769 (
            .O(N__82463),
            .I(\quad_counter1.millisecond_counter_1 ));
    InMux I__18768 (
            .O(N__82458),
            .I(N__82454));
    InMux I__18767 (
            .O(N__82457),
            .I(N__82451));
    LocalMux I__18766 (
            .O(N__82454),
            .I(N__82448));
    LocalMux I__18765 (
            .O(N__82451),
            .I(\quad_counter1.millisecond_counter_7 ));
    Odrv12 I__18764 (
            .O(N__82448),
            .I(\quad_counter1.millisecond_counter_7 ));
    CascadeMux I__18763 (
            .O(N__82443),
            .I(\quad_counter1.n34519_cascade_ ));
    InMux I__18762 (
            .O(N__82440),
            .I(N__82436));
    InMux I__18761 (
            .O(N__82439),
            .I(N__82433));
    LocalMux I__18760 (
            .O(N__82436),
            .I(N__82430));
    LocalMux I__18759 (
            .O(N__82433),
            .I(\quad_counter1.millisecond_counter_5 ));
    Odrv12 I__18758 (
            .O(N__82430),
            .I(\quad_counter1.millisecond_counter_5 ));
    InMux I__18757 (
            .O(N__82425),
            .I(N__82422));
    LocalMux I__18756 (
            .O(N__82422),
            .I(\quad_counter1.n12_adj_4467 ));
    InMux I__18755 (
            .O(N__82419),
            .I(N__82414));
    InMux I__18754 (
            .O(N__82418),
            .I(N__82411));
    InMux I__18753 (
            .O(N__82417),
            .I(N__82407));
    LocalMux I__18752 (
            .O(N__82414),
            .I(N__82402));
    LocalMux I__18751 (
            .O(N__82411),
            .I(N__82402));
    InMux I__18750 (
            .O(N__82410),
            .I(N__82399));
    LocalMux I__18749 (
            .O(N__82407),
            .I(N__82396));
    Span4Mux_v I__18748 (
            .O(N__82402),
            .I(N__82393));
    LocalMux I__18747 (
            .O(N__82399),
            .I(N__82388));
    Span4Mux_v I__18746 (
            .O(N__82396),
            .I(N__82388));
    Odrv4 I__18745 (
            .O(N__82393),
            .I(\quad_counter1.millisecond_counter_10 ));
    Odrv4 I__18744 (
            .O(N__82388),
            .I(\quad_counter1.millisecond_counter_10 ));
    InMux I__18743 (
            .O(N__82383),
            .I(bfn_22_13_0_));
    InMux I__18742 (
            .O(N__82380),
            .I(N__82376));
    InMux I__18741 (
            .O(N__82379),
            .I(N__82373));
    LocalMux I__18740 (
            .O(N__82376),
            .I(N__82368));
    LocalMux I__18739 (
            .O(N__82373),
            .I(N__82368));
    Span4Mux_v I__18738 (
            .O(N__82368),
            .I(N__82364));
    InMux I__18737 (
            .O(N__82367),
            .I(N__82361));
    Odrv4 I__18736 (
            .O(N__82364),
            .I(\quad_counter1.n3319 ));
    LocalMux I__18735 (
            .O(N__82361),
            .I(\quad_counter1.n3319 ));
    InMux I__18734 (
            .O(N__82356),
            .I(\quad_counter1.n30654 ));
    InMux I__18733 (
            .O(N__82353),
            .I(N__82349));
    InMux I__18732 (
            .O(N__82352),
            .I(N__82346));
    LocalMux I__18731 (
            .O(N__82349),
            .I(N__82340));
    LocalMux I__18730 (
            .O(N__82346),
            .I(N__82340));
    CascadeMux I__18729 (
            .O(N__82345),
            .I(N__82337));
    Span4Mux_v I__18728 (
            .O(N__82340),
            .I(N__82334));
    InMux I__18727 (
            .O(N__82337),
            .I(N__82331));
    Odrv4 I__18726 (
            .O(N__82334),
            .I(\quad_counter1.n3318 ));
    LocalMux I__18725 (
            .O(N__82331),
            .I(\quad_counter1.n3318 ));
    InMux I__18724 (
            .O(N__82326),
            .I(\quad_counter1.n30655 ));
    InMux I__18723 (
            .O(N__82323),
            .I(N__82319));
    InMux I__18722 (
            .O(N__82322),
            .I(N__82316));
    LocalMux I__18721 (
            .O(N__82319),
            .I(N__82311));
    LocalMux I__18720 (
            .O(N__82316),
            .I(N__82311));
    Span4Mux_v I__18719 (
            .O(N__82311),
            .I(N__82307));
    InMux I__18718 (
            .O(N__82310),
            .I(N__82304));
    Odrv4 I__18717 (
            .O(N__82307),
            .I(\quad_counter1.n3317 ));
    LocalMux I__18716 (
            .O(N__82304),
            .I(\quad_counter1.n3317 ));
    InMux I__18715 (
            .O(N__82299),
            .I(\quad_counter1.n30656 ));
    InMux I__18714 (
            .O(N__82296),
            .I(N__82292));
    InMux I__18713 (
            .O(N__82295),
            .I(N__82289));
    LocalMux I__18712 (
            .O(N__82292),
            .I(N__82284));
    LocalMux I__18711 (
            .O(N__82289),
            .I(N__82284));
    Span4Mux_v I__18710 (
            .O(N__82284),
            .I(N__82280));
    InMux I__18709 (
            .O(N__82283),
            .I(N__82277));
    Odrv4 I__18708 (
            .O(N__82280),
            .I(\quad_counter1.n3316 ));
    LocalMux I__18707 (
            .O(N__82277),
            .I(\quad_counter1.n3316 ));
    InMux I__18706 (
            .O(N__82272),
            .I(\quad_counter1.n30657 ));
    InMux I__18705 (
            .O(N__82269),
            .I(N__82265));
    InMux I__18704 (
            .O(N__82268),
            .I(N__82262));
    LocalMux I__18703 (
            .O(N__82265),
            .I(N__82257));
    LocalMux I__18702 (
            .O(N__82262),
            .I(N__82257));
    Span4Mux_h I__18701 (
            .O(N__82257),
            .I(N__82253));
    InMux I__18700 (
            .O(N__82256),
            .I(N__82250));
    Odrv4 I__18699 (
            .O(N__82253),
            .I(\quad_counter1.n3315 ));
    LocalMux I__18698 (
            .O(N__82250),
            .I(\quad_counter1.n3315 ));
    InMux I__18697 (
            .O(N__82245),
            .I(\quad_counter1.n30658 ));
    InMux I__18696 (
            .O(N__82242),
            .I(N__82238));
    InMux I__18695 (
            .O(N__82241),
            .I(N__82235));
    LocalMux I__18694 (
            .O(N__82238),
            .I(N__82229));
    LocalMux I__18693 (
            .O(N__82235),
            .I(N__82229));
    CascadeMux I__18692 (
            .O(N__82234),
            .I(N__82226));
    Span4Mux_v I__18691 (
            .O(N__82229),
            .I(N__82223));
    InMux I__18690 (
            .O(N__82226),
            .I(N__82220));
    Odrv4 I__18689 (
            .O(N__82223),
            .I(\quad_counter1.n3314 ));
    LocalMux I__18688 (
            .O(N__82220),
            .I(\quad_counter1.n3314 ));
    CascadeMux I__18687 (
            .O(N__82215),
            .I(N__82207));
    CascadeMux I__18686 (
            .O(N__82214),
            .I(N__82204));
    CascadeMux I__18685 (
            .O(N__82213),
            .I(N__82201));
    CascadeMux I__18684 (
            .O(N__82212),
            .I(N__82198));
    CascadeMux I__18683 (
            .O(N__82211),
            .I(N__82195));
    CascadeMux I__18682 (
            .O(N__82210),
            .I(N__82192));
    InMux I__18681 (
            .O(N__82207),
            .I(N__82187));
    InMux I__18680 (
            .O(N__82204),
            .I(N__82187));
    InMux I__18679 (
            .O(N__82201),
            .I(N__82178));
    InMux I__18678 (
            .O(N__82198),
            .I(N__82178));
    InMux I__18677 (
            .O(N__82195),
            .I(N__82178));
    InMux I__18676 (
            .O(N__82192),
            .I(N__82178));
    LocalMux I__18675 (
            .O(N__82187),
            .I(\quad_counter1.n36146 ));
    LocalMux I__18674 (
            .O(N__82178),
            .I(\quad_counter1.n36146 ));
    InMux I__18673 (
            .O(N__82173),
            .I(\quad_counter1.n30659 ));
    InMux I__18672 (
            .O(N__82170),
            .I(\quad_counter1.n30450 ));
    InMux I__18671 (
            .O(N__82167),
            .I(N__82164));
    LocalMux I__18670 (
            .O(N__82164),
            .I(\quad_counter1.n12935 ));
    InMux I__18669 (
            .O(N__82161),
            .I(N__82158));
    LocalMux I__18668 (
            .O(N__82158),
            .I(\quad_counter1.n8_adj_4453 ));
    InMux I__18667 (
            .O(N__82155),
            .I(\quad_counter1.n30451 ));
    InMux I__18666 (
            .O(N__82152),
            .I(N__82149));
    LocalMux I__18665 (
            .O(N__82149),
            .I(\quad_counter1.n12934 ));
    InMux I__18664 (
            .O(N__82146),
            .I(\quad_counter1.n30452 ));
    InMux I__18663 (
            .O(N__82143),
            .I(N__82140));
    LocalMux I__18662 (
            .O(N__82140),
            .I(\quad_counter1.n9_adj_4452 ));
    InMux I__18661 (
            .O(N__82137),
            .I(N__82134));
    LocalMux I__18660 (
            .O(N__82134),
            .I(\quad_counter1.n35987 ));
    InMux I__18659 (
            .O(N__82131),
            .I(N__82128));
    LocalMux I__18658 (
            .O(N__82128),
            .I(\quad_counter1.n10_adj_4454 ));
    CascadeMux I__18657 (
            .O(N__82125),
            .I(\quad_counter1.n31_adj_4461_cascade_ ));
    InMux I__18656 (
            .O(N__82122),
            .I(N__82119));
    LocalMux I__18655 (
            .O(N__82119),
            .I(\quad_counter1.n35986 ));
    CascadeMux I__18654 (
            .O(N__82116),
            .I(\quad_counter1.n34_adj_4465_cascade_ ));
    InMux I__18653 (
            .O(N__82113),
            .I(N__82109));
    InMux I__18652 (
            .O(N__82112),
            .I(N__82106));
    LocalMux I__18651 (
            .O(N__82109),
            .I(N__82103));
    LocalMux I__18650 (
            .O(N__82106),
            .I(\quad_counter1.millisecond_counter_3 ));
    Odrv12 I__18649 (
            .O(N__82103),
            .I(\quad_counter1.millisecond_counter_3 ));
    CascadeMux I__18648 (
            .O(N__82098),
            .I(\quad_counter1.n34207_cascade_ ));
    InMux I__18647 (
            .O(N__82095),
            .I(N__82092));
    LocalMux I__18646 (
            .O(N__82092),
            .I(N__82088));
    InMux I__18645 (
            .O(N__82091),
            .I(N__82085));
    Span4Mux_v I__18644 (
            .O(N__82088),
            .I(N__82082));
    LocalMux I__18643 (
            .O(N__82085),
            .I(\quad_counter1.millisecond_counter_0 ));
    Odrv4 I__18642 (
            .O(N__82082),
            .I(\quad_counter1.millisecond_counter_0 ));
    InMux I__18641 (
            .O(N__82077),
            .I(\quad_counter1.n30197 ));
    InMux I__18640 (
            .O(N__82074),
            .I(\quad_counter1.n30198 ));
    InMux I__18639 (
            .O(N__82071),
            .I(\quad_counter1.n30199 ));
    InMux I__18638 (
            .O(N__82068),
            .I(\quad_counter1.n30200 ));
    InMux I__18637 (
            .O(N__82065),
            .I(\quad_counter1.n30201 ));
    InMux I__18636 (
            .O(N__82062),
            .I(bfn_22_11_0_));
    InMux I__18635 (
            .O(N__82059),
            .I(\quad_counter1.n30447 ));
    InMux I__18634 (
            .O(N__82056),
            .I(\quad_counter1.n30448 ));
    InMux I__18633 (
            .O(N__82053),
            .I(N__82050));
    LocalMux I__18632 (
            .O(N__82050),
            .I(\quad_counter1.n12936 ));
    InMux I__18631 (
            .O(N__82047),
            .I(\quad_counter1.n30449 ));
    InMux I__18630 (
            .O(N__82044),
            .I(\quad_counter1.n30187 ));
    InMux I__18629 (
            .O(N__82041),
            .I(\quad_counter1.n30188 ));
    InMux I__18628 (
            .O(N__82038),
            .I(\quad_counter1.n30189 ));
    InMux I__18627 (
            .O(N__82035),
            .I(\quad_counter1.n30190 ));
    InMux I__18626 (
            .O(N__82032),
            .I(\quad_counter1.n30191 ));
    InMux I__18625 (
            .O(N__82029),
            .I(\quad_counter1.n30192 ));
    InMux I__18624 (
            .O(N__82026),
            .I(\quad_counter1.n30193 ));
    InMux I__18623 (
            .O(N__82023),
            .I(bfn_22_10_0_));
    InMux I__18622 (
            .O(N__82020),
            .I(\quad_counter1.n30195 ));
    InMux I__18621 (
            .O(N__82017),
            .I(\quad_counter1.n30196 ));
    InMux I__18620 (
            .O(N__82014),
            .I(\quad_counter1.n30179 ));
    InMux I__18619 (
            .O(N__82011),
            .I(\quad_counter1.n30180 ));
    InMux I__18618 (
            .O(N__82008),
            .I(N__82004));
    InMux I__18617 (
            .O(N__82007),
            .I(N__82001));
    LocalMux I__18616 (
            .O(N__82004),
            .I(N__81994));
    LocalMux I__18615 (
            .O(N__82001),
            .I(N__81994));
    InMux I__18614 (
            .O(N__82000),
            .I(N__81991));
    InMux I__18613 (
            .O(N__81999),
            .I(N__81988));
    Span4Mux_h I__18612 (
            .O(N__81994),
            .I(N__81985));
    LocalMux I__18611 (
            .O(N__81991),
            .I(N__81982));
    LocalMux I__18610 (
            .O(N__81988),
            .I(\quad_counter1.millisecond_counter_11 ));
    Odrv4 I__18609 (
            .O(N__81985),
            .I(\quad_counter1.millisecond_counter_11 ));
    Odrv4 I__18608 (
            .O(N__81982),
            .I(\quad_counter1.millisecond_counter_11 ));
    InMux I__18607 (
            .O(N__81975),
            .I(\quad_counter1.n30181 ));
    InMux I__18606 (
            .O(N__81972),
            .I(N__81967));
    InMux I__18605 (
            .O(N__81971),
            .I(N__81964));
    InMux I__18604 (
            .O(N__81970),
            .I(N__81961));
    LocalMux I__18603 (
            .O(N__81967),
            .I(N__81957));
    LocalMux I__18602 (
            .O(N__81964),
            .I(N__81954));
    LocalMux I__18601 (
            .O(N__81961),
            .I(N__81951));
    InMux I__18600 (
            .O(N__81960),
            .I(N__81948));
    Span4Mux_h I__18599 (
            .O(N__81957),
            .I(N__81943));
    Span4Mux_h I__18598 (
            .O(N__81954),
            .I(N__81943));
    Span4Mux_h I__18597 (
            .O(N__81951),
            .I(N__81940));
    LocalMux I__18596 (
            .O(N__81948),
            .I(\quad_counter1.millisecond_counter_12 ));
    Odrv4 I__18595 (
            .O(N__81943),
            .I(\quad_counter1.millisecond_counter_12 ));
    Odrv4 I__18594 (
            .O(N__81940),
            .I(\quad_counter1.millisecond_counter_12 ));
    InMux I__18593 (
            .O(N__81933),
            .I(\quad_counter1.n30182 ));
    InMux I__18592 (
            .O(N__81930),
            .I(N__81925));
    InMux I__18591 (
            .O(N__81929),
            .I(N__81922));
    InMux I__18590 (
            .O(N__81928),
            .I(N__81919));
    LocalMux I__18589 (
            .O(N__81925),
            .I(N__81916));
    LocalMux I__18588 (
            .O(N__81922),
            .I(N__81913));
    LocalMux I__18587 (
            .O(N__81919),
            .I(N__81910));
    Span4Mux_v I__18586 (
            .O(N__81916),
            .I(N__81906));
    Span4Mux_v I__18585 (
            .O(N__81913),
            .I(N__81903));
    Span4Mux_h I__18584 (
            .O(N__81910),
            .I(N__81900));
    InMux I__18583 (
            .O(N__81909),
            .I(N__81897));
    Span4Mux_v I__18582 (
            .O(N__81906),
            .I(N__81892));
    Span4Mux_h I__18581 (
            .O(N__81903),
            .I(N__81892));
    Span4Mux_h I__18580 (
            .O(N__81900),
            .I(N__81889));
    LocalMux I__18579 (
            .O(N__81897),
            .I(\quad_counter1.millisecond_counter_13 ));
    Odrv4 I__18578 (
            .O(N__81892),
            .I(\quad_counter1.millisecond_counter_13 ));
    Odrv4 I__18577 (
            .O(N__81889),
            .I(\quad_counter1.millisecond_counter_13 ));
    InMux I__18576 (
            .O(N__81882),
            .I(\quad_counter1.n30183 ));
    InMux I__18575 (
            .O(N__81879),
            .I(N__81874));
    InMux I__18574 (
            .O(N__81878),
            .I(N__81871));
    InMux I__18573 (
            .O(N__81877),
            .I(N__81868));
    LocalMux I__18572 (
            .O(N__81874),
            .I(N__81861));
    LocalMux I__18571 (
            .O(N__81871),
            .I(N__81861));
    LocalMux I__18570 (
            .O(N__81868),
            .I(N__81861));
    Span4Mux_v I__18569 (
            .O(N__81861),
            .I(N__81857));
    InMux I__18568 (
            .O(N__81860),
            .I(N__81854));
    Span4Mux_h I__18567 (
            .O(N__81857),
            .I(N__81851));
    LocalMux I__18566 (
            .O(N__81854),
            .I(\quad_counter1.millisecond_counter_14 ));
    Odrv4 I__18565 (
            .O(N__81851),
            .I(\quad_counter1.millisecond_counter_14 ));
    InMux I__18564 (
            .O(N__81846),
            .I(\quad_counter1.n30184 ));
    InMux I__18563 (
            .O(N__81843),
            .I(N__81838));
    InMux I__18562 (
            .O(N__81842),
            .I(N__81835));
    InMux I__18561 (
            .O(N__81841),
            .I(N__81832));
    LocalMux I__18560 (
            .O(N__81838),
            .I(N__81826));
    LocalMux I__18559 (
            .O(N__81835),
            .I(N__81826));
    LocalMux I__18558 (
            .O(N__81832),
            .I(N__81823));
    InMux I__18557 (
            .O(N__81831),
            .I(N__81820));
    Span12Mux_s7_v I__18556 (
            .O(N__81826),
            .I(N__81817));
    Span12Mux_h I__18555 (
            .O(N__81823),
            .I(N__81814));
    LocalMux I__18554 (
            .O(N__81820),
            .I(\quad_counter1.millisecond_counter_15 ));
    Odrv12 I__18553 (
            .O(N__81817),
            .I(\quad_counter1.millisecond_counter_15 ));
    Odrv12 I__18552 (
            .O(N__81814),
            .I(\quad_counter1.millisecond_counter_15 ));
    InMux I__18551 (
            .O(N__81807),
            .I(\quad_counter1.n30185 ));
    InMux I__18550 (
            .O(N__81804),
            .I(N__81800));
    InMux I__18549 (
            .O(N__81803),
            .I(N__81797));
    LocalMux I__18548 (
            .O(N__81800),
            .I(N__81791));
    LocalMux I__18547 (
            .O(N__81797),
            .I(N__81791));
    InMux I__18546 (
            .O(N__81796),
            .I(N__81788));
    Span4Mux_v I__18545 (
            .O(N__81791),
            .I(N__81784));
    LocalMux I__18544 (
            .O(N__81788),
            .I(N__81781));
    InMux I__18543 (
            .O(N__81787),
            .I(N__81778));
    Span4Mux_v I__18542 (
            .O(N__81784),
            .I(N__81775));
    Span4Mux_v I__18541 (
            .O(N__81781),
            .I(N__81772));
    LocalMux I__18540 (
            .O(N__81778),
            .I(\quad_counter1.millisecond_counter_16 ));
    Odrv4 I__18539 (
            .O(N__81775),
            .I(\quad_counter1.millisecond_counter_16 ));
    Odrv4 I__18538 (
            .O(N__81772),
            .I(\quad_counter1.millisecond_counter_16 ));
    InMux I__18537 (
            .O(N__81765),
            .I(bfn_22_9_0_));
    InMux I__18536 (
            .O(N__81762),
            .I(bfn_22_7_0_));
    InMux I__18535 (
            .O(N__81759),
            .I(\quad_counter1.n30171 ));
    InMux I__18534 (
            .O(N__81756),
            .I(N__81753));
    LocalMux I__18533 (
            .O(N__81753),
            .I(N__81750));
    Span4Mux_v I__18532 (
            .O(N__81750),
            .I(N__81746));
    InMux I__18531 (
            .O(N__81749),
            .I(N__81743));
    Odrv4 I__18530 (
            .O(N__81746),
            .I(\quad_counter1.millisecond_counter_2 ));
    LocalMux I__18529 (
            .O(N__81743),
            .I(\quad_counter1.millisecond_counter_2 ));
    InMux I__18528 (
            .O(N__81738),
            .I(\quad_counter1.n30172 ));
    InMux I__18527 (
            .O(N__81735),
            .I(\quad_counter1.n30173 ));
    CascadeMux I__18526 (
            .O(N__81732),
            .I(N__81729));
    InMux I__18525 (
            .O(N__81729),
            .I(N__81726));
    LocalMux I__18524 (
            .O(N__81726),
            .I(N__81723));
    Span4Mux_v I__18523 (
            .O(N__81723),
            .I(N__81719));
    InMux I__18522 (
            .O(N__81722),
            .I(N__81716));
    Odrv4 I__18521 (
            .O(N__81719),
            .I(\quad_counter1.millisecond_counter_4 ));
    LocalMux I__18520 (
            .O(N__81716),
            .I(\quad_counter1.millisecond_counter_4 ));
    InMux I__18519 (
            .O(N__81711),
            .I(\quad_counter1.n30174 ));
    InMux I__18518 (
            .O(N__81708),
            .I(\quad_counter1.n30175 ));
    InMux I__18517 (
            .O(N__81705),
            .I(N__81702));
    LocalMux I__18516 (
            .O(N__81702),
            .I(N__81699));
    Span4Mux_v I__18515 (
            .O(N__81699),
            .I(N__81695));
    InMux I__18514 (
            .O(N__81698),
            .I(N__81692));
    Odrv4 I__18513 (
            .O(N__81695),
            .I(\quad_counter1.millisecond_counter_6 ));
    LocalMux I__18512 (
            .O(N__81692),
            .I(\quad_counter1.millisecond_counter_6 ));
    InMux I__18511 (
            .O(N__81687),
            .I(\quad_counter1.n30176 ));
    InMux I__18510 (
            .O(N__81684),
            .I(\quad_counter1.n30177 ));
    InMux I__18509 (
            .O(N__81681),
            .I(bfn_22_8_0_));
    InMux I__18508 (
            .O(N__81678),
            .I(N__81673));
    InMux I__18507 (
            .O(N__81677),
            .I(N__81670));
    InMux I__18506 (
            .O(N__81676),
            .I(N__81667));
    LocalMux I__18505 (
            .O(N__81673),
            .I(\quad_counter1.n2706 ));
    LocalMux I__18504 (
            .O(N__81670),
            .I(\quad_counter1.n2706 ));
    LocalMux I__18503 (
            .O(N__81667),
            .I(\quad_counter1.n2706 ));
    InMux I__18502 (
            .O(N__81660),
            .I(N__81657));
    LocalMux I__18501 (
            .O(N__81657),
            .I(\quad_counter1.n14_adj_4470 ));
    CascadeMux I__18500 (
            .O(N__81654),
            .I(\quad_counter1.n18_adj_4471_cascade_ ));
    InMux I__18499 (
            .O(N__81651),
            .I(N__81646));
    InMux I__18498 (
            .O(N__81650),
            .I(N__81643));
    InMux I__18497 (
            .O(N__81649),
            .I(N__81640));
    LocalMux I__18496 (
            .O(N__81646),
            .I(\quad_counter1.n2710 ));
    LocalMux I__18495 (
            .O(N__81643),
            .I(\quad_counter1.n2710 ));
    LocalMux I__18494 (
            .O(N__81640),
            .I(\quad_counter1.n2710 ));
    CascadeMux I__18493 (
            .O(N__81633),
            .I(N__81621));
    CascadeMux I__18492 (
            .O(N__81632),
            .I(N__81618));
    CascadeMux I__18491 (
            .O(N__81631),
            .I(N__81615));
    CascadeMux I__18490 (
            .O(N__81630),
            .I(N__81612));
    CascadeMux I__18489 (
            .O(N__81629),
            .I(N__81609));
    CascadeMux I__18488 (
            .O(N__81628),
            .I(N__81606));
    CascadeMux I__18487 (
            .O(N__81627),
            .I(N__81603));
    CascadeMux I__18486 (
            .O(N__81626),
            .I(N__81600));
    CascadeMux I__18485 (
            .O(N__81625),
            .I(N__81597));
    CascadeMux I__18484 (
            .O(N__81624),
            .I(N__81594));
    InMux I__18483 (
            .O(N__81621),
            .I(N__81589));
    InMux I__18482 (
            .O(N__81618),
            .I(N__81589));
    InMux I__18481 (
            .O(N__81615),
            .I(N__81580));
    InMux I__18480 (
            .O(N__81612),
            .I(N__81580));
    InMux I__18479 (
            .O(N__81609),
            .I(N__81580));
    InMux I__18478 (
            .O(N__81606),
            .I(N__81580));
    InMux I__18477 (
            .O(N__81603),
            .I(N__81571));
    InMux I__18476 (
            .O(N__81600),
            .I(N__81571));
    InMux I__18475 (
            .O(N__81597),
            .I(N__81571));
    InMux I__18474 (
            .O(N__81594),
            .I(N__81571));
    LocalMux I__18473 (
            .O(N__81589),
            .I(N__81568));
    LocalMux I__18472 (
            .O(N__81580),
            .I(N__81562));
    LocalMux I__18471 (
            .O(N__81571),
            .I(N__81562));
    Span4Mux_h I__18470 (
            .O(N__81568),
            .I(N__81559));
    InMux I__18469 (
            .O(N__81567),
            .I(N__81556));
    Odrv4 I__18468 (
            .O(N__81562),
            .I(\quad_counter1.n2738 ));
    Odrv4 I__18467 (
            .O(N__81559),
            .I(\quad_counter1.n2738 ));
    LocalMux I__18466 (
            .O(N__81556),
            .I(\quad_counter1.n2738 ));
    InMux I__18465 (
            .O(N__81549),
            .I(N__81544));
    InMux I__18464 (
            .O(N__81548),
            .I(N__81541));
    InMux I__18463 (
            .O(N__81547),
            .I(N__81538));
    LocalMux I__18462 (
            .O(N__81544),
            .I(N__81533));
    LocalMux I__18461 (
            .O(N__81541),
            .I(N__81533));
    LocalMux I__18460 (
            .O(N__81538),
            .I(N__81530));
    Span4Mux_v I__18459 (
            .O(N__81533),
            .I(N__81525));
    Span4Mux_h I__18458 (
            .O(N__81530),
            .I(N__81525));
    Odrv4 I__18457 (
            .O(N__81525),
            .I(\quad_counter1.n3219 ));
    InMux I__18456 (
            .O(N__81522),
            .I(N__81517));
    InMux I__18455 (
            .O(N__81521),
            .I(N__81514));
    InMux I__18454 (
            .O(N__81520),
            .I(N__81511));
    LocalMux I__18453 (
            .O(N__81517),
            .I(N__81506));
    LocalMux I__18452 (
            .O(N__81514),
            .I(N__81506));
    LocalMux I__18451 (
            .O(N__81511),
            .I(N__81503));
    Span4Mux_v I__18450 (
            .O(N__81506),
            .I(N__81500));
    Span4Mux_h I__18449 (
            .O(N__81503),
            .I(N__81497));
    Odrv4 I__18448 (
            .O(N__81500),
            .I(\quad_counter1.n3218 ));
    Odrv4 I__18447 (
            .O(N__81497),
            .I(\quad_counter1.n3218 ));
    InMux I__18446 (
            .O(N__81492),
            .I(N__81487));
    InMux I__18445 (
            .O(N__81491),
            .I(N__81484));
    InMux I__18444 (
            .O(N__81490),
            .I(N__81481));
    LocalMux I__18443 (
            .O(N__81487),
            .I(N__81478));
    LocalMux I__18442 (
            .O(N__81484),
            .I(N__81475));
    LocalMux I__18441 (
            .O(N__81481),
            .I(N__81470));
    Span4Mux_h I__18440 (
            .O(N__81478),
            .I(N__81470));
    Span4Mux_v I__18439 (
            .O(N__81475),
            .I(N__81467));
    Odrv4 I__18438 (
            .O(N__81470),
            .I(\quad_counter1.n3214 ));
    Odrv4 I__18437 (
            .O(N__81467),
            .I(\quad_counter1.n3214 ));
    CascadeMux I__18436 (
            .O(N__81462),
            .I(\quad_counter1.n28243_cascade_ ));
    InMux I__18435 (
            .O(N__81459),
            .I(N__81455));
    InMux I__18434 (
            .O(N__81458),
            .I(N__81451));
    LocalMux I__18433 (
            .O(N__81455),
            .I(N__81448));
    InMux I__18432 (
            .O(N__81454),
            .I(N__81445));
    LocalMux I__18431 (
            .O(N__81451),
            .I(N__81442));
    Span4Mux_h I__18430 (
            .O(N__81448),
            .I(N__81437));
    LocalMux I__18429 (
            .O(N__81445),
            .I(N__81437));
    Span4Mux_h I__18428 (
            .O(N__81442),
            .I(N__81434));
    Odrv4 I__18427 (
            .O(N__81437),
            .I(\quad_counter1.n3217 ));
    Odrv4 I__18426 (
            .O(N__81434),
            .I(\quad_counter1.n3217 ));
    InMux I__18425 (
            .O(N__81429),
            .I(N__81426));
    LocalMux I__18424 (
            .O(N__81426),
            .I(N__81423));
    Span4Mux_h I__18423 (
            .O(N__81423),
            .I(N__81420));
    Odrv4 I__18422 (
            .O(N__81420),
            .I(\quad_counter1.n10_adj_4483 ));
    CascadeMux I__18421 (
            .O(N__81417),
            .I(\quad_counter1.n10_cascade_ ));
    CascadeMux I__18420 (
            .O(N__81414),
            .I(\quad_counter1.n16_cascade_ ));
    CascadeMux I__18419 (
            .O(N__81411),
            .I(N__81400));
    CascadeMux I__18418 (
            .O(N__81410),
            .I(N__81397));
    CascadeMux I__18417 (
            .O(N__81409),
            .I(N__81394));
    CascadeMux I__18416 (
            .O(N__81408),
            .I(N__81391));
    CascadeMux I__18415 (
            .O(N__81407),
            .I(N__81388));
    CascadeMux I__18414 (
            .O(N__81406),
            .I(N__81385));
    CascadeMux I__18413 (
            .O(N__81405),
            .I(N__81382));
    CascadeMux I__18412 (
            .O(N__81404),
            .I(N__81379));
    CascadeMux I__18411 (
            .O(N__81403),
            .I(N__81376));
    InMux I__18410 (
            .O(N__81400),
            .I(N__81369));
    InMux I__18409 (
            .O(N__81397),
            .I(N__81369));
    InMux I__18408 (
            .O(N__81394),
            .I(N__81369));
    InMux I__18407 (
            .O(N__81391),
            .I(N__81360));
    InMux I__18406 (
            .O(N__81388),
            .I(N__81360));
    InMux I__18405 (
            .O(N__81385),
            .I(N__81360));
    InMux I__18404 (
            .O(N__81382),
            .I(N__81360));
    InMux I__18403 (
            .O(N__81379),
            .I(N__81355));
    InMux I__18402 (
            .O(N__81376),
            .I(N__81355));
    LocalMux I__18401 (
            .O(N__81369),
            .I(\quad_counter1.n2639 ));
    LocalMux I__18400 (
            .O(N__81360),
            .I(\quad_counter1.n2639 ));
    LocalMux I__18399 (
            .O(N__81355),
            .I(\quad_counter1.n2639 ));
    CascadeMux I__18398 (
            .O(N__81348),
            .I(\quad_counter1.n2639_cascade_ ));
    CascadeMux I__18397 (
            .O(N__81345),
            .I(N__81337));
    CascadeMux I__18396 (
            .O(N__81344),
            .I(N__81334));
    CascadeMux I__18395 (
            .O(N__81343),
            .I(N__81331));
    CascadeMux I__18394 (
            .O(N__81342),
            .I(N__81328));
    CascadeMux I__18393 (
            .O(N__81341),
            .I(N__81325));
    CascadeMux I__18392 (
            .O(N__81340),
            .I(N__81322));
    InMux I__18391 (
            .O(N__81337),
            .I(N__81317));
    InMux I__18390 (
            .O(N__81334),
            .I(N__81317));
    InMux I__18389 (
            .O(N__81331),
            .I(N__81308));
    InMux I__18388 (
            .O(N__81328),
            .I(N__81308));
    InMux I__18387 (
            .O(N__81325),
            .I(N__81308));
    InMux I__18386 (
            .O(N__81322),
            .I(N__81308));
    LocalMux I__18385 (
            .O(N__81317),
            .I(\quad_counter1.n36132 ));
    LocalMux I__18384 (
            .O(N__81308),
            .I(\quad_counter1.n36132 ));
    InMux I__18383 (
            .O(N__81303),
            .I(N__81300));
    LocalMux I__18382 (
            .O(N__81300),
            .I(N__81297));
    Span4Mux_v I__18381 (
            .O(N__81297),
            .I(N__81294));
    Span4Mux_h I__18380 (
            .O(N__81294),
            .I(N__81290));
    InMux I__18379 (
            .O(N__81293),
            .I(N__81287));
    Span4Mux_v I__18378 (
            .O(N__81290),
            .I(N__81284));
    LocalMux I__18377 (
            .O(N__81287),
            .I(data_out_frame_11_3));
    Odrv4 I__18376 (
            .O(N__81284),
            .I(data_out_frame_11_3));
    InMux I__18375 (
            .O(N__81279),
            .I(N__81276));
    LocalMux I__18374 (
            .O(N__81276),
            .I(N__81272));
    InMux I__18373 (
            .O(N__81275),
            .I(N__81267));
    Span4Mux_v I__18372 (
            .O(N__81272),
            .I(N__81264));
    InMux I__18371 (
            .O(N__81271),
            .I(N__81261));
    InMux I__18370 (
            .O(N__81270),
            .I(N__81257));
    LocalMux I__18369 (
            .O(N__81267),
            .I(N__81254));
    Span4Mux_h I__18368 (
            .O(N__81264),
            .I(N__81249));
    LocalMux I__18367 (
            .O(N__81261),
            .I(N__81249));
    CascadeMux I__18366 (
            .O(N__81260),
            .I(N__81237));
    LocalMux I__18365 (
            .O(N__81257),
            .I(N__81234));
    Span4Mux_v I__18364 (
            .O(N__81254),
            .I(N__81229));
    Span4Mux_v I__18363 (
            .O(N__81249),
            .I(N__81229));
    InMux I__18362 (
            .O(N__81248),
            .I(N__81226));
    InMux I__18361 (
            .O(N__81247),
            .I(N__81217));
    InMux I__18360 (
            .O(N__81246),
            .I(N__81214));
    InMux I__18359 (
            .O(N__81245),
            .I(N__81210));
    InMux I__18358 (
            .O(N__81244),
            .I(N__81207));
    InMux I__18357 (
            .O(N__81243),
            .I(N__81204));
    InMux I__18356 (
            .O(N__81242),
            .I(N__81196));
    InMux I__18355 (
            .O(N__81241),
            .I(N__81196));
    InMux I__18354 (
            .O(N__81240),
            .I(N__81191));
    InMux I__18353 (
            .O(N__81237),
            .I(N__81191));
    Span4Mux_h I__18352 (
            .O(N__81234),
            .I(N__81184));
    Span4Mux_v I__18351 (
            .O(N__81229),
            .I(N__81184));
    LocalMux I__18350 (
            .O(N__81226),
            .I(N__81184));
    InMux I__18349 (
            .O(N__81225),
            .I(N__81181));
    InMux I__18348 (
            .O(N__81224),
            .I(N__81178));
    InMux I__18347 (
            .O(N__81223),
            .I(N__81175));
    InMux I__18346 (
            .O(N__81222),
            .I(N__81169));
    InMux I__18345 (
            .O(N__81221),
            .I(N__81166));
    InMux I__18344 (
            .O(N__81220),
            .I(N__81163));
    LocalMux I__18343 (
            .O(N__81217),
            .I(N__81160));
    LocalMux I__18342 (
            .O(N__81214),
            .I(N__81157));
    InMux I__18341 (
            .O(N__81213),
            .I(N__81154));
    LocalMux I__18340 (
            .O(N__81210),
            .I(N__81151));
    LocalMux I__18339 (
            .O(N__81207),
            .I(N__81148));
    LocalMux I__18338 (
            .O(N__81204),
            .I(N__81145));
    CascadeMux I__18337 (
            .O(N__81203),
            .I(N__81142));
    InMux I__18336 (
            .O(N__81202),
            .I(N__81139));
    InMux I__18335 (
            .O(N__81201),
            .I(N__81136));
    LocalMux I__18334 (
            .O(N__81196),
            .I(N__81133));
    LocalMux I__18333 (
            .O(N__81191),
            .I(N__81126));
    Span4Mux_h I__18332 (
            .O(N__81184),
            .I(N__81126));
    LocalMux I__18331 (
            .O(N__81181),
            .I(N__81126));
    LocalMux I__18330 (
            .O(N__81178),
            .I(N__81123));
    LocalMux I__18329 (
            .O(N__81175),
            .I(N__81120));
    CascadeMux I__18328 (
            .O(N__81174),
            .I(N__81117));
    InMux I__18327 (
            .O(N__81173),
            .I(N__81113));
    InMux I__18326 (
            .O(N__81172),
            .I(N__81110));
    LocalMux I__18325 (
            .O(N__81169),
            .I(N__81105));
    LocalMux I__18324 (
            .O(N__81166),
            .I(N__81105));
    LocalMux I__18323 (
            .O(N__81163),
            .I(N__81100));
    Span4Mux_v I__18322 (
            .O(N__81160),
            .I(N__81097));
    Span4Mux_v I__18321 (
            .O(N__81157),
            .I(N__81094));
    LocalMux I__18320 (
            .O(N__81154),
            .I(N__81089));
    Span4Mux_v I__18319 (
            .O(N__81151),
            .I(N__81089));
    Span4Mux_h I__18318 (
            .O(N__81148),
            .I(N__81084));
    Span4Mux_v I__18317 (
            .O(N__81145),
            .I(N__81084));
    InMux I__18316 (
            .O(N__81142),
            .I(N__81081));
    LocalMux I__18315 (
            .O(N__81139),
            .I(N__81076));
    LocalMux I__18314 (
            .O(N__81136),
            .I(N__81076));
    Span4Mux_v I__18313 (
            .O(N__81133),
            .I(N__81073));
    Span4Mux_h I__18312 (
            .O(N__81126),
            .I(N__81066));
    Span4Mux_h I__18311 (
            .O(N__81123),
            .I(N__81066));
    Span4Mux_v I__18310 (
            .O(N__81120),
            .I(N__81066));
    InMux I__18309 (
            .O(N__81117),
            .I(N__81063));
    InMux I__18308 (
            .O(N__81116),
            .I(N__81060));
    LocalMux I__18307 (
            .O(N__81113),
            .I(N__81055));
    LocalMux I__18306 (
            .O(N__81110),
            .I(N__81055));
    Span4Mux_h I__18305 (
            .O(N__81105),
            .I(N__81052));
    InMux I__18304 (
            .O(N__81104),
            .I(N__81047));
    InMux I__18303 (
            .O(N__81103),
            .I(N__81047));
    Span4Mux_v I__18302 (
            .O(N__81100),
            .I(N__81036));
    Span4Mux_h I__18301 (
            .O(N__81097),
            .I(N__81036));
    Span4Mux_v I__18300 (
            .O(N__81094),
            .I(N__81036));
    Span4Mux_v I__18299 (
            .O(N__81089),
            .I(N__81036));
    Span4Mux_v I__18298 (
            .O(N__81084),
            .I(N__81036));
    LocalMux I__18297 (
            .O(N__81081),
            .I(N__81027));
    Span4Mux_v I__18296 (
            .O(N__81076),
            .I(N__81027));
    Span4Mux_v I__18295 (
            .O(N__81073),
            .I(N__81027));
    Span4Mux_v I__18294 (
            .O(N__81066),
            .I(N__81027));
    LocalMux I__18293 (
            .O(N__81063),
            .I(N__81022));
    LocalMux I__18292 (
            .O(N__81060),
            .I(N__81015));
    Span4Mux_v I__18291 (
            .O(N__81055),
            .I(N__81015));
    Span4Mux_h I__18290 (
            .O(N__81052),
            .I(N__81015));
    LocalMux I__18289 (
            .O(N__81047),
            .I(N__81012));
    Sp12to4 I__18288 (
            .O(N__81036),
            .I(N__81007));
    Sp12to4 I__18287 (
            .O(N__81027),
            .I(N__81007));
    InMux I__18286 (
            .O(N__81026),
            .I(N__81004));
    InMux I__18285 (
            .O(N__81025),
            .I(N__81001));
    Span4Mux_h I__18284 (
            .O(N__81022),
            .I(N__80998));
    Span4Mux_h I__18283 (
            .O(N__81015),
            .I(N__80995));
    Span12Mux_s7_v I__18282 (
            .O(N__81012),
            .I(N__80990));
    Span12Mux_h I__18281 (
            .O(N__81007),
            .I(N__80990));
    LocalMux I__18280 (
            .O(N__81004),
            .I(\c0.n9 ));
    LocalMux I__18279 (
            .O(N__81001),
            .I(\c0.n9 ));
    Odrv4 I__18278 (
            .O(N__80998),
            .I(\c0.n9 ));
    Odrv4 I__18277 (
            .O(N__80995),
            .I(\c0.n9 ));
    Odrv12 I__18276 (
            .O(N__80990),
            .I(\c0.n9 ));
    CascadeMux I__18275 (
            .O(N__80979),
            .I(N__80971));
    InMux I__18274 (
            .O(N__80978),
            .I(N__80963));
    InMux I__18273 (
            .O(N__80977),
            .I(N__80963));
    InMux I__18272 (
            .O(N__80976),
            .I(N__80960));
    InMux I__18271 (
            .O(N__80975),
            .I(N__80957));
    InMux I__18270 (
            .O(N__80974),
            .I(N__80950));
    InMux I__18269 (
            .O(N__80971),
            .I(N__80943));
    InMux I__18268 (
            .O(N__80970),
            .I(N__80943));
    InMux I__18267 (
            .O(N__80969),
            .I(N__80943));
    InMux I__18266 (
            .O(N__80968),
            .I(N__80940));
    LocalMux I__18265 (
            .O(N__80963),
            .I(N__80937));
    LocalMux I__18264 (
            .O(N__80960),
            .I(N__80934));
    LocalMux I__18263 (
            .O(N__80957),
            .I(N__80927));
    InMux I__18262 (
            .O(N__80956),
            .I(N__80918));
    InMux I__18261 (
            .O(N__80955),
            .I(N__80915));
    InMux I__18260 (
            .O(N__80954),
            .I(N__80912));
    InMux I__18259 (
            .O(N__80953),
            .I(N__80907));
    LocalMux I__18258 (
            .O(N__80950),
            .I(N__80903));
    LocalMux I__18257 (
            .O(N__80943),
            .I(N__80900));
    LocalMux I__18256 (
            .O(N__80940),
            .I(N__80895));
    Span4Mux_v I__18255 (
            .O(N__80937),
            .I(N__80895));
    Span4Mux_v I__18254 (
            .O(N__80934),
            .I(N__80892));
    InMux I__18253 (
            .O(N__80933),
            .I(N__80889));
    InMux I__18252 (
            .O(N__80932),
            .I(N__80884));
    InMux I__18251 (
            .O(N__80931),
            .I(N__80884));
    InMux I__18250 (
            .O(N__80930),
            .I(N__80881));
    Span4Mux_v I__18249 (
            .O(N__80927),
            .I(N__80878));
    InMux I__18248 (
            .O(N__80926),
            .I(N__80873));
    InMux I__18247 (
            .O(N__80925),
            .I(N__80870));
    CascadeMux I__18246 (
            .O(N__80924),
            .I(N__80867));
    InMux I__18245 (
            .O(N__80923),
            .I(N__80862));
    InMux I__18244 (
            .O(N__80922),
            .I(N__80857));
    InMux I__18243 (
            .O(N__80921),
            .I(N__80857));
    LocalMux I__18242 (
            .O(N__80918),
            .I(N__80850));
    LocalMux I__18241 (
            .O(N__80915),
            .I(N__80850));
    LocalMux I__18240 (
            .O(N__80912),
            .I(N__80850));
    InMux I__18239 (
            .O(N__80911),
            .I(N__80845));
    InMux I__18238 (
            .O(N__80910),
            .I(N__80845));
    LocalMux I__18237 (
            .O(N__80907),
            .I(N__80842));
    InMux I__18236 (
            .O(N__80906),
            .I(N__80839));
    Span4Mux_h I__18235 (
            .O(N__80903),
            .I(N__80836));
    Span4Mux_h I__18234 (
            .O(N__80900),
            .I(N__80825));
    Span4Mux_h I__18233 (
            .O(N__80895),
            .I(N__80825));
    Span4Mux_h I__18232 (
            .O(N__80892),
            .I(N__80825));
    LocalMux I__18231 (
            .O(N__80889),
            .I(N__80825));
    LocalMux I__18230 (
            .O(N__80884),
            .I(N__80825));
    LocalMux I__18229 (
            .O(N__80881),
            .I(N__80822));
    Span4Mux_v I__18228 (
            .O(N__80878),
            .I(N__80819));
    InMux I__18227 (
            .O(N__80877),
            .I(N__80814));
    InMux I__18226 (
            .O(N__80876),
            .I(N__80814));
    LocalMux I__18225 (
            .O(N__80873),
            .I(N__80809));
    LocalMux I__18224 (
            .O(N__80870),
            .I(N__80809));
    InMux I__18223 (
            .O(N__80867),
            .I(N__80804));
    InMux I__18222 (
            .O(N__80866),
            .I(N__80799));
    InMux I__18221 (
            .O(N__80865),
            .I(N__80799));
    LocalMux I__18220 (
            .O(N__80862),
            .I(N__80796));
    LocalMux I__18219 (
            .O(N__80857),
            .I(N__80793));
    Span4Mux_v I__18218 (
            .O(N__80850),
            .I(N__80790));
    LocalMux I__18217 (
            .O(N__80845),
            .I(N__80785));
    Span4Mux_h I__18216 (
            .O(N__80842),
            .I(N__80785));
    LocalMux I__18215 (
            .O(N__80839),
            .I(N__80782));
    Span4Mux_h I__18214 (
            .O(N__80836),
            .I(N__80777));
    Span4Mux_v I__18213 (
            .O(N__80825),
            .I(N__80777));
    Span4Mux_v I__18212 (
            .O(N__80822),
            .I(N__80772));
    Span4Mux_h I__18211 (
            .O(N__80819),
            .I(N__80772));
    LocalMux I__18210 (
            .O(N__80814),
            .I(N__80767));
    Sp12to4 I__18209 (
            .O(N__80809),
            .I(N__80767));
    InMux I__18208 (
            .O(N__80808),
            .I(N__80764));
    InMux I__18207 (
            .O(N__80807),
            .I(N__80761));
    LocalMux I__18206 (
            .O(N__80804),
            .I(N__80758));
    LocalMux I__18205 (
            .O(N__80799),
            .I(N__80749));
    Span4Mux_h I__18204 (
            .O(N__80796),
            .I(N__80749));
    Span4Mux_v I__18203 (
            .O(N__80793),
            .I(N__80749));
    Span4Mux_h I__18202 (
            .O(N__80790),
            .I(N__80749));
    Span4Mux_h I__18201 (
            .O(N__80785),
            .I(N__80746));
    Span4Mux_v I__18200 (
            .O(N__80782),
            .I(N__80741));
    Span4Mux_v I__18199 (
            .O(N__80777),
            .I(N__80741));
    Sp12to4 I__18198 (
            .O(N__80772),
            .I(N__80736));
    Span12Mux_v I__18197 (
            .O(N__80767),
            .I(N__80736));
    LocalMux I__18196 (
            .O(N__80764),
            .I(rx_data_0));
    LocalMux I__18195 (
            .O(N__80761),
            .I(rx_data_0));
    Odrv12 I__18194 (
            .O(N__80758),
            .I(rx_data_0));
    Odrv4 I__18193 (
            .O(N__80749),
            .I(rx_data_0));
    Odrv4 I__18192 (
            .O(N__80746),
            .I(rx_data_0));
    Odrv4 I__18191 (
            .O(N__80741),
            .I(rx_data_0));
    Odrv12 I__18190 (
            .O(N__80736),
            .I(rx_data_0));
    InMux I__18189 (
            .O(N__80721),
            .I(N__80713));
    InMux I__18188 (
            .O(N__80720),
            .I(N__80713));
    InMux I__18187 (
            .O(N__80719),
            .I(N__80705));
    InMux I__18186 (
            .O(N__80718),
            .I(N__80702));
    LocalMux I__18185 (
            .O(N__80713),
            .I(N__80697));
    InMux I__18184 (
            .O(N__80712),
            .I(N__80694));
    InMux I__18183 (
            .O(N__80711),
            .I(N__80690));
    InMux I__18182 (
            .O(N__80710),
            .I(N__80685));
    InMux I__18181 (
            .O(N__80709),
            .I(N__80681));
    InMux I__18180 (
            .O(N__80708),
            .I(N__80677));
    LocalMux I__18179 (
            .O(N__80705),
            .I(N__80671));
    LocalMux I__18178 (
            .O(N__80702),
            .I(N__80671));
    InMux I__18177 (
            .O(N__80701),
            .I(N__80668));
    InMux I__18176 (
            .O(N__80700),
            .I(N__80665));
    Span4Mux_h I__18175 (
            .O(N__80697),
            .I(N__80658));
    LocalMux I__18174 (
            .O(N__80694),
            .I(N__80658));
    InMux I__18173 (
            .O(N__80693),
            .I(N__80655));
    LocalMux I__18172 (
            .O(N__80690),
            .I(N__80652));
    InMux I__18171 (
            .O(N__80689),
            .I(N__80647));
    InMux I__18170 (
            .O(N__80688),
            .I(N__80647));
    LocalMux I__18169 (
            .O(N__80685),
            .I(N__80644));
    InMux I__18168 (
            .O(N__80684),
            .I(N__80641));
    LocalMux I__18167 (
            .O(N__80681),
            .I(N__80637));
    InMux I__18166 (
            .O(N__80680),
            .I(N__80634));
    LocalMux I__18165 (
            .O(N__80677),
            .I(N__80630));
    InMux I__18164 (
            .O(N__80676),
            .I(N__80627));
    Span4Mux_v I__18163 (
            .O(N__80671),
            .I(N__80624));
    LocalMux I__18162 (
            .O(N__80668),
            .I(N__80619));
    LocalMux I__18161 (
            .O(N__80665),
            .I(N__80619));
    InMux I__18160 (
            .O(N__80664),
            .I(N__80612));
    InMux I__18159 (
            .O(N__80663),
            .I(N__80612));
    Span4Mux_v I__18158 (
            .O(N__80658),
            .I(N__80607));
    LocalMux I__18157 (
            .O(N__80655),
            .I(N__80607));
    Span4Mux_v I__18156 (
            .O(N__80652),
            .I(N__80602));
    LocalMux I__18155 (
            .O(N__80647),
            .I(N__80602));
    Span4Mux_v I__18154 (
            .O(N__80644),
            .I(N__80596));
    LocalMux I__18153 (
            .O(N__80641),
            .I(N__80596));
    CascadeMux I__18152 (
            .O(N__80640),
            .I(N__80593));
    Span4Mux_v I__18151 (
            .O(N__80637),
            .I(N__80587));
    LocalMux I__18150 (
            .O(N__80634),
            .I(N__80587));
    InMux I__18149 (
            .O(N__80633),
            .I(N__80584));
    Span4Mux_v I__18148 (
            .O(N__80630),
            .I(N__80575));
    LocalMux I__18147 (
            .O(N__80627),
            .I(N__80575));
    Span4Mux_h I__18146 (
            .O(N__80624),
            .I(N__80575));
    Span4Mux_v I__18145 (
            .O(N__80619),
            .I(N__80575));
    CascadeMux I__18144 (
            .O(N__80618),
            .I(N__80572));
    InMux I__18143 (
            .O(N__80617),
            .I(N__80569));
    LocalMux I__18142 (
            .O(N__80612),
            .I(N__80564));
    Span4Mux_v I__18141 (
            .O(N__80607),
            .I(N__80564));
    Span4Mux_v I__18140 (
            .O(N__80602),
            .I(N__80561));
    InMux I__18139 (
            .O(N__80601),
            .I(N__80558));
    Span4Mux_v I__18138 (
            .O(N__80596),
            .I(N__80555));
    InMux I__18137 (
            .O(N__80593),
            .I(N__80548));
    InMux I__18136 (
            .O(N__80592),
            .I(N__80548));
    Span4Mux_h I__18135 (
            .O(N__80587),
            .I(N__80544));
    LocalMux I__18134 (
            .O(N__80584),
            .I(N__80541));
    Span4Mux_h I__18133 (
            .O(N__80575),
            .I(N__80538));
    InMux I__18132 (
            .O(N__80572),
            .I(N__80534));
    LocalMux I__18131 (
            .O(N__80569),
            .I(N__80531));
    Span4Mux_v I__18130 (
            .O(N__80564),
            .I(N__80526));
    Span4Mux_h I__18129 (
            .O(N__80561),
            .I(N__80526));
    LocalMux I__18128 (
            .O(N__80558),
            .I(N__80523));
    Sp12to4 I__18127 (
            .O(N__80555),
            .I(N__80520));
    InMux I__18126 (
            .O(N__80554),
            .I(N__80514));
    InMux I__18125 (
            .O(N__80553),
            .I(N__80514));
    LocalMux I__18124 (
            .O(N__80548),
            .I(N__80511));
    InMux I__18123 (
            .O(N__80547),
            .I(N__80508));
    Span4Mux_h I__18122 (
            .O(N__80544),
            .I(N__80505));
    Span4Mux_v I__18121 (
            .O(N__80541),
            .I(N__80500));
    Span4Mux_h I__18120 (
            .O(N__80538),
            .I(N__80500));
    InMux I__18119 (
            .O(N__80537),
            .I(N__80495));
    LocalMux I__18118 (
            .O(N__80534),
            .I(N__80492));
    Span4Mux_h I__18117 (
            .O(N__80531),
            .I(N__80487));
    Span4Mux_h I__18116 (
            .O(N__80526),
            .I(N__80487));
    Span12Mux_h I__18115 (
            .O(N__80523),
            .I(N__80482));
    Span12Mux_h I__18114 (
            .O(N__80520),
            .I(N__80482));
    InMux I__18113 (
            .O(N__80519),
            .I(N__80479));
    LocalMux I__18112 (
            .O(N__80514),
            .I(N__80476));
    Span4Mux_v I__18111 (
            .O(N__80511),
            .I(N__80473));
    LocalMux I__18110 (
            .O(N__80508),
            .I(N__80466));
    Span4Mux_v I__18109 (
            .O(N__80505),
            .I(N__80466));
    Span4Mux_h I__18108 (
            .O(N__80500),
            .I(N__80466));
    InMux I__18107 (
            .O(N__80499),
            .I(N__80463));
    InMux I__18106 (
            .O(N__80498),
            .I(N__80460));
    LocalMux I__18105 (
            .O(N__80495),
            .I(N__80457));
    Span4Mux_v I__18104 (
            .O(N__80492),
            .I(N__80452));
    Span4Mux_v I__18103 (
            .O(N__80487),
            .I(N__80452));
    Span12Mux_v I__18102 (
            .O(N__80482),
            .I(N__80449));
    LocalMux I__18101 (
            .O(N__80479),
            .I(N__80440));
    Span4Mux_v I__18100 (
            .O(N__80476),
            .I(N__80440));
    Span4Mux_h I__18099 (
            .O(N__80473),
            .I(N__80440));
    Span4Mux_v I__18098 (
            .O(N__80466),
            .I(N__80440));
    LocalMux I__18097 (
            .O(N__80463),
            .I(rx_data_2));
    LocalMux I__18096 (
            .O(N__80460),
            .I(rx_data_2));
    Odrv4 I__18095 (
            .O(N__80457),
            .I(rx_data_2));
    Odrv4 I__18094 (
            .O(N__80452),
            .I(rx_data_2));
    Odrv12 I__18093 (
            .O(N__80449),
            .I(rx_data_2));
    Odrv4 I__18092 (
            .O(N__80440),
            .I(rx_data_2));
    CascadeMux I__18091 (
            .O(N__80427),
            .I(N__80424));
    InMux I__18090 (
            .O(N__80424),
            .I(N__80419));
    InMux I__18089 (
            .O(N__80423),
            .I(N__80416));
    InMux I__18088 (
            .O(N__80422),
            .I(N__80413));
    LocalMux I__18087 (
            .O(N__80419),
            .I(N__80403));
    LocalMux I__18086 (
            .O(N__80416),
            .I(N__80398));
    LocalMux I__18085 (
            .O(N__80413),
            .I(N__80398));
    CascadeMux I__18084 (
            .O(N__80412),
            .I(N__80392));
    InMux I__18083 (
            .O(N__80411),
            .I(N__80387));
    InMux I__18082 (
            .O(N__80410),
            .I(N__80387));
    CascadeMux I__18081 (
            .O(N__80409),
            .I(N__80382));
    InMux I__18080 (
            .O(N__80408),
            .I(N__80375));
    InMux I__18079 (
            .O(N__80407),
            .I(N__80375));
    InMux I__18078 (
            .O(N__80406),
            .I(N__80375));
    Span4Mux_v I__18077 (
            .O(N__80403),
            .I(N__80370));
    Span4Mux_v I__18076 (
            .O(N__80398),
            .I(N__80370));
    InMux I__18075 (
            .O(N__80397),
            .I(N__80367));
    CascadeMux I__18074 (
            .O(N__80396),
            .I(N__80363));
    CascadeMux I__18073 (
            .O(N__80395),
            .I(N__80358));
    InMux I__18072 (
            .O(N__80392),
            .I(N__80355));
    LocalMux I__18071 (
            .O(N__80387),
            .I(N__80352));
    InMux I__18070 (
            .O(N__80386),
            .I(N__80349));
    InMux I__18069 (
            .O(N__80385),
            .I(N__80344));
    InMux I__18068 (
            .O(N__80382),
            .I(N__80344));
    LocalMux I__18067 (
            .O(N__80375),
            .I(N__80337));
    Span4Mux_h I__18066 (
            .O(N__80370),
            .I(N__80337));
    LocalMux I__18065 (
            .O(N__80367),
            .I(N__80337));
    CascadeMux I__18064 (
            .O(N__80366),
            .I(N__80333));
    InMux I__18063 (
            .O(N__80363),
            .I(N__80328));
    InMux I__18062 (
            .O(N__80362),
            .I(N__80325));
    CascadeMux I__18061 (
            .O(N__80361),
            .I(N__80322));
    InMux I__18060 (
            .O(N__80358),
            .I(N__80316));
    LocalMux I__18059 (
            .O(N__80355),
            .I(N__80313));
    Span4Mux_v I__18058 (
            .O(N__80352),
            .I(N__80308));
    LocalMux I__18057 (
            .O(N__80349),
            .I(N__80308));
    LocalMux I__18056 (
            .O(N__80344),
            .I(N__80303));
    Span4Mux_v I__18055 (
            .O(N__80337),
            .I(N__80303));
    InMux I__18054 (
            .O(N__80336),
            .I(N__80300));
    InMux I__18053 (
            .O(N__80333),
            .I(N__80295));
    InMux I__18052 (
            .O(N__80332),
            .I(N__80292));
    InMux I__18051 (
            .O(N__80331),
            .I(N__80289));
    LocalMux I__18050 (
            .O(N__80328),
            .I(N__80286));
    LocalMux I__18049 (
            .O(N__80325),
            .I(N__80283));
    InMux I__18048 (
            .O(N__80322),
            .I(N__80280));
    InMux I__18047 (
            .O(N__80321),
            .I(N__80277));
    InMux I__18046 (
            .O(N__80320),
            .I(N__80274));
    CascadeMux I__18045 (
            .O(N__80319),
            .I(N__80270));
    LocalMux I__18044 (
            .O(N__80316),
            .I(N__80258));
    Span4Mux_v I__18043 (
            .O(N__80313),
            .I(N__80258));
    Span4Mux_h I__18042 (
            .O(N__80308),
            .I(N__80258));
    Span4Mux_v I__18041 (
            .O(N__80303),
            .I(N__80253));
    LocalMux I__18040 (
            .O(N__80300),
            .I(N__80253));
    InMux I__18039 (
            .O(N__80299),
            .I(N__80250));
    InMux I__18038 (
            .O(N__80298),
            .I(N__80247));
    LocalMux I__18037 (
            .O(N__80295),
            .I(N__80242));
    LocalMux I__18036 (
            .O(N__80292),
            .I(N__80242));
    LocalMux I__18035 (
            .O(N__80289),
            .I(N__80235));
    Span4Mux_v I__18034 (
            .O(N__80286),
            .I(N__80235));
    Span4Mux_h I__18033 (
            .O(N__80283),
            .I(N__80235));
    LocalMux I__18032 (
            .O(N__80280),
            .I(N__80232));
    LocalMux I__18031 (
            .O(N__80277),
            .I(N__80227));
    LocalMux I__18030 (
            .O(N__80274),
            .I(N__80227));
    InMux I__18029 (
            .O(N__80273),
            .I(N__80222));
    InMux I__18028 (
            .O(N__80270),
            .I(N__80222));
    InMux I__18027 (
            .O(N__80269),
            .I(N__80217));
    InMux I__18026 (
            .O(N__80268),
            .I(N__80217));
    InMux I__18025 (
            .O(N__80267),
            .I(N__80212));
    InMux I__18024 (
            .O(N__80266),
            .I(N__80212));
    InMux I__18023 (
            .O(N__80265),
            .I(N__80209));
    Span4Mux_h I__18022 (
            .O(N__80258),
            .I(N__80206));
    Span4Mux_v I__18021 (
            .O(N__80253),
            .I(N__80203));
    LocalMux I__18020 (
            .O(N__80250),
            .I(N__80200));
    LocalMux I__18019 (
            .O(N__80247),
            .I(N__80197));
    Span4Mux_v I__18018 (
            .O(N__80242),
            .I(N__80192));
    Span4Mux_h I__18017 (
            .O(N__80235),
            .I(N__80192));
    Span4Mux_v I__18016 (
            .O(N__80232),
            .I(N__80187));
    Span4Mux_v I__18015 (
            .O(N__80227),
            .I(N__80187));
    LocalMux I__18014 (
            .O(N__80222),
            .I(N__80182));
    LocalMux I__18013 (
            .O(N__80217),
            .I(N__80182));
    LocalMux I__18012 (
            .O(N__80212),
            .I(N__80175));
    LocalMux I__18011 (
            .O(N__80209),
            .I(N__80175));
    Span4Mux_h I__18010 (
            .O(N__80206),
            .I(N__80175));
    Sp12to4 I__18009 (
            .O(N__80203),
            .I(N__80172));
    Span4Mux_v I__18008 (
            .O(N__80200),
            .I(N__80165));
    Span4Mux_v I__18007 (
            .O(N__80197),
            .I(N__80165));
    Span4Mux_h I__18006 (
            .O(N__80192),
            .I(N__80165));
    Span4Mux_v I__18005 (
            .O(N__80187),
            .I(N__80162));
    Span12Mux_h I__18004 (
            .O(N__80182),
            .I(N__80155));
    Sp12to4 I__18003 (
            .O(N__80175),
            .I(N__80155));
    Span12Mux_h I__18002 (
            .O(N__80172),
            .I(N__80155));
    Span4Mux_h I__18001 (
            .O(N__80165),
            .I(N__80152));
    Odrv4 I__18000 (
            .O(N__80162),
            .I(\c0.n9_adj_4530 ));
    Odrv12 I__17999 (
            .O(N__80155),
            .I(\c0.n9_adj_4530 ));
    Odrv4 I__17998 (
            .O(N__80152),
            .I(\c0.n9_adj_4530 ));
    InMux I__17997 (
            .O(N__80145),
            .I(N__80141));
    InMux I__17996 (
            .O(N__80144),
            .I(N__80138));
    LocalMux I__17995 (
            .O(N__80141),
            .I(N__80132));
    LocalMux I__17994 (
            .O(N__80138),
            .I(N__80129));
    CascadeMux I__17993 (
            .O(N__80137),
            .I(N__80124));
    InMux I__17992 (
            .O(N__80136),
            .I(N__80116));
    InMux I__17991 (
            .O(N__80135),
            .I(N__80113));
    Span4Mux_h I__17990 (
            .O(N__80132),
            .I(N__80106));
    Span4Mux_v I__17989 (
            .O(N__80129),
            .I(N__80106));
    InMux I__17988 (
            .O(N__80128),
            .I(N__80103));
    InMux I__17987 (
            .O(N__80127),
            .I(N__80093));
    InMux I__17986 (
            .O(N__80124),
            .I(N__80093));
    InMux I__17985 (
            .O(N__80123),
            .I(N__80088));
    InMux I__17984 (
            .O(N__80122),
            .I(N__80088));
    InMux I__17983 (
            .O(N__80121),
            .I(N__80083));
    InMux I__17982 (
            .O(N__80120),
            .I(N__80083));
    InMux I__17981 (
            .O(N__80119),
            .I(N__80079));
    LocalMux I__17980 (
            .O(N__80116),
            .I(N__80074));
    LocalMux I__17979 (
            .O(N__80113),
            .I(N__80074));
    InMux I__17978 (
            .O(N__80112),
            .I(N__80071));
    InMux I__17977 (
            .O(N__80111),
            .I(N__80068));
    Span4Mux_h I__17976 (
            .O(N__80106),
            .I(N__80063));
    LocalMux I__17975 (
            .O(N__80103),
            .I(N__80063));
    InMux I__17974 (
            .O(N__80102),
            .I(N__80058));
    InMux I__17973 (
            .O(N__80101),
            .I(N__80058));
    InMux I__17972 (
            .O(N__80100),
            .I(N__80054));
    InMux I__17971 (
            .O(N__80099),
            .I(N__80048));
    InMux I__17970 (
            .O(N__80098),
            .I(N__80045));
    LocalMux I__17969 (
            .O(N__80093),
            .I(N__80042));
    LocalMux I__17968 (
            .O(N__80088),
            .I(N__80039));
    LocalMux I__17967 (
            .O(N__80083),
            .I(N__80036));
    CascadeMux I__17966 (
            .O(N__80082),
            .I(N__80033));
    LocalMux I__17965 (
            .O(N__80079),
            .I(N__80028));
    Span4Mux_v I__17964 (
            .O(N__80074),
            .I(N__80028));
    LocalMux I__17963 (
            .O(N__80071),
            .I(N__80023));
    LocalMux I__17962 (
            .O(N__80068),
            .I(N__80023));
    Span4Mux_v I__17961 (
            .O(N__80063),
            .I(N__80018));
    LocalMux I__17960 (
            .O(N__80058),
            .I(N__80018));
    InMux I__17959 (
            .O(N__80057),
            .I(N__80013));
    LocalMux I__17958 (
            .O(N__80054),
            .I(N__80010));
    InMux I__17957 (
            .O(N__80053),
            .I(N__80005));
    InMux I__17956 (
            .O(N__80052),
            .I(N__80002));
    InMux I__17955 (
            .O(N__80051),
            .I(N__79999));
    LocalMux I__17954 (
            .O(N__80048),
            .I(N__79994));
    LocalMux I__17953 (
            .O(N__80045),
            .I(N__79989));
    Span4Mux_v I__17952 (
            .O(N__80042),
            .I(N__79989));
    Span4Mux_v I__17951 (
            .O(N__80039),
            .I(N__79984));
    Span4Mux_v I__17950 (
            .O(N__80036),
            .I(N__79984));
    InMux I__17949 (
            .O(N__80033),
            .I(N__79981));
    Span4Mux_v I__17948 (
            .O(N__80028),
            .I(N__79978));
    Span4Mux_v I__17947 (
            .O(N__80023),
            .I(N__79973));
    Span4Mux_v I__17946 (
            .O(N__80018),
            .I(N__79973));
    InMux I__17945 (
            .O(N__80017),
            .I(N__79970));
    InMux I__17944 (
            .O(N__80016),
            .I(N__79967));
    LocalMux I__17943 (
            .O(N__80013),
            .I(N__79962));
    Span4Mux_h I__17942 (
            .O(N__80010),
            .I(N__79962));
    InMux I__17941 (
            .O(N__80009),
            .I(N__79957));
    InMux I__17940 (
            .O(N__80008),
            .I(N__79954));
    LocalMux I__17939 (
            .O(N__80005),
            .I(N__79951));
    LocalMux I__17938 (
            .O(N__80002),
            .I(N__79948));
    LocalMux I__17937 (
            .O(N__79999),
            .I(N__79945));
    InMux I__17936 (
            .O(N__79998),
            .I(N__79942));
    InMux I__17935 (
            .O(N__79997),
            .I(N__79939));
    Span4Mux_v I__17934 (
            .O(N__79994),
            .I(N__79932));
    Span4Mux_v I__17933 (
            .O(N__79989),
            .I(N__79932));
    Span4Mux_v I__17932 (
            .O(N__79984),
            .I(N__79932));
    LocalMux I__17931 (
            .O(N__79981),
            .I(N__79925));
    Span4Mux_h I__17930 (
            .O(N__79978),
            .I(N__79925));
    Span4Mux_v I__17929 (
            .O(N__79973),
            .I(N__79925));
    LocalMux I__17928 (
            .O(N__79970),
            .I(N__79918));
    LocalMux I__17927 (
            .O(N__79967),
            .I(N__79918));
    Sp12to4 I__17926 (
            .O(N__79962),
            .I(N__79918));
    InMux I__17925 (
            .O(N__79961),
            .I(N__79913));
    InMux I__17924 (
            .O(N__79960),
            .I(N__79913));
    LocalMux I__17923 (
            .O(N__79957),
            .I(N__79906));
    LocalMux I__17922 (
            .O(N__79954),
            .I(N__79906));
    Span4Mux_h I__17921 (
            .O(N__79951),
            .I(N__79906));
    Span4Mux_h I__17920 (
            .O(N__79948),
            .I(N__79901));
    Span4Mux_h I__17919 (
            .O(N__79945),
            .I(N__79901));
    LocalMux I__17918 (
            .O(N__79942),
            .I(N__79890));
    LocalMux I__17917 (
            .O(N__79939),
            .I(N__79890));
    Sp12to4 I__17916 (
            .O(N__79932),
            .I(N__79890));
    Sp12to4 I__17915 (
            .O(N__79925),
            .I(N__79890));
    Span12Mux_s11_v I__17914 (
            .O(N__79918),
            .I(N__79890));
    LocalMux I__17913 (
            .O(N__79913),
            .I(rx_data_7));
    Odrv4 I__17912 (
            .O(N__79906),
            .I(rx_data_7));
    Odrv4 I__17911 (
            .O(N__79901),
            .I(rx_data_7));
    Odrv12 I__17910 (
            .O(N__79890),
            .I(rx_data_7));
    CascadeMux I__17909 (
            .O(N__79881),
            .I(N__79875));
    InMux I__17908 (
            .O(N__79880),
            .I(N__79872));
    CascadeMux I__17907 (
            .O(N__79879),
            .I(N__79856));
    CascadeMux I__17906 (
            .O(N__79878),
            .I(N__79851));
    InMux I__17905 (
            .O(N__79875),
            .I(N__79839));
    LocalMux I__17904 (
            .O(N__79872),
            .I(N__79835));
    InMux I__17903 (
            .O(N__79871),
            .I(N__79830));
    InMux I__17902 (
            .O(N__79870),
            .I(N__79823));
    InMux I__17901 (
            .O(N__79869),
            .I(N__79823));
    InMux I__17900 (
            .O(N__79868),
            .I(N__79823));
    InMux I__17899 (
            .O(N__79867),
            .I(N__79809));
    InMux I__17898 (
            .O(N__79866),
            .I(N__79809));
    InMux I__17897 (
            .O(N__79865),
            .I(N__79809));
    InMux I__17896 (
            .O(N__79864),
            .I(N__79794));
    InMux I__17895 (
            .O(N__79863),
            .I(N__79794));
    InMux I__17894 (
            .O(N__79862),
            .I(N__79794));
    InMux I__17893 (
            .O(N__79861),
            .I(N__79794));
    InMux I__17892 (
            .O(N__79860),
            .I(N__79794));
    InMux I__17891 (
            .O(N__79859),
            .I(N__79794));
    InMux I__17890 (
            .O(N__79856),
            .I(N__79791));
    InMux I__17889 (
            .O(N__79855),
            .I(N__79786));
    InMux I__17888 (
            .O(N__79854),
            .I(N__79786));
    InMux I__17887 (
            .O(N__79851),
            .I(N__79783));
    InMux I__17886 (
            .O(N__79850),
            .I(N__79776));
    InMux I__17885 (
            .O(N__79849),
            .I(N__79776));
    InMux I__17884 (
            .O(N__79848),
            .I(N__79776));
    InMux I__17883 (
            .O(N__79847),
            .I(N__79773));
    InMux I__17882 (
            .O(N__79846),
            .I(N__79770));
    InMux I__17881 (
            .O(N__79845),
            .I(N__79767));
    InMux I__17880 (
            .O(N__79844),
            .I(N__79764));
    InMux I__17879 (
            .O(N__79843),
            .I(N__79759));
    InMux I__17878 (
            .O(N__79842),
            .I(N__79759));
    LocalMux I__17877 (
            .O(N__79839),
            .I(N__79756));
    InMux I__17876 (
            .O(N__79838),
            .I(N__79753));
    Span4Mux_h I__17875 (
            .O(N__79835),
            .I(N__79750));
    InMux I__17874 (
            .O(N__79834),
            .I(N__79747));
    InMux I__17873 (
            .O(N__79833),
            .I(N__79744));
    LocalMux I__17872 (
            .O(N__79830),
            .I(N__79739));
    LocalMux I__17871 (
            .O(N__79823),
            .I(N__79739));
    InMux I__17870 (
            .O(N__79822),
            .I(N__79734));
    InMux I__17869 (
            .O(N__79821),
            .I(N__79734));
    InMux I__17868 (
            .O(N__79820),
            .I(N__79727));
    InMux I__17867 (
            .O(N__79819),
            .I(N__79727));
    InMux I__17866 (
            .O(N__79818),
            .I(N__79727));
    InMux I__17865 (
            .O(N__79817),
            .I(N__79722));
    InMux I__17864 (
            .O(N__79816),
            .I(N__79722));
    LocalMux I__17863 (
            .O(N__79809),
            .I(N__79719));
    InMux I__17862 (
            .O(N__79808),
            .I(N__79714));
    InMux I__17861 (
            .O(N__79807),
            .I(N__79714));
    LocalMux I__17860 (
            .O(N__79794),
            .I(N__79711));
    LocalMux I__17859 (
            .O(N__79791),
            .I(N__79702));
    LocalMux I__17858 (
            .O(N__79786),
            .I(N__79702));
    LocalMux I__17857 (
            .O(N__79783),
            .I(N__79702));
    LocalMux I__17856 (
            .O(N__79776),
            .I(N__79702));
    LocalMux I__17855 (
            .O(N__79773),
            .I(N__79697));
    LocalMux I__17854 (
            .O(N__79770),
            .I(N__79697));
    LocalMux I__17853 (
            .O(N__79767),
            .I(N__79692));
    LocalMux I__17852 (
            .O(N__79764),
            .I(N__79692));
    LocalMux I__17851 (
            .O(N__79759),
            .I(N__79687));
    Span4Mux_h I__17850 (
            .O(N__79756),
            .I(N__79687));
    LocalMux I__17849 (
            .O(N__79753),
            .I(N__79684));
    Span4Mux_h I__17848 (
            .O(N__79750),
            .I(N__79667));
    LocalMux I__17847 (
            .O(N__79747),
            .I(N__79667));
    LocalMux I__17846 (
            .O(N__79744),
            .I(N__79667));
    Span4Mux_h I__17845 (
            .O(N__79739),
            .I(N__79667));
    LocalMux I__17844 (
            .O(N__79734),
            .I(N__79667));
    LocalMux I__17843 (
            .O(N__79727),
            .I(N__79667));
    LocalMux I__17842 (
            .O(N__79722),
            .I(N__79667));
    Span4Mux_v I__17841 (
            .O(N__79719),
            .I(N__79667));
    LocalMux I__17840 (
            .O(N__79714),
            .I(N__79664));
    Span4Mux_h I__17839 (
            .O(N__79711),
            .I(N__79659));
    Span4Mux_v I__17838 (
            .O(N__79702),
            .I(N__79659));
    Sp12to4 I__17837 (
            .O(N__79697),
            .I(N__79654));
    Span12Mux_h I__17836 (
            .O(N__79692),
            .I(N__79654));
    Span4Mux_v I__17835 (
            .O(N__79687),
            .I(N__79649));
    Span4Mux_h I__17834 (
            .O(N__79684),
            .I(N__79649));
    Span4Mux_v I__17833 (
            .O(N__79667),
            .I(N__79646));
    Span4Mux_v I__17832 (
            .O(N__79664),
            .I(N__79641));
    Span4Mux_h I__17831 (
            .O(N__79659),
            .I(N__79641));
    Odrv12 I__17830 (
            .O(N__79654),
            .I(\c0.n33257 ));
    Odrv4 I__17829 (
            .O(N__79649),
            .I(\c0.n33257 ));
    Odrv4 I__17828 (
            .O(N__79646),
            .I(\c0.n33257 ));
    Odrv4 I__17827 (
            .O(N__79641),
            .I(\c0.n33257 ));
    CascadeMux I__17826 (
            .O(N__79632),
            .I(N__79629));
    InMux I__17825 (
            .O(N__79629),
            .I(N__79624));
    CascadeMux I__17824 (
            .O(N__79628),
            .I(N__79620));
    InMux I__17823 (
            .O(N__79627),
            .I(N__79617));
    LocalMux I__17822 (
            .O(N__79624),
            .I(N__79614));
    InMux I__17821 (
            .O(N__79623),
            .I(N__79611));
    InMux I__17820 (
            .O(N__79620),
            .I(N__79608));
    LocalMux I__17819 (
            .O(N__79617),
            .I(N__79605));
    Span4Mux_h I__17818 (
            .O(N__79614),
            .I(N__79600));
    LocalMux I__17817 (
            .O(N__79611),
            .I(N__79600));
    LocalMux I__17816 (
            .O(N__79608),
            .I(\c0.data_in_frame_26_7 ));
    Odrv4 I__17815 (
            .O(N__79605),
            .I(\c0.data_in_frame_26_7 ));
    Odrv4 I__17814 (
            .O(N__79600),
            .I(\c0.data_in_frame_26_7 ));
    CascadeMux I__17813 (
            .O(N__79593),
            .I(N__79590));
    InMux I__17812 (
            .O(N__79590),
            .I(N__79586));
    InMux I__17811 (
            .O(N__79589),
            .I(N__79583));
    LocalMux I__17810 (
            .O(N__79586),
            .I(\c0.data_in_frame_26_2 ));
    LocalMux I__17809 (
            .O(N__79583),
            .I(\c0.data_in_frame_26_2 ));
    InMux I__17808 (
            .O(N__79578),
            .I(N__79573));
    CascadeMux I__17807 (
            .O(N__79577),
            .I(N__79570));
    InMux I__17806 (
            .O(N__79576),
            .I(N__79567));
    LocalMux I__17805 (
            .O(N__79573),
            .I(N__79564));
    InMux I__17804 (
            .O(N__79570),
            .I(N__79560));
    LocalMux I__17803 (
            .O(N__79567),
            .I(N__79555));
    Span12Mux_s6_v I__17802 (
            .O(N__79564),
            .I(N__79555));
    InMux I__17801 (
            .O(N__79563),
            .I(N__79552));
    LocalMux I__17800 (
            .O(N__79560),
            .I(\c0.data_in_frame_24_0 ));
    Odrv12 I__17799 (
            .O(N__79555),
            .I(\c0.data_in_frame_24_0 ));
    LocalMux I__17798 (
            .O(N__79552),
            .I(\c0.data_in_frame_24_0 ));
    InMux I__17797 (
            .O(N__79545),
            .I(N__79541));
    InMux I__17796 (
            .O(N__79544),
            .I(N__79538));
    LocalMux I__17795 (
            .O(N__79541),
            .I(N__79535));
    LocalMux I__17794 (
            .O(N__79538),
            .I(N__79532));
    Span4Mux_v I__17793 (
            .O(N__79535),
            .I(N__79529));
    Span4Mux_h I__17792 (
            .O(N__79532),
            .I(N__79526));
    Span4Mux_h I__17791 (
            .O(N__79529),
            .I(N__79522));
    Span4Mux_h I__17790 (
            .O(N__79526),
            .I(N__79519));
    InMux I__17789 (
            .O(N__79525),
            .I(N__79516));
    Odrv4 I__17788 (
            .O(N__79522),
            .I(\c0.n17627 ));
    Odrv4 I__17787 (
            .O(N__79519),
            .I(\c0.n17627 ));
    LocalMux I__17786 (
            .O(N__79516),
            .I(\c0.n17627 ));
    InMux I__17785 (
            .O(N__79509),
            .I(N__79505));
    InMux I__17784 (
            .O(N__79508),
            .I(N__79502));
    LocalMux I__17783 (
            .O(N__79505),
            .I(N__79497));
    LocalMux I__17782 (
            .O(N__79502),
            .I(N__79497));
    Span4Mux_h I__17781 (
            .O(N__79497),
            .I(N__79494));
    Span4Mux_h I__17780 (
            .O(N__79494),
            .I(N__79491));
    Odrv4 I__17779 (
            .O(N__79491),
            .I(\c0.n31545 ));
    CascadeMux I__17778 (
            .O(N__79488),
            .I(\c0.n31545_cascade_ ));
    InMux I__17777 (
            .O(N__79485),
            .I(N__79481));
    InMux I__17776 (
            .O(N__79484),
            .I(N__79478));
    LocalMux I__17775 (
            .O(N__79481),
            .I(N__79470));
    LocalMux I__17774 (
            .O(N__79478),
            .I(N__79470));
    InMux I__17773 (
            .O(N__79477),
            .I(N__79464));
    InMux I__17772 (
            .O(N__79476),
            .I(N__79464));
    InMux I__17771 (
            .O(N__79475),
            .I(N__79460));
    Span4Mux_v I__17770 (
            .O(N__79470),
            .I(N__79457));
    InMux I__17769 (
            .O(N__79469),
            .I(N__79454));
    LocalMux I__17768 (
            .O(N__79464),
            .I(N__79449));
    InMux I__17767 (
            .O(N__79463),
            .I(N__79446));
    LocalMux I__17766 (
            .O(N__79460),
            .I(N__79439));
    Sp12to4 I__17765 (
            .O(N__79457),
            .I(N__79439));
    LocalMux I__17764 (
            .O(N__79454),
            .I(N__79439));
    InMux I__17763 (
            .O(N__79453),
            .I(N__79434));
    InMux I__17762 (
            .O(N__79452),
            .I(N__79434));
    Span4Mux_h I__17761 (
            .O(N__79449),
            .I(N__79431));
    LocalMux I__17760 (
            .O(N__79446),
            .I(\c0.n18578 ));
    Odrv12 I__17759 (
            .O(N__79439),
            .I(\c0.n18578 ));
    LocalMux I__17758 (
            .O(N__79434),
            .I(\c0.n18578 ));
    Odrv4 I__17757 (
            .O(N__79431),
            .I(\c0.n18578 ));
    InMux I__17756 (
            .O(N__79422),
            .I(N__79415));
    InMux I__17755 (
            .O(N__79421),
            .I(N__79415));
    InMux I__17754 (
            .O(N__79420),
            .I(N__79412));
    LocalMux I__17753 (
            .O(N__79415),
            .I(\c0.data_in_frame_24_6 ));
    LocalMux I__17752 (
            .O(N__79412),
            .I(\c0.data_in_frame_24_6 ));
    InMux I__17751 (
            .O(N__79407),
            .I(N__79404));
    LocalMux I__17750 (
            .O(N__79404),
            .I(N__79401));
    Odrv12 I__17749 (
            .O(N__79401),
            .I(\c0.n20_adj_4698 ));
    CascadeMux I__17748 (
            .O(N__79398),
            .I(\c0.n19_adj_4699_cascade_ ));
    InMux I__17747 (
            .O(N__79395),
            .I(N__79391));
    InMux I__17746 (
            .O(N__79394),
            .I(N__79388));
    LocalMux I__17745 (
            .O(N__79391),
            .I(N__79383));
    LocalMux I__17744 (
            .O(N__79388),
            .I(N__79383));
    Span4Mux_h I__17743 (
            .O(N__79383),
            .I(N__79380));
    Odrv4 I__17742 (
            .O(N__79380),
            .I(\c0.n33819 ));
    InMux I__17741 (
            .O(N__79377),
            .I(N__79374));
    LocalMux I__17740 (
            .O(N__79374),
            .I(N__79371));
    Span4Mux_h I__17739 (
            .O(N__79371),
            .I(N__79368));
    Span4Mux_h I__17738 (
            .O(N__79368),
            .I(N__79365));
    Odrv4 I__17737 (
            .O(N__79365),
            .I(\c0.n32_adj_4705 ));
    InMux I__17736 (
            .O(N__79362),
            .I(N__79357));
    InMux I__17735 (
            .O(N__79361),
            .I(N__79354));
    InMux I__17734 (
            .O(N__79360),
            .I(N__79351));
    LocalMux I__17733 (
            .O(N__79357),
            .I(\quad_counter1.n2713 ));
    LocalMux I__17732 (
            .O(N__79354),
            .I(\quad_counter1.n2713 ));
    LocalMux I__17731 (
            .O(N__79351),
            .I(\quad_counter1.n2713 ));
    InMux I__17730 (
            .O(N__79344),
            .I(N__79339));
    InMux I__17729 (
            .O(N__79343),
            .I(N__79336));
    InMux I__17728 (
            .O(N__79342),
            .I(N__79333));
    LocalMux I__17727 (
            .O(N__79339),
            .I(\quad_counter1.n2705 ));
    LocalMux I__17726 (
            .O(N__79336),
            .I(\quad_counter1.n2705 ));
    LocalMux I__17725 (
            .O(N__79333),
            .I(\quad_counter1.n2705 ));
    CascadeMux I__17724 (
            .O(N__79326),
            .I(N__79321));
    InMux I__17723 (
            .O(N__79325),
            .I(N__79318));
    InMux I__17722 (
            .O(N__79324),
            .I(N__79315));
    InMux I__17721 (
            .O(N__79321),
            .I(N__79312));
    LocalMux I__17720 (
            .O(N__79318),
            .I(\quad_counter1.n2707 ));
    LocalMux I__17719 (
            .O(N__79315),
            .I(\quad_counter1.n2707 ));
    LocalMux I__17718 (
            .O(N__79312),
            .I(\quad_counter1.n2707 ));
    InMux I__17717 (
            .O(N__79305),
            .I(N__79300));
    InMux I__17716 (
            .O(N__79304),
            .I(N__79297));
    InMux I__17715 (
            .O(N__79303),
            .I(N__79294));
    LocalMux I__17714 (
            .O(N__79300),
            .I(\quad_counter1.n2709 ));
    LocalMux I__17713 (
            .O(N__79297),
            .I(\quad_counter1.n2709 ));
    LocalMux I__17712 (
            .O(N__79294),
            .I(\quad_counter1.n2709 ));
    InMux I__17711 (
            .O(N__79287),
            .I(N__79282));
    InMux I__17710 (
            .O(N__79286),
            .I(N__79279));
    InMux I__17709 (
            .O(N__79285),
            .I(N__79276));
    LocalMux I__17708 (
            .O(N__79282),
            .I(\quad_counter1.n2708 ));
    LocalMux I__17707 (
            .O(N__79279),
            .I(\quad_counter1.n2708 ));
    LocalMux I__17706 (
            .O(N__79276),
            .I(\quad_counter1.n2708 ));
    CascadeMux I__17705 (
            .O(N__79269),
            .I(\quad_counter1.n16_adj_4469_cascade_ ));
    InMux I__17704 (
            .O(N__79266),
            .I(N__79261));
    InMux I__17703 (
            .O(N__79265),
            .I(N__79258));
    InMux I__17702 (
            .O(N__79264),
            .I(N__79255));
    LocalMux I__17701 (
            .O(N__79261),
            .I(\quad_counter1.n2711 ));
    LocalMux I__17700 (
            .O(N__79258),
            .I(\quad_counter1.n2711 ));
    LocalMux I__17699 (
            .O(N__79255),
            .I(\quad_counter1.n2711 ));
    CascadeMux I__17698 (
            .O(N__79248),
            .I(N__79245));
    InMux I__17697 (
            .O(N__79245),
            .I(N__79240));
    InMux I__17696 (
            .O(N__79244),
            .I(N__79237));
    InMux I__17695 (
            .O(N__79243),
            .I(N__79234));
    LocalMux I__17694 (
            .O(N__79240),
            .I(N__79230));
    LocalMux I__17693 (
            .O(N__79237),
            .I(N__79227));
    LocalMux I__17692 (
            .O(N__79234),
            .I(N__79223));
    InMux I__17691 (
            .O(N__79233),
            .I(N__79218));
    Span4Mux_v I__17690 (
            .O(N__79230),
            .I(N__79213));
    Span4Mux_h I__17689 (
            .O(N__79227),
            .I(N__79213));
    InMux I__17688 (
            .O(N__79226),
            .I(N__79210));
    Span4Mux_h I__17687 (
            .O(N__79223),
            .I(N__79207));
    InMux I__17686 (
            .O(N__79222),
            .I(N__79202));
    InMux I__17685 (
            .O(N__79221),
            .I(N__79202));
    LocalMux I__17684 (
            .O(N__79218),
            .I(encoder0_position_12));
    Odrv4 I__17683 (
            .O(N__79213),
            .I(encoder0_position_12));
    LocalMux I__17682 (
            .O(N__79210),
            .I(encoder0_position_12));
    Odrv4 I__17681 (
            .O(N__79207),
            .I(encoder0_position_12));
    LocalMux I__17680 (
            .O(N__79202),
            .I(encoder0_position_12));
    InMux I__17679 (
            .O(N__79191),
            .I(N__79187));
    InMux I__17678 (
            .O(N__79190),
            .I(N__79184));
    LocalMux I__17677 (
            .O(N__79187),
            .I(N__79181));
    LocalMux I__17676 (
            .O(N__79184),
            .I(N__79176));
    Span4Mux_h I__17675 (
            .O(N__79181),
            .I(N__79173));
    InMux I__17674 (
            .O(N__79180),
            .I(N__79170));
    InMux I__17673 (
            .O(N__79179),
            .I(N__79167));
    Span4Mux_h I__17672 (
            .O(N__79176),
            .I(N__79162));
    Span4Mux_v I__17671 (
            .O(N__79173),
            .I(N__79162));
    LocalMux I__17670 (
            .O(N__79170),
            .I(encoder1_position_16));
    LocalMux I__17669 (
            .O(N__79167),
            .I(encoder1_position_16));
    Odrv4 I__17668 (
            .O(N__79162),
            .I(encoder1_position_16));
    CascadeMux I__17667 (
            .O(N__79155),
            .I(N__79149));
    InMux I__17666 (
            .O(N__79154),
            .I(N__79141));
    InMux I__17665 (
            .O(N__79153),
            .I(N__79141));
    InMux I__17664 (
            .O(N__79152),
            .I(N__79138));
    InMux I__17663 (
            .O(N__79149),
            .I(N__79133));
    InMux I__17662 (
            .O(N__79148),
            .I(N__79133));
    InMux I__17661 (
            .O(N__79147),
            .I(N__79130));
    CascadeMux I__17660 (
            .O(N__79146),
            .I(N__79127));
    LocalMux I__17659 (
            .O(N__79141),
            .I(N__79124));
    LocalMux I__17658 (
            .O(N__79138),
            .I(N__79121));
    LocalMux I__17657 (
            .O(N__79133),
            .I(N__79118));
    LocalMux I__17656 (
            .O(N__79130),
            .I(N__79114));
    InMux I__17655 (
            .O(N__79127),
            .I(N__79111));
    Span4Mux_v I__17654 (
            .O(N__79124),
            .I(N__79108));
    Span4Mux_h I__17653 (
            .O(N__79121),
            .I(N__79103));
    Span4Mux_h I__17652 (
            .O(N__79118),
            .I(N__79103));
    InMux I__17651 (
            .O(N__79117),
            .I(N__79100));
    Span12Mux_v I__17650 (
            .O(N__79114),
            .I(N__79097));
    LocalMux I__17649 (
            .O(N__79111),
            .I(N__79092));
    Span4Mux_h I__17648 (
            .O(N__79108),
            .I(N__79092));
    Span4Mux_h I__17647 (
            .O(N__79103),
            .I(N__79089));
    LocalMux I__17646 (
            .O(N__79100),
            .I(encoder0_position_27));
    Odrv12 I__17645 (
            .O(N__79097),
            .I(encoder0_position_27));
    Odrv4 I__17644 (
            .O(N__79092),
            .I(encoder0_position_27));
    Odrv4 I__17643 (
            .O(N__79089),
            .I(encoder0_position_27));
    InMux I__17642 (
            .O(N__79080),
            .I(N__79077));
    LocalMux I__17641 (
            .O(N__79077),
            .I(\c0.n33807 ));
    CascadeMux I__17640 (
            .O(N__79074),
            .I(\c0.n6_adj_4566_cascade_ ));
    InMux I__17639 (
            .O(N__79071),
            .I(N__79066));
    CascadeMux I__17638 (
            .O(N__79070),
            .I(N__79061));
    CascadeMux I__17637 (
            .O(N__79069),
            .I(N__79057));
    LocalMux I__17636 (
            .O(N__79066),
            .I(N__79054));
    InMux I__17635 (
            .O(N__79065),
            .I(N__79051));
    InMux I__17634 (
            .O(N__79064),
            .I(N__79048));
    InMux I__17633 (
            .O(N__79061),
            .I(N__79045));
    InMux I__17632 (
            .O(N__79060),
            .I(N__79042));
    InMux I__17631 (
            .O(N__79057),
            .I(N__79039));
    Span4Mux_h I__17630 (
            .O(N__79054),
            .I(N__79036));
    LocalMux I__17629 (
            .O(N__79051),
            .I(N__79031));
    LocalMux I__17628 (
            .O(N__79048),
            .I(N__79031));
    LocalMux I__17627 (
            .O(N__79045),
            .I(N__79027));
    LocalMux I__17626 (
            .O(N__79042),
            .I(N__79018));
    LocalMux I__17625 (
            .O(N__79039),
            .I(N__79018));
    Span4Mux_v I__17624 (
            .O(N__79036),
            .I(N__79018));
    Span4Mux_h I__17623 (
            .O(N__79031),
            .I(N__79018));
    InMux I__17622 (
            .O(N__79030),
            .I(N__79015));
    Span4Mux_v I__17621 (
            .O(N__79027),
            .I(N__79012));
    Span4Mux_h I__17620 (
            .O(N__79018),
            .I(N__79009));
    LocalMux I__17619 (
            .O(N__79015),
            .I(encoder0_position_29));
    Odrv4 I__17618 (
            .O(N__79012),
            .I(encoder0_position_29));
    Odrv4 I__17617 (
            .O(N__79009),
            .I(encoder0_position_29));
    InMux I__17616 (
            .O(N__79002),
            .I(N__78999));
    LocalMux I__17615 (
            .O(N__78999),
            .I(\c0.n18572 ));
    CascadeMux I__17614 (
            .O(N__78996),
            .I(N__78992));
    InMux I__17613 (
            .O(N__78995),
            .I(N__78983));
    InMux I__17612 (
            .O(N__78992),
            .I(N__78971));
    InMux I__17611 (
            .O(N__78991),
            .I(N__78971));
    InMux I__17610 (
            .O(N__78990),
            .I(N__78971));
    InMux I__17609 (
            .O(N__78989),
            .I(N__78966));
    InMux I__17608 (
            .O(N__78988),
            .I(N__78966));
    InMux I__17607 (
            .O(N__78987),
            .I(N__78958));
    InMux I__17606 (
            .O(N__78986),
            .I(N__78955));
    LocalMux I__17605 (
            .O(N__78983),
            .I(N__78952));
    InMux I__17604 (
            .O(N__78982),
            .I(N__78949));
    InMux I__17603 (
            .O(N__78981),
            .I(N__78943));
    InMux I__17602 (
            .O(N__78980),
            .I(N__78940));
    InMux I__17601 (
            .O(N__78979),
            .I(N__78937));
    InMux I__17600 (
            .O(N__78978),
            .I(N__78934));
    LocalMux I__17599 (
            .O(N__78971),
            .I(N__78931));
    LocalMux I__17598 (
            .O(N__78966),
            .I(N__78928));
    InMux I__17597 (
            .O(N__78965),
            .I(N__78925));
    InMux I__17596 (
            .O(N__78964),
            .I(N__78922));
    InMux I__17595 (
            .O(N__78963),
            .I(N__78917));
    InMux I__17594 (
            .O(N__78962),
            .I(N__78917));
    CascadeMux I__17593 (
            .O(N__78961),
            .I(N__78910));
    LocalMux I__17592 (
            .O(N__78958),
            .I(N__78900));
    LocalMux I__17591 (
            .O(N__78955),
            .I(N__78900));
    Span4Mux_h I__17590 (
            .O(N__78952),
            .I(N__78900));
    LocalMux I__17589 (
            .O(N__78949),
            .I(N__78897));
    InMux I__17588 (
            .O(N__78948),
            .I(N__78894));
    InMux I__17587 (
            .O(N__78947),
            .I(N__78889));
    InMux I__17586 (
            .O(N__78946),
            .I(N__78889));
    LocalMux I__17585 (
            .O(N__78943),
            .I(N__78886));
    LocalMux I__17584 (
            .O(N__78940),
            .I(N__78881));
    LocalMux I__17583 (
            .O(N__78937),
            .I(N__78881));
    LocalMux I__17582 (
            .O(N__78934),
            .I(N__78874));
    Span4Mux_h I__17581 (
            .O(N__78931),
            .I(N__78874));
    Span4Mux_v I__17580 (
            .O(N__78928),
            .I(N__78874));
    LocalMux I__17579 (
            .O(N__78925),
            .I(N__78871));
    LocalMux I__17578 (
            .O(N__78922),
            .I(N__78866));
    LocalMux I__17577 (
            .O(N__78917),
            .I(N__78866));
    InMux I__17576 (
            .O(N__78916),
            .I(N__78861));
    InMux I__17575 (
            .O(N__78915),
            .I(N__78861));
    InMux I__17574 (
            .O(N__78914),
            .I(N__78858));
    InMux I__17573 (
            .O(N__78913),
            .I(N__78853));
    InMux I__17572 (
            .O(N__78910),
            .I(N__78853));
    InMux I__17571 (
            .O(N__78909),
            .I(N__78848));
    InMux I__17570 (
            .O(N__78908),
            .I(N__78845));
    InMux I__17569 (
            .O(N__78907),
            .I(N__78842));
    Span4Mux_h I__17568 (
            .O(N__78900),
            .I(N__78839));
    Span4Mux_h I__17567 (
            .O(N__78897),
            .I(N__78834));
    LocalMux I__17566 (
            .O(N__78894),
            .I(N__78834));
    LocalMux I__17565 (
            .O(N__78889),
            .I(N__78831));
    Span4Mux_v I__17564 (
            .O(N__78886),
            .I(N__78828));
    Span4Mux_v I__17563 (
            .O(N__78881),
            .I(N__78825));
    Span4Mux_v I__17562 (
            .O(N__78874),
            .I(N__78822));
    Span4Mux_h I__17561 (
            .O(N__78871),
            .I(N__78815));
    Span4Mux_v I__17560 (
            .O(N__78866),
            .I(N__78815));
    LocalMux I__17559 (
            .O(N__78861),
            .I(N__78815));
    LocalMux I__17558 (
            .O(N__78858),
            .I(N__78812));
    LocalMux I__17557 (
            .O(N__78853),
            .I(N__78809));
    CascadeMux I__17556 (
            .O(N__78852),
            .I(N__78805));
    CascadeMux I__17555 (
            .O(N__78851),
            .I(N__78802));
    LocalMux I__17554 (
            .O(N__78848),
            .I(N__78798));
    LocalMux I__17553 (
            .O(N__78845),
            .I(N__78793));
    LocalMux I__17552 (
            .O(N__78842),
            .I(N__78793));
    Span4Mux_h I__17551 (
            .O(N__78839),
            .I(N__78788));
    Span4Mux_h I__17550 (
            .O(N__78834),
            .I(N__78788));
    Span4Mux_v I__17549 (
            .O(N__78831),
            .I(N__78785));
    Span4Mux_h I__17548 (
            .O(N__78828),
            .I(N__78778));
    Span4Mux_v I__17547 (
            .O(N__78825),
            .I(N__78778));
    Span4Mux_h I__17546 (
            .O(N__78822),
            .I(N__78778));
    Span4Mux_h I__17545 (
            .O(N__78815),
            .I(N__78775));
    Span4Mux_v I__17544 (
            .O(N__78812),
            .I(N__78770));
    Span4Mux_h I__17543 (
            .O(N__78809),
            .I(N__78770));
    InMux I__17542 (
            .O(N__78808),
            .I(N__78767));
    InMux I__17541 (
            .O(N__78805),
            .I(N__78764));
    InMux I__17540 (
            .O(N__78802),
            .I(N__78759));
    InMux I__17539 (
            .O(N__78801),
            .I(N__78759));
    Span4Mux_h I__17538 (
            .O(N__78798),
            .I(N__78752));
    Span4Mux_h I__17537 (
            .O(N__78793),
            .I(N__78752));
    Span4Mux_h I__17536 (
            .O(N__78788),
            .I(N__78752));
    Sp12to4 I__17535 (
            .O(N__78785),
            .I(N__78747));
    Sp12to4 I__17534 (
            .O(N__78778),
            .I(N__78747));
    Span4Mux_h I__17533 (
            .O(N__78775),
            .I(N__78742));
    Span4Mux_h I__17532 (
            .O(N__78770),
            .I(N__78742));
    LocalMux I__17531 (
            .O(N__78767),
            .I(rx_data_3));
    LocalMux I__17530 (
            .O(N__78764),
            .I(rx_data_3));
    LocalMux I__17529 (
            .O(N__78759),
            .I(rx_data_3));
    Odrv4 I__17528 (
            .O(N__78752),
            .I(rx_data_3));
    Odrv12 I__17527 (
            .O(N__78747),
            .I(rx_data_3));
    Odrv4 I__17526 (
            .O(N__78742),
            .I(rx_data_3));
    CascadeMux I__17525 (
            .O(N__78729),
            .I(N__78726));
    InMux I__17524 (
            .O(N__78726),
            .I(N__78719));
    InMux I__17523 (
            .O(N__78725),
            .I(N__78719));
    InMux I__17522 (
            .O(N__78724),
            .I(N__78716));
    LocalMux I__17521 (
            .O(N__78719),
            .I(N__78710));
    LocalMux I__17520 (
            .O(N__78716),
            .I(N__78710));
    CascadeMux I__17519 (
            .O(N__78715),
            .I(N__78707));
    Span4Mux_h I__17518 (
            .O(N__78710),
            .I(N__78703));
    InMux I__17517 (
            .O(N__78707),
            .I(N__78698));
    InMux I__17516 (
            .O(N__78706),
            .I(N__78698));
    Odrv4 I__17515 (
            .O(N__78703),
            .I(\c0.data_in_frame_21_3 ));
    LocalMux I__17514 (
            .O(N__78698),
            .I(\c0.data_in_frame_21_3 ));
    InMux I__17513 (
            .O(N__78693),
            .I(N__78690));
    LocalMux I__17512 (
            .O(N__78690),
            .I(N__78686));
    InMux I__17511 (
            .O(N__78689),
            .I(N__78682));
    Span4Mux_v I__17510 (
            .O(N__78686),
            .I(N__78679));
    InMux I__17509 (
            .O(N__78685),
            .I(N__78676));
    LocalMux I__17508 (
            .O(N__78682),
            .I(N__78673));
    Span4Mux_h I__17507 (
            .O(N__78679),
            .I(N__78670));
    LocalMux I__17506 (
            .O(N__78676),
            .I(N__78667));
    Span4Mux_h I__17505 (
            .O(N__78673),
            .I(N__78664));
    Odrv4 I__17504 (
            .O(N__78670),
            .I(\c0.n27890 ));
    Odrv4 I__17503 (
            .O(N__78667),
            .I(\c0.n27890 ));
    Odrv4 I__17502 (
            .O(N__78664),
            .I(\c0.n27890 ));
    CascadeMux I__17501 (
            .O(N__78657),
            .I(N__78651));
    InMux I__17500 (
            .O(N__78656),
            .I(N__78642));
    InMux I__17499 (
            .O(N__78655),
            .I(N__78642));
    InMux I__17498 (
            .O(N__78654),
            .I(N__78642));
    InMux I__17497 (
            .O(N__78651),
            .I(N__78642));
    LocalMux I__17496 (
            .O(N__78642),
            .I(N__78635));
    InMux I__17495 (
            .O(N__78641),
            .I(N__78632));
    InMux I__17494 (
            .O(N__78640),
            .I(N__78629));
    CascadeMux I__17493 (
            .O(N__78639),
            .I(N__78625));
    CascadeMux I__17492 (
            .O(N__78638),
            .I(N__78622));
    Span4Mux_v I__17491 (
            .O(N__78635),
            .I(N__78612));
    LocalMux I__17490 (
            .O(N__78632),
            .I(N__78612));
    LocalMux I__17489 (
            .O(N__78629),
            .I(N__78612));
    InMux I__17488 (
            .O(N__78628),
            .I(N__78609));
    InMux I__17487 (
            .O(N__78625),
            .I(N__78604));
    InMux I__17486 (
            .O(N__78622),
            .I(N__78604));
    InMux I__17485 (
            .O(N__78621),
            .I(N__78601));
    InMux I__17484 (
            .O(N__78620),
            .I(N__78596));
    InMux I__17483 (
            .O(N__78619),
            .I(N__78596));
    Span4Mux_v I__17482 (
            .O(N__78612),
            .I(N__78585));
    LocalMux I__17481 (
            .O(N__78609),
            .I(N__78585));
    LocalMux I__17480 (
            .O(N__78604),
            .I(N__78585));
    LocalMux I__17479 (
            .O(N__78601),
            .I(N__78585));
    LocalMux I__17478 (
            .O(N__78596),
            .I(N__78582));
    InMux I__17477 (
            .O(N__78595),
            .I(N__78576));
    InMux I__17476 (
            .O(N__78594),
            .I(N__78576));
    Span4Mux_h I__17475 (
            .O(N__78585),
            .I(N__78567));
    Span4Mux_v I__17474 (
            .O(N__78582),
            .I(N__78567));
    InMux I__17473 (
            .O(N__78581),
            .I(N__78564));
    LocalMux I__17472 (
            .O(N__78576),
            .I(N__78561));
    InMux I__17471 (
            .O(N__78575),
            .I(N__78553));
    InMux I__17470 (
            .O(N__78574),
            .I(N__78550));
    InMux I__17469 (
            .O(N__78573),
            .I(N__78545));
    InMux I__17468 (
            .O(N__78572),
            .I(N__78545));
    Span4Mux_h I__17467 (
            .O(N__78567),
            .I(N__78540));
    LocalMux I__17466 (
            .O(N__78564),
            .I(N__78540));
    Span4Mux_v I__17465 (
            .O(N__78561),
            .I(N__78537));
    InMux I__17464 (
            .O(N__78560),
            .I(N__78533));
    InMux I__17463 (
            .O(N__78559),
            .I(N__78528));
    InMux I__17462 (
            .O(N__78558),
            .I(N__78528));
    InMux I__17461 (
            .O(N__78557),
            .I(N__78525));
    InMux I__17460 (
            .O(N__78556),
            .I(N__78522));
    LocalMux I__17459 (
            .O(N__78553),
            .I(N__78517));
    LocalMux I__17458 (
            .O(N__78550),
            .I(N__78517));
    LocalMux I__17457 (
            .O(N__78545),
            .I(N__78512));
    Span4Mux_v I__17456 (
            .O(N__78540),
            .I(N__78507));
    Span4Mux_v I__17455 (
            .O(N__78537),
            .I(N__78507));
    InMux I__17454 (
            .O(N__78536),
            .I(N__78500));
    LocalMux I__17453 (
            .O(N__78533),
            .I(N__78497));
    LocalMux I__17452 (
            .O(N__78528),
            .I(N__78494));
    LocalMux I__17451 (
            .O(N__78525),
            .I(N__78491));
    LocalMux I__17450 (
            .O(N__78522),
            .I(N__78486));
    Span4Mux_h I__17449 (
            .O(N__78517),
            .I(N__78486));
    InMux I__17448 (
            .O(N__78516),
            .I(N__78481));
    InMux I__17447 (
            .O(N__78515),
            .I(N__78481));
    Span4Mux_h I__17446 (
            .O(N__78512),
            .I(N__78478));
    Sp12to4 I__17445 (
            .O(N__78507),
            .I(N__78475));
    InMux I__17444 (
            .O(N__78506),
            .I(N__78470));
    InMux I__17443 (
            .O(N__78505),
            .I(N__78470));
    InMux I__17442 (
            .O(N__78504),
            .I(N__78465));
    InMux I__17441 (
            .O(N__78503),
            .I(N__78465));
    LocalMux I__17440 (
            .O(N__78500),
            .I(N__78458));
    Span4Mux_v I__17439 (
            .O(N__78497),
            .I(N__78458));
    Span4Mux_v I__17438 (
            .O(N__78494),
            .I(N__78458));
    Span4Mux_h I__17437 (
            .O(N__78491),
            .I(N__78453));
    Span4Mux_h I__17436 (
            .O(N__78486),
            .I(N__78453));
    LocalMux I__17435 (
            .O(N__78481),
            .I(N__78448));
    Span4Mux_v I__17434 (
            .O(N__78478),
            .I(N__78448));
    Span12Mux_h I__17433 (
            .O(N__78475),
            .I(N__78445));
    LocalMux I__17432 (
            .O(N__78470),
            .I(\c0.n33224 ));
    LocalMux I__17431 (
            .O(N__78465),
            .I(\c0.n33224 ));
    Odrv4 I__17430 (
            .O(N__78458),
            .I(\c0.n33224 ));
    Odrv4 I__17429 (
            .O(N__78453),
            .I(\c0.n33224 ));
    Odrv4 I__17428 (
            .O(N__78448),
            .I(\c0.n33224 ));
    Odrv12 I__17427 (
            .O(N__78445),
            .I(\c0.n33224 ));
    CascadeMux I__17426 (
            .O(N__78432),
            .I(N__78426));
    InMux I__17425 (
            .O(N__78431),
            .I(N__78418));
    InMux I__17424 (
            .O(N__78430),
            .I(N__78415));
    InMux I__17423 (
            .O(N__78429),
            .I(N__78410));
    InMux I__17422 (
            .O(N__78426),
            .I(N__78410));
    InMux I__17421 (
            .O(N__78425),
            .I(N__78405));
    InMux I__17420 (
            .O(N__78424),
            .I(N__78405));
    InMux I__17419 (
            .O(N__78423),
            .I(N__78400));
    InMux I__17418 (
            .O(N__78422),
            .I(N__78400));
    InMux I__17417 (
            .O(N__78421),
            .I(N__78397));
    LocalMux I__17416 (
            .O(N__78418),
            .I(N__78394));
    LocalMux I__17415 (
            .O(N__78415),
            .I(N__78391));
    LocalMux I__17414 (
            .O(N__78410),
            .I(N__78388));
    LocalMux I__17413 (
            .O(N__78405),
            .I(N__78383));
    LocalMux I__17412 (
            .O(N__78400),
            .I(N__78383));
    LocalMux I__17411 (
            .O(N__78397),
            .I(N__78380));
    Span4Mux_v I__17410 (
            .O(N__78394),
            .I(N__78377));
    Span4Mux_v I__17409 (
            .O(N__78391),
            .I(N__78370));
    Span4Mux_v I__17408 (
            .O(N__78388),
            .I(N__78370));
    Span4Mux_v I__17407 (
            .O(N__78383),
            .I(N__78370));
    Span4Mux_h I__17406 (
            .O(N__78380),
            .I(N__78365));
    Span4Mux_h I__17405 (
            .O(N__78377),
            .I(N__78365));
    Odrv4 I__17404 (
            .O(N__78370),
            .I(\c0.n12_adj_4519 ));
    Odrv4 I__17403 (
            .O(N__78365),
            .I(\c0.n12_adj_4519 ));
    CascadeMux I__17402 (
            .O(N__78360),
            .I(\c0.n33224_cascade_ ));
    InMux I__17401 (
            .O(N__78357),
            .I(N__78351));
    InMux I__17400 (
            .O(N__78356),
            .I(N__78351));
    LocalMux I__17399 (
            .O(N__78351),
            .I(N__78346));
    InMux I__17398 (
            .O(N__78350),
            .I(N__78341));
    InMux I__17397 (
            .O(N__78349),
            .I(N__78341));
    Odrv12 I__17396 (
            .O(N__78346),
            .I(\c0.data_in_frame_21_4 ));
    LocalMux I__17395 (
            .O(N__78341),
            .I(\c0.data_in_frame_21_4 ));
    CascadeMux I__17394 (
            .O(N__78336),
            .I(N__78328));
    InMux I__17393 (
            .O(N__78335),
            .I(N__78322));
    InMux I__17392 (
            .O(N__78334),
            .I(N__78315));
    InMux I__17391 (
            .O(N__78333),
            .I(N__78315));
    InMux I__17390 (
            .O(N__78332),
            .I(N__78312));
    InMux I__17389 (
            .O(N__78331),
            .I(N__78309));
    InMux I__17388 (
            .O(N__78328),
            .I(N__78306));
    CascadeMux I__17387 (
            .O(N__78327),
            .I(N__78303));
    InMux I__17386 (
            .O(N__78326),
            .I(N__78300));
    CascadeMux I__17385 (
            .O(N__78325),
            .I(N__78297));
    LocalMux I__17384 (
            .O(N__78322),
            .I(N__78293));
    InMux I__17383 (
            .O(N__78321),
            .I(N__78290));
    CascadeMux I__17382 (
            .O(N__78320),
            .I(N__78282));
    LocalMux I__17381 (
            .O(N__78315),
            .I(N__78279));
    LocalMux I__17380 (
            .O(N__78312),
            .I(N__78276));
    LocalMux I__17379 (
            .O(N__78309),
            .I(N__78271));
    LocalMux I__17378 (
            .O(N__78306),
            .I(N__78271));
    InMux I__17377 (
            .O(N__78303),
            .I(N__78267));
    LocalMux I__17376 (
            .O(N__78300),
            .I(N__78264));
    InMux I__17375 (
            .O(N__78297),
            .I(N__78261));
    CascadeMux I__17374 (
            .O(N__78296),
            .I(N__78256));
    Span4Mux_v I__17373 (
            .O(N__78293),
            .I(N__78252));
    LocalMux I__17372 (
            .O(N__78290),
            .I(N__78249));
    CascadeMux I__17371 (
            .O(N__78289),
            .I(N__78246));
    InMux I__17370 (
            .O(N__78288),
            .I(N__78241));
    InMux I__17369 (
            .O(N__78287),
            .I(N__78241));
    InMux I__17368 (
            .O(N__78286),
            .I(N__78235));
    InMux I__17367 (
            .O(N__78285),
            .I(N__78235));
    InMux I__17366 (
            .O(N__78282),
            .I(N__78232));
    Span4Mux_h I__17365 (
            .O(N__78279),
            .I(N__78225));
    Span4Mux_v I__17364 (
            .O(N__78276),
            .I(N__78225));
    Span4Mux_v I__17363 (
            .O(N__78271),
            .I(N__78225));
    InMux I__17362 (
            .O(N__78270),
            .I(N__78222));
    LocalMux I__17361 (
            .O(N__78267),
            .I(N__78216));
    Span4Mux_v I__17360 (
            .O(N__78264),
            .I(N__78211));
    LocalMux I__17359 (
            .O(N__78261),
            .I(N__78211));
    InMux I__17358 (
            .O(N__78260),
            .I(N__78204));
    InMux I__17357 (
            .O(N__78259),
            .I(N__78201));
    InMux I__17356 (
            .O(N__78256),
            .I(N__78198));
    InMux I__17355 (
            .O(N__78255),
            .I(N__78195));
    Span4Mux_v I__17354 (
            .O(N__78252),
            .I(N__78190));
    Span4Mux_h I__17353 (
            .O(N__78249),
            .I(N__78190));
    InMux I__17352 (
            .O(N__78246),
            .I(N__78187));
    LocalMux I__17351 (
            .O(N__78241),
            .I(N__78184));
    InMux I__17350 (
            .O(N__78240),
            .I(N__78181));
    LocalMux I__17349 (
            .O(N__78235),
            .I(N__78176));
    LocalMux I__17348 (
            .O(N__78232),
            .I(N__78176));
    Span4Mux_h I__17347 (
            .O(N__78225),
            .I(N__78171));
    LocalMux I__17346 (
            .O(N__78222),
            .I(N__78171));
    CascadeMux I__17345 (
            .O(N__78221),
            .I(N__78168));
    InMux I__17344 (
            .O(N__78220),
            .I(N__78163));
    InMux I__17343 (
            .O(N__78219),
            .I(N__78160));
    Span4Mux_h I__17342 (
            .O(N__78216),
            .I(N__78155));
    Span4Mux_v I__17341 (
            .O(N__78211),
            .I(N__78155));
    InMux I__17340 (
            .O(N__78210),
            .I(N__78152));
    InMux I__17339 (
            .O(N__78209),
            .I(N__78145));
    InMux I__17338 (
            .O(N__78208),
            .I(N__78145));
    InMux I__17337 (
            .O(N__78207),
            .I(N__78145));
    LocalMux I__17336 (
            .O(N__78204),
            .I(N__78140));
    LocalMux I__17335 (
            .O(N__78201),
            .I(N__78140));
    LocalMux I__17334 (
            .O(N__78198),
            .I(N__78136));
    LocalMux I__17333 (
            .O(N__78195),
            .I(N__78131));
    Span4Mux_h I__17332 (
            .O(N__78190),
            .I(N__78131));
    LocalMux I__17331 (
            .O(N__78187),
            .I(N__78124));
    Span4Mux_h I__17330 (
            .O(N__78184),
            .I(N__78124));
    LocalMux I__17329 (
            .O(N__78181),
            .I(N__78124));
    Span12Mux_v I__17328 (
            .O(N__78176),
            .I(N__78119));
    Sp12to4 I__17327 (
            .O(N__78171),
            .I(N__78119));
    InMux I__17326 (
            .O(N__78168),
            .I(N__78116));
    InMux I__17325 (
            .O(N__78167),
            .I(N__78111));
    InMux I__17324 (
            .O(N__78166),
            .I(N__78111));
    LocalMux I__17323 (
            .O(N__78163),
            .I(N__78104));
    LocalMux I__17322 (
            .O(N__78160),
            .I(N__78104));
    Sp12to4 I__17321 (
            .O(N__78155),
            .I(N__78104));
    LocalMux I__17320 (
            .O(N__78152),
            .I(N__78097));
    LocalMux I__17319 (
            .O(N__78145),
            .I(N__78097));
    Span12Mux_v I__17318 (
            .O(N__78140),
            .I(N__78097));
    InMux I__17317 (
            .O(N__78139),
            .I(N__78094));
    Span4Mux_h I__17316 (
            .O(N__78136),
            .I(N__78091));
    Span4Mux_h I__17315 (
            .O(N__78131),
            .I(N__78088));
    Sp12to4 I__17314 (
            .O(N__78124),
            .I(N__78083));
    Span12Mux_h I__17313 (
            .O(N__78119),
            .I(N__78083));
    LocalMux I__17312 (
            .O(N__78116),
            .I(N__78076));
    LocalMux I__17311 (
            .O(N__78111),
            .I(N__78076));
    Span12Mux_s7_v I__17310 (
            .O(N__78104),
            .I(N__78076));
    Span12Mux_h I__17309 (
            .O(N__78097),
            .I(N__78073));
    LocalMux I__17308 (
            .O(N__78094),
            .I(\c0.n9_adj_4628 ));
    Odrv4 I__17307 (
            .O(N__78091),
            .I(\c0.n9_adj_4628 ));
    Odrv4 I__17306 (
            .O(N__78088),
            .I(\c0.n9_adj_4628 ));
    Odrv12 I__17305 (
            .O(N__78083),
            .I(\c0.n9_adj_4628 ));
    Odrv12 I__17304 (
            .O(N__78076),
            .I(\c0.n9_adj_4628 ));
    Odrv12 I__17303 (
            .O(N__78073),
            .I(\c0.n9_adj_4628 ));
    InMux I__17302 (
            .O(N__78060),
            .I(N__78057));
    LocalMux I__17301 (
            .O(N__78057),
            .I(N__78054));
    Span4Mux_h I__17300 (
            .O(N__78054),
            .I(N__78051));
    Odrv4 I__17299 (
            .O(N__78051),
            .I(n2321));
    CascadeMux I__17298 (
            .O(N__78048),
            .I(N__78045));
    InMux I__17297 (
            .O(N__78045),
            .I(N__78042));
    LocalMux I__17296 (
            .O(N__78042),
            .I(N__78039));
    Span4Mux_v I__17295 (
            .O(N__78039),
            .I(N__78032));
    InMux I__17294 (
            .O(N__78038),
            .I(N__78029));
    InMux I__17293 (
            .O(N__78037),
            .I(N__78026));
    InMux I__17292 (
            .O(N__78036),
            .I(N__78021));
    InMux I__17291 (
            .O(N__78035),
            .I(N__78017));
    Sp12to4 I__17290 (
            .O(N__78032),
            .I(N__78012));
    LocalMux I__17289 (
            .O(N__78029),
            .I(N__78012));
    LocalMux I__17288 (
            .O(N__78026),
            .I(N__78009));
    InMux I__17287 (
            .O(N__78025),
            .I(N__78004));
    InMux I__17286 (
            .O(N__78024),
            .I(N__78004));
    LocalMux I__17285 (
            .O(N__78021),
            .I(N__78001));
    InMux I__17284 (
            .O(N__78020),
            .I(N__77998));
    LocalMux I__17283 (
            .O(N__78017),
            .I(N__77995));
    Span12Mux_h I__17282 (
            .O(N__78012),
            .I(N__77992));
    Span4Mux_v I__17281 (
            .O(N__78009),
            .I(N__77985));
    LocalMux I__17280 (
            .O(N__78004),
            .I(N__77985));
    Span4Mux_h I__17279 (
            .O(N__78001),
            .I(N__77985));
    LocalMux I__17278 (
            .O(N__77998),
            .I(encoder0_position_24));
    Odrv12 I__17277 (
            .O(N__77995),
            .I(encoder0_position_24));
    Odrv12 I__17276 (
            .O(N__77992),
            .I(encoder0_position_24));
    Odrv4 I__17275 (
            .O(N__77985),
            .I(encoder0_position_24));
    InMux I__17274 (
            .O(N__77976),
            .I(N__77973));
    LocalMux I__17273 (
            .O(N__77973),
            .I(N__77970));
    Span4Mux_v I__17272 (
            .O(N__77970),
            .I(N__77967));
    Span4Mux_h I__17271 (
            .O(N__77967),
            .I(N__77964));
    Odrv4 I__17270 (
            .O(N__77964),
            .I(n2340));
    InMux I__17269 (
            .O(N__77961),
            .I(N__77958));
    LocalMux I__17268 (
            .O(N__77958),
            .I(N__77955));
    Odrv12 I__17267 (
            .O(N__77955),
            .I(n2333));
    CascadeMux I__17266 (
            .O(N__77952),
            .I(N__77949));
    InMux I__17265 (
            .O(N__77949),
            .I(N__77944));
    InMux I__17264 (
            .O(N__77948),
            .I(N__77940));
    InMux I__17263 (
            .O(N__77947),
            .I(N__77937));
    LocalMux I__17262 (
            .O(N__77944),
            .I(N__77933));
    CascadeMux I__17261 (
            .O(N__77943),
            .I(N__77930));
    LocalMux I__17260 (
            .O(N__77940),
            .I(N__77925));
    LocalMux I__17259 (
            .O(N__77937),
            .I(N__77925));
    InMux I__17258 (
            .O(N__77936),
            .I(N__77922));
    Span4Mux_v I__17257 (
            .O(N__77933),
            .I(N__77919));
    InMux I__17256 (
            .O(N__77930),
            .I(N__77916));
    Span12Mux_h I__17255 (
            .O(N__77925),
            .I(N__77913));
    LocalMux I__17254 (
            .O(N__77922),
            .I(encoder1_position_29));
    Odrv4 I__17253 (
            .O(N__77919),
            .I(encoder1_position_29));
    LocalMux I__17252 (
            .O(N__77916),
            .I(encoder1_position_29));
    Odrv12 I__17251 (
            .O(N__77913),
            .I(encoder1_position_29));
    InMux I__17250 (
            .O(N__77904),
            .I(N__77896));
    InMux I__17249 (
            .O(N__77903),
            .I(N__77896));
    InMux I__17248 (
            .O(N__77902),
            .I(N__77893));
    InMux I__17247 (
            .O(N__77901),
            .I(N__77890));
    LocalMux I__17246 (
            .O(N__77896),
            .I(N__77883));
    LocalMux I__17245 (
            .O(N__77893),
            .I(N__77883));
    LocalMux I__17244 (
            .O(N__77890),
            .I(N__77883));
    Span4Mux_v I__17243 (
            .O(N__77883),
            .I(N__77880));
    Odrv4 I__17242 (
            .O(N__77880),
            .I(\c0.n18214 ));
    CascadeMux I__17241 (
            .O(N__77877),
            .I(N__77874));
    InMux I__17240 (
            .O(N__77874),
            .I(N__77870));
    CascadeMux I__17239 (
            .O(N__77873),
            .I(N__77867));
    LocalMux I__17238 (
            .O(N__77870),
            .I(N__77863));
    InMux I__17237 (
            .O(N__77867),
            .I(N__77860));
    InMux I__17236 (
            .O(N__77866),
            .I(N__77857));
    Span4Mux_v I__17235 (
            .O(N__77863),
            .I(N__77853));
    LocalMux I__17234 (
            .O(N__77860),
            .I(N__77850));
    LocalMux I__17233 (
            .O(N__77857),
            .I(N__77847));
    InMux I__17232 (
            .O(N__77856),
            .I(N__77844));
    Span4Mux_h I__17231 (
            .O(N__77853),
            .I(N__77841));
    Span4Mux_h I__17230 (
            .O(N__77850),
            .I(N__77838));
    Span4Mux_v I__17229 (
            .O(N__77847),
            .I(N__77835));
    LocalMux I__17228 (
            .O(N__77844),
            .I(encoder1_position_17));
    Odrv4 I__17227 (
            .O(N__77841),
            .I(encoder1_position_17));
    Odrv4 I__17226 (
            .O(N__77838),
            .I(encoder1_position_17));
    Odrv4 I__17225 (
            .O(N__77835),
            .I(encoder1_position_17));
    CascadeMux I__17224 (
            .O(N__77826),
            .I(N__77822));
    InMux I__17223 (
            .O(N__77825),
            .I(N__77816));
    InMux I__17222 (
            .O(N__77822),
            .I(N__77813));
    InMux I__17221 (
            .O(N__77821),
            .I(N__77810));
    InMux I__17220 (
            .O(N__77820),
            .I(N__77807));
    InMux I__17219 (
            .O(N__77819),
            .I(N__77804));
    LocalMux I__17218 (
            .O(N__77816),
            .I(N__77801));
    LocalMux I__17217 (
            .O(N__77813),
            .I(N__77798));
    LocalMux I__17216 (
            .O(N__77810),
            .I(N__77795));
    LocalMux I__17215 (
            .O(N__77807),
            .I(N__77792));
    LocalMux I__17214 (
            .O(N__77804),
            .I(encoder0_position_13));
    Odrv12 I__17213 (
            .O(N__77801),
            .I(encoder0_position_13));
    Odrv4 I__17212 (
            .O(N__77798),
            .I(encoder0_position_13));
    Odrv4 I__17211 (
            .O(N__77795),
            .I(encoder0_position_13));
    Odrv4 I__17210 (
            .O(N__77792),
            .I(encoder0_position_13));
    InMux I__17209 (
            .O(N__77781),
            .I(N__77778));
    LocalMux I__17208 (
            .O(N__77778),
            .I(N__77775));
    Odrv4 I__17207 (
            .O(N__77775),
            .I(\c0.n33896 ));
    CascadeMux I__17206 (
            .O(N__77772),
            .I(\c0.n33896_cascade_ ));
    InMux I__17205 (
            .O(N__77769),
            .I(N__77766));
    LocalMux I__17204 (
            .O(N__77766),
            .I(N__77763));
    Odrv4 I__17203 (
            .O(N__77763),
            .I(\c0.n6_adj_4541 ));
    InMux I__17202 (
            .O(N__77760),
            .I(N__77756));
    InMux I__17201 (
            .O(N__77759),
            .I(N__77753));
    LocalMux I__17200 (
            .O(N__77756),
            .I(N__77750));
    LocalMux I__17199 (
            .O(N__77753),
            .I(N__77747));
    Span4Mux_h I__17198 (
            .O(N__77750),
            .I(N__77744));
    Span4Mux_h I__17197 (
            .O(N__77747),
            .I(N__77741));
    Odrv4 I__17196 (
            .O(N__77744),
            .I(\c0.n18892 ));
    Odrv4 I__17195 (
            .O(N__77741),
            .I(\c0.n18892 ));
    CascadeMux I__17194 (
            .O(N__77736),
            .I(\c0.n33360_cascade_ ));
    InMux I__17193 (
            .O(N__77733),
            .I(N__77728));
    InMux I__17192 (
            .O(N__77732),
            .I(N__77723));
    InMux I__17191 (
            .O(N__77731),
            .I(N__77723));
    LocalMux I__17190 (
            .O(N__77728),
            .I(\c0.n18181 ));
    LocalMux I__17189 (
            .O(N__77723),
            .I(\c0.n18181 ));
    InMux I__17188 (
            .O(N__77718),
            .I(N__77715));
    LocalMux I__17187 (
            .O(N__77715),
            .I(\c0.n18740 ));
    InMux I__17186 (
            .O(N__77712),
            .I(N__77706));
    InMux I__17185 (
            .O(N__77711),
            .I(N__77706));
    LocalMux I__17184 (
            .O(N__77706),
            .I(\c0.data_out_frame_29__7__N_734 ));
    CascadeMux I__17183 (
            .O(N__77703),
            .I(\c0.n33425_cascade_ ));
    CascadeMux I__17182 (
            .O(N__77700),
            .I(N__77696));
    CascadeMux I__17181 (
            .O(N__77699),
            .I(N__77693));
    InMux I__17180 (
            .O(N__77696),
            .I(N__77688));
    InMux I__17179 (
            .O(N__77693),
            .I(N__77685));
    InMux I__17178 (
            .O(N__77692),
            .I(N__77682));
    InMux I__17177 (
            .O(N__77691),
            .I(N__77679));
    LocalMux I__17176 (
            .O(N__77688),
            .I(N__77673));
    LocalMux I__17175 (
            .O(N__77685),
            .I(N__77670));
    LocalMux I__17174 (
            .O(N__77682),
            .I(N__77667));
    LocalMux I__17173 (
            .O(N__77679),
            .I(N__77664));
    InMux I__17172 (
            .O(N__77678),
            .I(N__77659));
    InMux I__17171 (
            .O(N__77677),
            .I(N__77659));
    InMux I__17170 (
            .O(N__77676),
            .I(N__77656));
    Span4Mux_h I__17169 (
            .O(N__77673),
            .I(N__77651));
    Span4Mux_h I__17168 (
            .O(N__77670),
            .I(N__77651));
    Span12Mux_v I__17167 (
            .O(N__77667),
            .I(N__77648));
    Span4Mux_h I__17166 (
            .O(N__77664),
            .I(N__77645));
    LocalMux I__17165 (
            .O(N__77659),
            .I(N__77642));
    LocalMux I__17164 (
            .O(N__77656),
            .I(encoder0_position_18));
    Odrv4 I__17163 (
            .O(N__77651),
            .I(encoder0_position_18));
    Odrv12 I__17162 (
            .O(N__77648),
            .I(encoder0_position_18));
    Odrv4 I__17161 (
            .O(N__77645),
            .I(encoder0_position_18));
    Odrv4 I__17160 (
            .O(N__77642),
            .I(encoder0_position_18));
    InMux I__17159 (
            .O(N__77631),
            .I(N__77623));
    InMux I__17158 (
            .O(N__77630),
            .I(N__77620));
    InMux I__17157 (
            .O(N__77629),
            .I(N__77613));
    InMux I__17156 (
            .O(N__77628),
            .I(N__77613));
    InMux I__17155 (
            .O(N__77627),
            .I(N__77610));
    InMux I__17154 (
            .O(N__77626),
            .I(N__77607));
    LocalMux I__17153 (
            .O(N__77623),
            .I(N__77604));
    LocalMux I__17152 (
            .O(N__77620),
            .I(N__77601));
    InMux I__17151 (
            .O(N__77619),
            .I(N__77596));
    InMux I__17150 (
            .O(N__77618),
            .I(N__77596));
    LocalMux I__17149 (
            .O(N__77613),
            .I(N__77593));
    LocalMux I__17148 (
            .O(N__77610),
            .I(N__77588));
    LocalMux I__17147 (
            .O(N__77607),
            .I(N__77588));
    Span4Mux_v I__17146 (
            .O(N__77604),
            .I(N__77585));
    Span4Mux_v I__17145 (
            .O(N__77601),
            .I(N__77582));
    LocalMux I__17144 (
            .O(N__77596),
            .I(N__77579));
    Span4Mux_h I__17143 (
            .O(N__77593),
            .I(N__77576));
    Span4Mux_h I__17142 (
            .O(N__77588),
            .I(N__77573));
    Span4Mux_v I__17141 (
            .O(N__77585),
            .I(N__77568));
    Span4Mux_v I__17140 (
            .O(N__77582),
            .I(N__77568));
    Odrv12 I__17139 (
            .O(N__77579),
            .I(n35693));
    Odrv4 I__17138 (
            .O(N__77576),
            .I(n35693));
    Odrv4 I__17137 (
            .O(N__77573),
            .I(n35693));
    Odrv4 I__17136 (
            .O(N__77568),
            .I(n35693));
    CascadeMux I__17135 (
            .O(N__77559),
            .I(N__77555));
    InMux I__17134 (
            .O(N__77558),
            .I(N__77550));
    InMux I__17133 (
            .O(N__77555),
            .I(N__77547));
    InMux I__17132 (
            .O(N__77554),
            .I(N__77544));
    InMux I__17131 (
            .O(N__77553),
            .I(N__77539));
    LocalMux I__17130 (
            .O(N__77550),
            .I(N__77536));
    LocalMux I__17129 (
            .O(N__77547),
            .I(N__77533));
    LocalMux I__17128 (
            .O(N__77544),
            .I(N__77530));
    InMux I__17127 (
            .O(N__77543),
            .I(N__77525));
    InMux I__17126 (
            .O(N__77542),
            .I(N__77525));
    LocalMux I__17125 (
            .O(N__77539),
            .I(N__77522));
    Span4Mux_h I__17124 (
            .O(N__77536),
            .I(N__77519));
    Odrv4 I__17123 (
            .O(N__77533),
            .I(control_mode_4));
    Odrv4 I__17122 (
            .O(N__77530),
            .I(control_mode_4));
    LocalMux I__17121 (
            .O(N__77525),
            .I(control_mode_4));
    Odrv4 I__17120 (
            .O(N__77522),
            .I(control_mode_4));
    Odrv4 I__17119 (
            .O(N__77519),
            .I(control_mode_4));
    InMux I__17118 (
            .O(N__77508),
            .I(N__77505));
    LocalMux I__17117 (
            .O(N__77505),
            .I(N__77501));
    InMux I__17116 (
            .O(N__77504),
            .I(N__77496));
    Span4Mux_v I__17115 (
            .O(N__77501),
            .I(N__77493));
    InMux I__17114 (
            .O(N__77500),
            .I(N__77490));
    CascadeMux I__17113 (
            .O(N__77499),
            .I(N__77486));
    LocalMux I__17112 (
            .O(N__77496),
            .I(N__77483));
    Span4Mux_h I__17111 (
            .O(N__77493),
            .I(N__77478));
    LocalMux I__17110 (
            .O(N__77490),
            .I(N__77478));
    InMux I__17109 (
            .O(N__77489),
            .I(N__77475));
    InMux I__17108 (
            .O(N__77486),
            .I(N__77472));
    Span4Mux_v I__17107 (
            .O(N__77483),
            .I(N__77467));
    Span4Mux_h I__17106 (
            .O(N__77478),
            .I(N__77467));
    LocalMux I__17105 (
            .O(N__77475),
            .I(encoder1_position_27));
    LocalMux I__17104 (
            .O(N__77472),
            .I(encoder1_position_27));
    Odrv4 I__17103 (
            .O(N__77467),
            .I(encoder1_position_27));
    CascadeMux I__17102 (
            .O(N__77460),
            .I(N__77457));
    InMux I__17101 (
            .O(N__77457),
            .I(N__77454));
    LocalMux I__17100 (
            .O(N__77454),
            .I(N__77450));
    CascadeMux I__17099 (
            .O(N__77453),
            .I(N__77447));
    Span4Mux_h I__17098 (
            .O(N__77450),
            .I(N__77444));
    InMux I__17097 (
            .O(N__77447),
            .I(N__77441));
    Span4Mux_v I__17096 (
            .O(N__77444),
            .I(N__77436));
    LocalMux I__17095 (
            .O(N__77441),
            .I(N__77436));
    Span4Mux_v I__17094 (
            .O(N__77436),
            .I(N__77432));
    InMux I__17093 (
            .O(N__77435),
            .I(N__77429));
    Span4Mux_h I__17092 (
            .O(N__77432),
            .I(N__77424));
    LocalMux I__17091 (
            .O(N__77429),
            .I(N__77421));
    InMux I__17090 (
            .O(N__77428),
            .I(N__77416));
    InMux I__17089 (
            .O(N__77427),
            .I(N__77416));
    Odrv4 I__17088 (
            .O(N__77424),
            .I(encoder0_position_9));
    Odrv4 I__17087 (
            .O(N__77421),
            .I(encoder0_position_9));
    LocalMux I__17086 (
            .O(N__77416),
            .I(encoder0_position_9));
    InMux I__17085 (
            .O(N__77409),
            .I(N__77405));
    InMux I__17084 (
            .O(N__77408),
            .I(N__77402));
    LocalMux I__17083 (
            .O(N__77405),
            .I(N__77399));
    LocalMux I__17082 (
            .O(N__77402),
            .I(\c0.n17510 ));
    Odrv4 I__17081 (
            .O(N__77399),
            .I(\c0.n17510 ));
    CascadeMux I__17080 (
            .O(N__77394),
            .I(N__77391));
    InMux I__17079 (
            .O(N__77391),
            .I(N__77382));
    InMux I__17078 (
            .O(N__77390),
            .I(N__77382));
    InMux I__17077 (
            .O(N__77389),
            .I(N__77382));
    LocalMux I__17076 (
            .O(N__77382),
            .I(N__77379));
    Span4Mux_v I__17075 (
            .O(N__77379),
            .I(N__77376));
    Odrv4 I__17074 (
            .O(N__77376),
            .I(\c0.n33393 ));
    CascadeMux I__17073 (
            .O(N__77373),
            .I(N__77370));
    InMux I__17072 (
            .O(N__77370),
            .I(N__77367));
    LocalMux I__17071 (
            .O(N__77367),
            .I(N__77363));
    InMux I__17070 (
            .O(N__77366),
            .I(N__77360));
    Span4Mux_h I__17069 (
            .O(N__77363),
            .I(N__77357));
    LocalMux I__17068 (
            .O(N__77360),
            .I(\c0.n33280 ));
    Odrv4 I__17067 (
            .O(N__77357),
            .I(\c0.n33280 ));
    CascadeMux I__17066 (
            .O(N__77352),
            .I(N__77348));
    InMux I__17065 (
            .O(N__77351),
            .I(N__77345));
    InMux I__17064 (
            .O(N__77348),
            .I(N__77340));
    LocalMux I__17063 (
            .O(N__77345),
            .I(N__77337));
    InMux I__17062 (
            .O(N__77344),
            .I(N__77333));
    InMux I__17061 (
            .O(N__77343),
            .I(N__77330));
    LocalMux I__17060 (
            .O(N__77340),
            .I(N__77325));
    Span4Mux_h I__17059 (
            .O(N__77337),
            .I(N__77325));
    InMux I__17058 (
            .O(N__77336),
            .I(N__77322));
    LocalMux I__17057 (
            .O(N__77333),
            .I(encoder1_position_28));
    LocalMux I__17056 (
            .O(N__77330),
            .I(encoder1_position_28));
    Odrv4 I__17055 (
            .O(N__77325),
            .I(encoder1_position_28));
    LocalMux I__17054 (
            .O(N__77322),
            .I(encoder1_position_28));
    InMux I__17053 (
            .O(N__77313),
            .I(N__77307));
    InMux I__17052 (
            .O(N__77312),
            .I(N__77307));
    LocalMux I__17051 (
            .O(N__77307),
            .I(N__77304));
    Span4Mux_h I__17050 (
            .O(N__77304),
            .I(N__77301));
    Odrv4 I__17049 (
            .O(N__77301),
            .I(\c0.n33496 ));
    CascadeMux I__17048 (
            .O(N__77298),
            .I(\c0.n33496_cascade_ ));
    CascadeMux I__17047 (
            .O(N__77295),
            .I(N__77291));
    InMux I__17046 (
            .O(N__77294),
            .I(N__77288));
    InMux I__17045 (
            .O(N__77291),
            .I(N__77282));
    LocalMux I__17044 (
            .O(N__77288),
            .I(N__77278));
    InMux I__17043 (
            .O(N__77287),
            .I(N__77273));
    InMux I__17042 (
            .O(N__77286),
            .I(N__77273));
    InMux I__17041 (
            .O(N__77285),
            .I(N__77269));
    LocalMux I__17040 (
            .O(N__77282),
            .I(N__77266));
    InMux I__17039 (
            .O(N__77281),
            .I(N__77263));
    Span4Mux_v I__17038 (
            .O(N__77278),
            .I(N__77260));
    LocalMux I__17037 (
            .O(N__77273),
            .I(N__77257));
    InMux I__17036 (
            .O(N__77272),
            .I(N__77254));
    LocalMux I__17035 (
            .O(N__77269),
            .I(encoder1_position_14));
    Odrv12 I__17034 (
            .O(N__77266),
            .I(encoder1_position_14));
    LocalMux I__17033 (
            .O(N__77263),
            .I(encoder1_position_14));
    Odrv4 I__17032 (
            .O(N__77260),
            .I(encoder1_position_14));
    Odrv12 I__17031 (
            .O(N__77257),
            .I(encoder1_position_14));
    LocalMux I__17030 (
            .O(N__77254),
            .I(encoder1_position_14));
    CascadeMux I__17029 (
            .O(N__77241),
            .I(\c0.n6_adj_4544_cascade_ ));
    InMux I__17028 (
            .O(N__77238),
            .I(N__77235));
    LocalMux I__17027 (
            .O(N__77235),
            .I(N__77232));
    Span4Mux_h I__17026 (
            .O(N__77232),
            .I(N__77229));
    Odrv4 I__17025 (
            .O(N__77229),
            .I(n36176));
    InMux I__17024 (
            .O(N__77226),
            .I(N__77223));
    LocalMux I__17023 (
            .O(N__77223),
            .I(N__77220));
    Span4Mux_v I__17022 (
            .O(N__77220),
            .I(N__77217));
    Odrv4 I__17021 (
            .O(N__77217),
            .I(n36099));
    CascadeMux I__17020 (
            .O(N__77214),
            .I(N__77211));
    InMux I__17019 (
            .O(N__77211),
            .I(N__77207));
    InMux I__17018 (
            .O(N__77210),
            .I(N__77204));
    LocalMux I__17017 (
            .O(N__77207),
            .I(N__77197));
    LocalMux I__17016 (
            .O(N__77204),
            .I(N__77197));
    InMux I__17015 (
            .O(N__77203),
            .I(N__77194));
    InMux I__17014 (
            .O(N__77202),
            .I(N__77191));
    Span4Mux_h I__17013 (
            .O(N__77197),
            .I(N__77186));
    LocalMux I__17012 (
            .O(N__77194),
            .I(N__77186));
    LocalMux I__17011 (
            .O(N__77191),
            .I(N__77181));
    Span4Mux_h I__17010 (
            .O(N__77186),
            .I(N__77178));
    InMux I__17009 (
            .O(N__77185),
            .I(N__77175));
    InMux I__17008 (
            .O(N__77184),
            .I(N__77172));
    Span12Mux_h I__17007 (
            .O(N__77181),
            .I(N__77169));
    Span4Mux_v I__17006 (
            .O(N__77178),
            .I(N__77166));
    LocalMux I__17005 (
            .O(N__77175),
            .I(data_in_frame_1_7));
    LocalMux I__17004 (
            .O(N__77172),
            .I(data_in_frame_1_7));
    Odrv12 I__17003 (
            .O(N__77169),
            .I(data_in_frame_1_7));
    Odrv4 I__17002 (
            .O(N__77166),
            .I(data_in_frame_1_7));
    InMux I__17001 (
            .O(N__77157),
            .I(N__77154));
    LocalMux I__17000 (
            .O(N__77154),
            .I(N__77151));
    Span4Mux_h I__16999 (
            .O(N__77151),
            .I(N__77148));
    Odrv4 I__16998 (
            .O(N__77148),
            .I(n2334));
    CascadeMux I__16997 (
            .O(N__77145),
            .I(N__77142));
    InMux I__16996 (
            .O(N__77142),
            .I(N__77138));
    CascadeMux I__16995 (
            .O(N__77141),
            .I(N__77135));
    LocalMux I__16994 (
            .O(N__77138),
            .I(N__77132));
    InMux I__16993 (
            .O(N__77135),
            .I(N__77129));
    Span4Mux_v I__16992 (
            .O(N__77132),
            .I(N__77125));
    LocalMux I__16991 (
            .O(N__77129),
            .I(N__77122));
    InMux I__16990 (
            .O(N__77128),
            .I(N__77118));
    Span4Mux_h I__16989 (
            .O(N__77125),
            .I(N__77113));
    Span4Mux_h I__16988 (
            .O(N__77122),
            .I(N__77113));
    InMux I__16987 (
            .O(N__77121),
            .I(N__77110));
    LocalMux I__16986 (
            .O(N__77118),
            .I(encoder0_position_11));
    Odrv4 I__16985 (
            .O(N__77113),
            .I(encoder0_position_11));
    LocalMux I__16984 (
            .O(N__77110),
            .I(encoder0_position_11));
    InMux I__16983 (
            .O(N__77103),
            .I(N__77100));
    LocalMux I__16982 (
            .O(N__77100),
            .I(N__77097));
    Span4Mux_h I__16981 (
            .O(N__77097),
            .I(N__77091));
    InMux I__16980 (
            .O(N__77096),
            .I(N__77084));
    InMux I__16979 (
            .O(N__77095),
            .I(N__77084));
    InMux I__16978 (
            .O(N__77094),
            .I(N__77084));
    Span4Mux_h I__16977 (
            .O(N__77091),
            .I(N__77076));
    LocalMux I__16976 (
            .O(N__77084),
            .I(N__77076));
    InMux I__16975 (
            .O(N__77083),
            .I(N__77073));
    InMux I__16974 (
            .O(N__77082),
            .I(N__77068));
    InMux I__16973 (
            .O(N__77081),
            .I(N__77068));
    Span4Mux_h I__16972 (
            .O(N__77076),
            .I(N__77065));
    LocalMux I__16971 (
            .O(N__77073),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__16970 (
            .O(N__77068),
            .I(\c0.rx.r_Clock_Count_4 ));
    Odrv4 I__16969 (
            .O(N__77065),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__16968 (
            .O(N__77058),
            .I(N__77055));
    LocalMux I__16967 (
            .O(N__77055),
            .I(N__77052));
    Span4Mux_v I__16966 (
            .O(N__77052),
            .I(N__77049));
    Sp12to4 I__16965 (
            .O(N__77049),
            .I(N__77043));
    InMux I__16964 (
            .O(N__77048),
            .I(N__77036));
    InMux I__16963 (
            .O(N__77047),
            .I(N__77036));
    InMux I__16962 (
            .O(N__77046),
            .I(N__77036));
    Odrv12 I__16961 (
            .O(N__77043),
            .I(\c0.rx.n18092 ));
    LocalMux I__16960 (
            .O(N__77036),
            .I(\c0.rx.n18092 ));
    InMux I__16959 (
            .O(N__77031),
            .I(N__77027));
    CascadeMux I__16958 (
            .O(N__77030),
            .I(N__77022));
    LocalMux I__16957 (
            .O(N__77027),
            .I(N__77017));
    InMux I__16956 (
            .O(N__77026),
            .I(N__77014));
    InMux I__16955 (
            .O(N__77025),
            .I(N__77011));
    InMux I__16954 (
            .O(N__77022),
            .I(N__77004));
    InMux I__16953 (
            .O(N__77021),
            .I(N__77004));
    InMux I__16952 (
            .O(N__77020),
            .I(N__77004));
    Odrv12 I__16951 (
            .O(N__77017),
            .I(\c0.rx.n33168 ));
    LocalMux I__16950 (
            .O(N__77014),
            .I(\c0.rx.n33168 ));
    LocalMux I__16949 (
            .O(N__77011),
            .I(\c0.rx.n33168 ));
    LocalMux I__16948 (
            .O(N__77004),
            .I(\c0.rx.n33168 ));
    InMux I__16947 (
            .O(N__76995),
            .I(N__76985));
    InMux I__16946 (
            .O(N__76994),
            .I(N__76985));
    InMux I__16945 (
            .O(N__76993),
            .I(N__76982));
    InMux I__16944 (
            .O(N__76992),
            .I(N__76976));
    InMux I__16943 (
            .O(N__76991),
            .I(N__76971));
    InMux I__16942 (
            .O(N__76990),
            .I(N__76971));
    LocalMux I__16941 (
            .O(N__76985),
            .I(N__76968));
    LocalMux I__16940 (
            .O(N__76982),
            .I(N__76965));
    InMux I__16939 (
            .O(N__76981),
            .I(N__76958));
    InMux I__16938 (
            .O(N__76980),
            .I(N__76958));
    InMux I__16937 (
            .O(N__76979),
            .I(N__76958));
    LocalMux I__16936 (
            .O(N__76976),
            .I(N__76955));
    LocalMux I__16935 (
            .O(N__76971),
            .I(N__76952));
    Span4Mux_v I__16934 (
            .O(N__76968),
            .I(N__76945));
    Span4Mux_h I__16933 (
            .O(N__76965),
            .I(N__76945));
    LocalMux I__16932 (
            .O(N__76958),
            .I(N__76945));
    Span4Mux_h I__16931 (
            .O(N__76955),
            .I(N__76942));
    Span12Mux_h I__16930 (
            .O(N__76952),
            .I(N__76937));
    Sp12to4 I__16929 (
            .O(N__76945),
            .I(N__76937));
    Odrv4 I__16928 (
            .O(N__76942),
            .I(r_SM_Main_2));
    Odrv12 I__16927 (
            .O(N__76937),
            .I(r_SM_Main_2));
    SRMux I__16926 (
            .O(N__76932),
            .I(N__76929));
    LocalMux I__16925 (
            .O(N__76929),
            .I(N__76926));
    Span4Mux_v I__16924 (
            .O(N__76926),
            .I(N__76923));
    Span4Mux_h I__16923 (
            .O(N__76923),
            .I(N__76920));
    Sp12to4 I__16922 (
            .O(N__76920),
            .I(N__76917));
    Odrv12 I__16921 (
            .O(N__76917),
            .I(\c0.rx.n34953 ));
    CascadeMux I__16920 (
            .O(N__76914),
            .I(N__76911));
    InMux I__16919 (
            .O(N__76911),
            .I(N__76907));
    InMux I__16918 (
            .O(N__76910),
            .I(N__76901));
    LocalMux I__16917 (
            .O(N__76907),
            .I(N__76898));
    InMux I__16916 (
            .O(N__76906),
            .I(N__76895));
    InMux I__16915 (
            .O(N__76905),
            .I(N__76890));
    InMux I__16914 (
            .O(N__76904),
            .I(N__76890));
    LocalMux I__16913 (
            .O(N__76901),
            .I(N__76886));
    Span4Mux_h I__16912 (
            .O(N__76898),
            .I(N__76881));
    LocalMux I__16911 (
            .O(N__76895),
            .I(N__76881));
    LocalMux I__16910 (
            .O(N__76890),
            .I(N__76878));
    InMux I__16909 (
            .O(N__76889),
            .I(N__76875));
    Span4Mux_v I__16908 (
            .O(N__76886),
            .I(N__76870));
    Span4Mux_v I__16907 (
            .O(N__76881),
            .I(N__76870));
    Span4Mux_h I__16906 (
            .O(N__76878),
            .I(N__76867));
    LocalMux I__16905 (
            .O(N__76875),
            .I(encoder0_position_31));
    Odrv4 I__16904 (
            .O(N__76870),
            .I(encoder0_position_31));
    Odrv4 I__16903 (
            .O(N__76867),
            .I(encoder0_position_31));
    CascadeMux I__16902 (
            .O(N__76860),
            .I(N__76857));
    InMux I__16901 (
            .O(N__76857),
            .I(N__76852));
    InMux I__16900 (
            .O(N__76856),
            .I(N__76847));
    InMux I__16899 (
            .O(N__76855),
            .I(N__76847));
    LocalMux I__16898 (
            .O(N__76852),
            .I(N__76843));
    LocalMux I__16897 (
            .O(N__76847),
            .I(N__76840));
    InMux I__16896 (
            .O(N__76846),
            .I(N__76836));
    Span4Mux_h I__16895 (
            .O(N__76843),
            .I(N__76831));
    Span4Mux_h I__16894 (
            .O(N__76840),
            .I(N__76831));
    InMux I__16893 (
            .O(N__76839),
            .I(N__76828));
    LocalMux I__16892 (
            .O(N__76836),
            .I(N__76825));
    Span4Mux_v I__16891 (
            .O(N__76831),
            .I(N__76822));
    LocalMux I__16890 (
            .O(N__76828),
            .I(encoder0_position_30));
    Odrv4 I__16889 (
            .O(N__76825),
            .I(encoder0_position_30));
    Odrv4 I__16888 (
            .O(N__76822),
            .I(encoder0_position_30));
    CascadeMux I__16887 (
            .O(N__76815),
            .I(N__76812));
    InMux I__16886 (
            .O(N__76812),
            .I(N__76809));
    LocalMux I__16885 (
            .O(N__76809),
            .I(N__76804));
    InMux I__16884 (
            .O(N__76808),
            .I(N__76801));
    InMux I__16883 (
            .O(N__76807),
            .I(N__76798));
    Span4Mux_h I__16882 (
            .O(N__76804),
            .I(N__76795));
    LocalMux I__16881 (
            .O(N__76801),
            .I(N__76792));
    LocalMux I__16880 (
            .O(N__76798),
            .I(N__76785));
    Span4Mux_v I__16879 (
            .O(N__76795),
            .I(N__76782));
    Span4Mux_h I__16878 (
            .O(N__76792),
            .I(N__76779));
    InMux I__16877 (
            .O(N__76791),
            .I(N__76776));
    InMux I__16876 (
            .O(N__76790),
            .I(N__76773));
    InMux I__16875 (
            .O(N__76789),
            .I(N__76768));
    InMux I__16874 (
            .O(N__76788),
            .I(N__76768));
    Span4Mux_h I__16873 (
            .O(N__76785),
            .I(N__76765));
    Odrv4 I__16872 (
            .O(N__76782),
            .I(control_mode_5));
    Odrv4 I__16871 (
            .O(N__76779),
            .I(control_mode_5));
    LocalMux I__16870 (
            .O(N__76776),
            .I(control_mode_5));
    LocalMux I__16869 (
            .O(N__76773),
            .I(control_mode_5));
    LocalMux I__16868 (
            .O(N__76768),
            .I(control_mode_5));
    Odrv4 I__16867 (
            .O(N__76765),
            .I(control_mode_5));
    CascadeMux I__16866 (
            .O(N__76752),
            .I(N__76747));
    CascadeMux I__16865 (
            .O(N__76751),
            .I(N__76743));
    CascadeMux I__16864 (
            .O(N__76750),
            .I(N__76740));
    InMux I__16863 (
            .O(N__76747),
            .I(N__76735));
    CascadeMux I__16862 (
            .O(N__76746),
            .I(N__76732));
    InMux I__16861 (
            .O(N__76743),
            .I(N__76729));
    InMux I__16860 (
            .O(N__76740),
            .I(N__76726));
    InMux I__16859 (
            .O(N__76739),
            .I(N__76723));
    InMux I__16858 (
            .O(N__76738),
            .I(N__76720));
    LocalMux I__16857 (
            .O(N__76735),
            .I(N__76717));
    InMux I__16856 (
            .O(N__76732),
            .I(N__76714));
    LocalMux I__16855 (
            .O(N__76729),
            .I(N__76710));
    LocalMux I__16854 (
            .O(N__76726),
            .I(N__76707));
    LocalMux I__16853 (
            .O(N__76723),
            .I(N__76702));
    LocalMux I__16852 (
            .O(N__76720),
            .I(N__76702));
    Span4Mux_v I__16851 (
            .O(N__76717),
            .I(N__76697));
    LocalMux I__16850 (
            .O(N__76714),
            .I(N__76697));
    InMux I__16849 (
            .O(N__76713),
            .I(N__76694));
    Span12Mux_h I__16848 (
            .O(N__76710),
            .I(N__76691));
    Span4Mux_h I__16847 (
            .O(N__76707),
            .I(N__76684));
    Span4Mux_h I__16846 (
            .O(N__76702),
            .I(N__76684));
    Span4Mux_h I__16845 (
            .O(N__76697),
            .I(N__76684));
    LocalMux I__16844 (
            .O(N__76694),
            .I(encoder0_position_22));
    Odrv12 I__16843 (
            .O(N__76691),
            .I(encoder0_position_22));
    Odrv4 I__16842 (
            .O(N__76684),
            .I(encoder0_position_22));
    InMux I__16841 (
            .O(N__76677),
            .I(N__76674));
    LocalMux I__16840 (
            .O(N__76674),
            .I(N__76670));
    InMux I__16839 (
            .O(N__76673),
            .I(N__76667));
    Odrv12 I__16838 (
            .O(N__76670),
            .I(\c0.n18199 ));
    LocalMux I__16837 (
            .O(N__76667),
            .I(\c0.n18199 ));
    InMux I__16836 (
            .O(N__76662),
            .I(N__76659));
    LocalMux I__16835 (
            .O(N__76659),
            .I(N__76656));
    Span4Mux_v I__16834 (
            .O(N__76656),
            .I(N__76653));
    Span4Mux_h I__16833 (
            .O(N__76653),
            .I(N__76648));
    InMux I__16832 (
            .O(N__76652),
            .I(N__76645));
    InMux I__16831 (
            .O(N__76651),
            .I(N__76641));
    Span4Mux_h I__16830 (
            .O(N__76648),
            .I(N__76636));
    LocalMux I__16829 (
            .O(N__76645),
            .I(N__76636));
    InMux I__16828 (
            .O(N__76644),
            .I(N__76632));
    LocalMux I__16827 (
            .O(N__76641),
            .I(N__76629));
    Span4Mux_v I__16826 (
            .O(N__76636),
            .I(N__76626));
    InMux I__16825 (
            .O(N__76635),
            .I(N__76623));
    LocalMux I__16824 (
            .O(N__76632),
            .I(encoder1_position_20));
    Odrv4 I__16823 (
            .O(N__76629),
            .I(encoder1_position_20));
    Odrv4 I__16822 (
            .O(N__76626),
            .I(encoder1_position_20));
    LocalMux I__16821 (
            .O(N__76623),
            .I(encoder1_position_20));
    CascadeMux I__16820 (
            .O(N__76614),
            .I(N__76611));
    InMux I__16819 (
            .O(N__76611),
            .I(N__76608));
    LocalMux I__16818 (
            .O(N__76608),
            .I(\c0.data_out_frame_29__7__N_756 ));
    CascadeMux I__16817 (
            .O(N__76605),
            .I(\c0.n18232_cascade_ ));
    InMux I__16816 (
            .O(N__76602),
            .I(N__76599));
    LocalMux I__16815 (
            .O(N__76599),
            .I(N__76596));
    Span4Mux_h I__16814 (
            .O(N__76596),
            .I(N__76593));
    Odrv4 I__16813 (
            .O(N__76593),
            .I(n2273));
    CascadeMux I__16812 (
            .O(N__76590),
            .I(N__76586));
    InMux I__16811 (
            .O(N__76589),
            .I(N__76580));
    InMux I__16810 (
            .O(N__76586),
            .I(N__76576));
    InMux I__16809 (
            .O(N__76585),
            .I(N__76573));
    InMux I__16808 (
            .O(N__76584),
            .I(N__76569));
    CascadeMux I__16807 (
            .O(N__76583),
            .I(N__76566));
    LocalMux I__16806 (
            .O(N__76580),
            .I(N__76558));
    InMux I__16805 (
            .O(N__76579),
            .I(N__76555));
    LocalMux I__16804 (
            .O(N__76576),
            .I(N__76552));
    LocalMux I__16803 (
            .O(N__76573),
            .I(N__76549));
    InMux I__16802 (
            .O(N__76572),
            .I(N__76546));
    LocalMux I__16801 (
            .O(N__76569),
            .I(N__76537));
    InMux I__16800 (
            .O(N__76566),
            .I(N__76532));
    InMux I__16799 (
            .O(N__76565),
            .I(N__76532));
    InMux I__16798 (
            .O(N__76564),
            .I(N__76529));
    InMux I__16797 (
            .O(N__76563),
            .I(N__76524));
    InMux I__16796 (
            .O(N__76562),
            .I(N__76524));
    InMux I__16795 (
            .O(N__76561),
            .I(N__76517));
    Span4Mux_h I__16794 (
            .O(N__76558),
            .I(N__76508));
    LocalMux I__16793 (
            .O(N__76555),
            .I(N__76508));
    Span4Mux_v I__16792 (
            .O(N__76552),
            .I(N__76508));
    Span4Mux_v I__16791 (
            .O(N__76549),
            .I(N__76508));
    LocalMux I__16790 (
            .O(N__76546),
            .I(N__76505));
    InMux I__16789 (
            .O(N__76545),
            .I(N__76500));
    InMux I__16788 (
            .O(N__76544),
            .I(N__76500));
    InMux I__16787 (
            .O(N__76543),
            .I(N__76497));
    InMux I__16786 (
            .O(N__76542),
            .I(N__76490));
    InMux I__16785 (
            .O(N__76541),
            .I(N__76490));
    InMux I__16784 (
            .O(N__76540),
            .I(N__76490));
    Span4Mux_h I__16783 (
            .O(N__76537),
            .I(N__76483));
    LocalMux I__16782 (
            .O(N__76532),
            .I(N__76483));
    LocalMux I__16781 (
            .O(N__76529),
            .I(N__76483));
    LocalMux I__16780 (
            .O(N__76524),
            .I(N__76470));
    InMux I__16779 (
            .O(N__76523),
            .I(N__76467));
    InMux I__16778 (
            .O(N__76522),
            .I(N__76462));
    InMux I__16777 (
            .O(N__76521),
            .I(N__76462));
    InMux I__16776 (
            .O(N__76520),
            .I(N__76459));
    LocalMux I__16775 (
            .O(N__76517),
            .I(N__76452));
    Span4Mux_h I__16774 (
            .O(N__76508),
            .I(N__76452));
    Span4Mux_h I__16773 (
            .O(N__76505),
            .I(N__76452));
    LocalMux I__16772 (
            .O(N__76500),
            .I(N__76447));
    LocalMux I__16771 (
            .O(N__76497),
            .I(N__76447));
    LocalMux I__16770 (
            .O(N__76490),
            .I(N__76442));
    Span4Mux_v I__16769 (
            .O(N__76483),
            .I(N__76442));
    InMux I__16768 (
            .O(N__76482),
            .I(N__76439));
    InMux I__16767 (
            .O(N__76481),
            .I(N__76436));
    InMux I__16766 (
            .O(N__76480),
            .I(N__76433));
    InMux I__16765 (
            .O(N__76479),
            .I(N__76430));
    InMux I__16764 (
            .O(N__76478),
            .I(N__76423));
    InMux I__16763 (
            .O(N__76477),
            .I(N__76423));
    InMux I__16762 (
            .O(N__76476),
            .I(N__76423));
    InMux I__16761 (
            .O(N__76475),
            .I(N__76420));
    InMux I__16760 (
            .O(N__76474),
            .I(N__76415));
    InMux I__16759 (
            .O(N__76473),
            .I(N__76415));
    Span4Mux_h I__16758 (
            .O(N__76470),
            .I(N__76410));
    LocalMux I__16757 (
            .O(N__76467),
            .I(N__76410));
    LocalMux I__16756 (
            .O(N__76462),
            .I(N__76405));
    LocalMux I__16755 (
            .O(N__76459),
            .I(N__76405));
    Span4Mux_v I__16754 (
            .O(N__76452),
            .I(N__76402));
    Span4Mux_h I__16753 (
            .O(N__76447),
            .I(N__76397));
    Span4Mux_v I__16752 (
            .O(N__76442),
            .I(N__76397));
    LocalMux I__16751 (
            .O(N__76439),
            .I(N__76380));
    LocalMux I__16750 (
            .O(N__76436),
            .I(N__76380));
    LocalMux I__16749 (
            .O(N__76433),
            .I(N__76380));
    LocalMux I__16748 (
            .O(N__76430),
            .I(N__76380));
    LocalMux I__16747 (
            .O(N__76423),
            .I(N__76380));
    LocalMux I__16746 (
            .O(N__76420),
            .I(N__76380));
    LocalMux I__16745 (
            .O(N__76415),
            .I(N__76380));
    Sp12to4 I__16744 (
            .O(N__76410),
            .I(N__76380));
    Span4Mux_v I__16743 (
            .O(N__76405),
            .I(N__76375));
    Span4Mux_v I__16742 (
            .O(N__76402),
            .I(N__76375));
    Span4Mux_v I__16741 (
            .O(N__76397),
            .I(N__76372));
    Span12Mux_v I__16740 (
            .O(N__76380),
            .I(N__76369));
    Span4Mux_v I__16739 (
            .O(N__76375),
            .I(N__76366));
    Span4Mux_v I__16738 (
            .O(N__76372),
            .I(N__76363));
    Odrv12 I__16737 (
            .O(N__76369),
            .I(count_enable_adj_4814));
    Odrv4 I__16736 (
            .O(N__76366),
            .I(count_enable_adj_4814));
    Odrv4 I__16735 (
            .O(N__76363),
            .I(count_enable_adj_4814));
    InMux I__16734 (
            .O(N__76356),
            .I(N__76353));
    LocalMux I__16733 (
            .O(N__76353),
            .I(N__76349));
    InMux I__16732 (
            .O(N__76352),
            .I(N__76346));
    Span4Mux_v I__16731 (
            .O(N__76349),
            .I(N__76341));
    LocalMux I__16730 (
            .O(N__76346),
            .I(N__76341));
    Odrv4 I__16729 (
            .O(N__76341),
            .I(\c0.n33902 ));
    CascadeMux I__16728 (
            .O(N__76338),
            .I(\c0.data_out_frame_29__7__N_976_cascade_ ));
    InMux I__16727 (
            .O(N__76335),
            .I(N__76331));
    InMux I__16726 (
            .O(N__76334),
            .I(N__76328));
    LocalMux I__16725 (
            .O(N__76331),
            .I(N__76325));
    LocalMux I__16724 (
            .O(N__76328),
            .I(N__76322));
    Span4Mux_v I__16723 (
            .O(N__76325),
            .I(N__76319));
    Odrv12 I__16722 (
            .O(N__76322),
            .I(\c0.n33772 ));
    Odrv4 I__16721 (
            .O(N__76319),
            .I(\c0.n33772 ));
    InMux I__16720 (
            .O(N__76314),
            .I(N__76311));
    LocalMux I__16719 (
            .O(N__76311),
            .I(\c0.n42_adj_4570 ));
    InMux I__16718 (
            .O(N__76308),
            .I(N__76305));
    LocalMux I__16717 (
            .O(N__76305),
            .I(N__76302));
    Span4Mux_h I__16716 (
            .O(N__76302),
            .I(N__76298));
    InMux I__16715 (
            .O(N__76301),
            .I(N__76295));
    Odrv4 I__16714 (
            .O(N__76298),
            .I(\c0.n33305 ));
    LocalMux I__16713 (
            .O(N__76295),
            .I(\c0.n33305 ));
    InMux I__16712 (
            .O(N__76290),
            .I(N__76287));
    LocalMux I__16711 (
            .O(N__76287),
            .I(\c0.data_out_frame_29__7__N_740 ));
    CascadeMux I__16710 (
            .O(N__76284),
            .I(N__76281));
    InMux I__16709 (
            .O(N__76281),
            .I(N__76278));
    LocalMux I__16708 (
            .O(N__76278),
            .I(N__76275));
    Odrv4 I__16707 (
            .O(N__76275),
            .I(\c0.n18689 ));
    InMux I__16706 (
            .O(N__76272),
            .I(N__76269));
    LocalMux I__16705 (
            .O(N__76269),
            .I(\c0.n6_adj_4560 ));
    InMux I__16704 (
            .O(N__76266),
            .I(N__76263));
    LocalMux I__16703 (
            .O(N__76263),
            .I(N__76258));
    InMux I__16702 (
            .O(N__76262),
            .I(N__76255));
    CascadeMux I__16701 (
            .O(N__76261),
            .I(N__76252));
    Span4Mux_h I__16700 (
            .O(N__76258),
            .I(N__76247));
    LocalMux I__16699 (
            .O(N__76255),
            .I(N__76247));
    InMux I__16698 (
            .O(N__76252),
            .I(N__76244));
    Odrv4 I__16697 (
            .O(N__76247),
            .I(\c0.n18523 ));
    LocalMux I__16696 (
            .O(N__76244),
            .I(\c0.n18523 ));
    CascadeMux I__16695 (
            .O(N__76239),
            .I(\c0.n35113_cascade_ ));
    InMux I__16694 (
            .O(N__76236),
            .I(N__76232));
    InMux I__16693 (
            .O(N__76235),
            .I(N__76229));
    LocalMux I__16692 (
            .O(N__76232),
            .I(\c0.n31401 ));
    LocalMux I__16691 (
            .O(N__76229),
            .I(\c0.n31401 ));
    CascadeMux I__16690 (
            .O(N__76224),
            .I(\c0.n12_adj_4561_cascade_ ));
    InMux I__16689 (
            .O(N__76221),
            .I(N__76218));
    LocalMux I__16688 (
            .O(N__76218),
            .I(N__76215));
    Span4Mux_h I__16687 (
            .O(N__76215),
            .I(N__76211));
    InMux I__16686 (
            .O(N__76214),
            .I(N__76208));
    Span4Mux_v I__16685 (
            .O(N__76211),
            .I(N__76205));
    LocalMux I__16684 (
            .O(N__76208),
            .I(N__76202));
    Odrv4 I__16683 (
            .O(N__76205),
            .I(\c0.n33615 ));
    Odrv4 I__16682 (
            .O(N__76202),
            .I(\c0.n33615 ));
    CascadeMux I__16681 (
            .O(N__76197),
            .I(\c0.n12_adj_4553_cascade_ ));
    InMux I__16680 (
            .O(N__76194),
            .I(N__76191));
    LocalMux I__16679 (
            .O(N__76191),
            .I(N__76187));
    InMux I__16678 (
            .O(N__76190),
            .I(N__76184));
    Span4Mux_h I__16677 (
            .O(N__76187),
            .I(N__76181));
    LocalMux I__16676 (
            .O(N__76184),
            .I(data_out_frame_13_3));
    Odrv4 I__16675 (
            .O(N__76181),
            .I(data_out_frame_13_3));
    InMux I__16674 (
            .O(N__76176),
            .I(N__76172));
    InMux I__16673 (
            .O(N__76175),
            .I(N__76169));
    LocalMux I__16672 (
            .O(N__76172),
            .I(N__76166));
    LocalMux I__16671 (
            .O(N__76169),
            .I(data_out_frame_29_6));
    Odrv4 I__16670 (
            .O(N__76166),
            .I(data_out_frame_29_6));
    InMux I__16669 (
            .O(N__76161),
            .I(N__76158));
    LocalMux I__16668 (
            .O(N__76158),
            .I(N__76155));
    Odrv4 I__16667 (
            .O(N__76155),
            .I(n2267));
    InMux I__16666 (
            .O(N__76152),
            .I(N__76149));
    LocalMux I__16665 (
            .O(N__76149),
            .I(N__76146));
    Span4Mux_h I__16664 (
            .O(N__76146),
            .I(N__76139));
    InMux I__16663 (
            .O(N__76145),
            .I(N__76134));
    InMux I__16662 (
            .O(N__76144),
            .I(N__76134));
    CascadeMux I__16661 (
            .O(N__76143),
            .I(N__76131));
    InMux I__16660 (
            .O(N__76142),
            .I(N__76128));
    Span4Mux_h I__16659 (
            .O(N__76139),
            .I(N__76123));
    LocalMux I__16658 (
            .O(N__76134),
            .I(N__76123));
    InMux I__16657 (
            .O(N__76131),
            .I(N__76119));
    LocalMux I__16656 (
            .O(N__76128),
            .I(N__76116));
    Span4Mux_h I__16655 (
            .O(N__76123),
            .I(N__76113));
    InMux I__16654 (
            .O(N__76122),
            .I(N__76110));
    LocalMux I__16653 (
            .O(N__76119),
            .I(data_in_frame_1_0));
    Odrv12 I__16652 (
            .O(N__76116),
            .I(data_in_frame_1_0));
    Odrv4 I__16651 (
            .O(N__76113),
            .I(data_in_frame_1_0));
    LocalMux I__16650 (
            .O(N__76110),
            .I(data_in_frame_1_0));
    CascadeMux I__16649 (
            .O(N__76101),
            .I(N__76097));
    InMux I__16648 (
            .O(N__76100),
            .I(N__76091));
    InMux I__16647 (
            .O(N__76097),
            .I(N__76091));
    CascadeMux I__16646 (
            .O(N__76096),
            .I(N__76087));
    LocalMux I__16645 (
            .O(N__76091),
            .I(N__76084));
    InMux I__16644 (
            .O(N__76090),
            .I(N__76079));
    InMux I__16643 (
            .O(N__76087),
            .I(N__76076));
    Span4Mux_h I__16642 (
            .O(N__76084),
            .I(N__76073));
    InMux I__16641 (
            .O(N__76083),
            .I(N__76068));
    InMux I__16640 (
            .O(N__76082),
            .I(N__76068));
    LocalMux I__16639 (
            .O(N__76079),
            .I(encoder1_position_13));
    LocalMux I__16638 (
            .O(N__76076),
            .I(encoder1_position_13));
    Odrv4 I__16637 (
            .O(N__76073),
            .I(encoder1_position_13));
    LocalMux I__16636 (
            .O(N__76068),
            .I(encoder1_position_13));
    InMux I__16635 (
            .O(N__76059),
            .I(N__76055));
    InMux I__16634 (
            .O(N__76058),
            .I(N__76051));
    LocalMux I__16633 (
            .O(N__76055),
            .I(N__76047));
    InMux I__16632 (
            .O(N__76054),
            .I(N__76044));
    LocalMux I__16631 (
            .O(N__76051),
            .I(N__76040));
    InMux I__16630 (
            .O(N__76050),
            .I(N__76037));
    Span4Mux_v I__16629 (
            .O(N__76047),
            .I(N__76034));
    LocalMux I__16628 (
            .O(N__76044),
            .I(N__76031));
    InMux I__16627 (
            .O(N__76043),
            .I(N__76028));
    Sp12to4 I__16626 (
            .O(N__76040),
            .I(N__76025));
    LocalMux I__16625 (
            .O(N__76037),
            .I(encoder1_position_12));
    Odrv4 I__16624 (
            .O(N__76034),
            .I(encoder1_position_12));
    Odrv12 I__16623 (
            .O(N__76031),
            .I(encoder1_position_12));
    LocalMux I__16622 (
            .O(N__76028),
            .I(encoder1_position_12));
    Odrv12 I__16621 (
            .O(N__76025),
            .I(encoder1_position_12));
    InMux I__16620 (
            .O(N__76014),
            .I(N__76011));
    LocalMux I__16619 (
            .O(N__76011),
            .I(\quad_counter1.n7_adj_4425 ));
    CascadeMux I__16618 (
            .O(N__76008),
            .I(\quad_counter1.n8_adj_4424_cascade_ ));
    InMux I__16617 (
            .O(N__76005),
            .I(N__76002));
    LocalMux I__16616 (
            .O(N__76002),
            .I(\quad_counter1.n25 ));
    InMux I__16615 (
            .O(N__75999),
            .I(N__75996));
    LocalMux I__16614 (
            .O(N__75996),
            .I(\quad_counter1.n26 ));
    CascadeMux I__16613 (
            .O(N__75993),
            .I(N__75990));
    InMux I__16612 (
            .O(N__75990),
            .I(N__75987));
    LocalMux I__16611 (
            .O(N__75987),
            .I(\quad_counter1.n28 ));
    InMux I__16610 (
            .O(N__75984),
            .I(N__75981));
    LocalMux I__16609 (
            .O(N__75981),
            .I(\quad_counter1.n27 ));
    CascadeMux I__16608 (
            .O(N__75978),
            .I(\quad_counter1.n3332_cascade_ ));
    InMux I__16607 (
            .O(N__75975),
            .I(N__75972));
    LocalMux I__16606 (
            .O(N__75972),
            .I(N__75969));
    Odrv4 I__16605 (
            .O(N__75969),
            .I(n2275));
    InMux I__16604 (
            .O(N__75966),
            .I(N__75963));
    LocalMux I__16603 (
            .O(N__75963),
            .I(N__75960));
    Odrv12 I__16602 (
            .O(N__75960),
            .I(n2277));
    InMux I__16601 (
            .O(N__75957),
            .I(N__75954));
    LocalMux I__16600 (
            .O(N__75954),
            .I(N__75951));
    Odrv12 I__16599 (
            .O(N__75951),
            .I(\c0.n26_adj_4516 ));
    CascadeMux I__16598 (
            .O(N__75948),
            .I(N__75945));
    InMux I__16597 (
            .O(N__75945),
            .I(N__75940));
    CascadeMux I__16596 (
            .O(N__75944),
            .I(N__75937));
    InMux I__16595 (
            .O(N__75943),
            .I(N__75934));
    LocalMux I__16594 (
            .O(N__75940),
            .I(N__75931));
    InMux I__16593 (
            .O(N__75937),
            .I(N__75927));
    LocalMux I__16592 (
            .O(N__75934),
            .I(N__75924));
    Span12Mux_h I__16591 (
            .O(N__75931),
            .I(N__75919));
    InMux I__16590 (
            .O(N__75930),
            .I(N__75916));
    LocalMux I__16589 (
            .O(N__75927),
            .I(N__75913));
    Span4Mux_v I__16588 (
            .O(N__75924),
            .I(N__75910));
    InMux I__16587 (
            .O(N__75923),
            .I(N__75905));
    InMux I__16586 (
            .O(N__75922),
            .I(N__75905));
    Span12Mux_v I__16585 (
            .O(N__75919),
            .I(N__75902));
    LocalMux I__16584 (
            .O(N__75916),
            .I(N__75895));
    Span4Mux_h I__16583 (
            .O(N__75913),
            .I(N__75895));
    Span4Mux_v I__16582 (
            .O(N__75910),
            .I(N__75895));
    LocalMux I__16581 (
            .O(N__75905),
            .I(N__75892));
    Odrv12 I__16580 (
            .O(N__75902),
            .I(encoder0_position_7));
    Odrv4 I__16579 (
            .O(N__75895),
            .I(encoder0_position_7));
    Odrv4 I__16578 (
            .O(N__75892),
            .I(encoder0_position_7));
    CascadeMux I__16577 (
            .O(N__75885),
            .I(N__75882));
    InMux I__16576 (
            .O(N__75882),
            .I(N__75879));
    LocalMux I__16575 (
            .O(N__75879),
            .I(N__75876));
    Span4Mux_h I__16574 (
            .O(N__75876),
            .I(N__75870));
    InMux I__16573 (
            .O(N__75875),
            .I(N__75867));
    CascadeMux I__16572 (
            .O(N__75874),
            .I(N__75864));
    InMux I__16571 (
            .O(N__75873),
            .I(N__75860));
    Span4Mux_h I__16570 (
            .O(N__75870),
            .I(N__75857));
    LocalMux I__16569 (
            .O(N__75867),
            .I(N__75854));
    InMux I__16568 (
            .O(N__75864),
            .I(N__75851));
    InMux I__16567 (
            .O(N__75863),
            .I(N__75848));
    LocalMux I__16566 (
            .O(N__75860),
            .I(encoder1_position_8));
    Odrv4 I__16565 (
            .O(N__75857),
            .I(encoder1_position_8));
    Odrv4 I__16564 (
            .O(N__75854),
            .I(encoder1_position_8));
    LocalMux I__16563 (
            .O(N__75851),
            .I(encoder1_position_8));
    LocalMux I__16562 (
            .O(N__75848),
            .I(encoder1_position_8));
    InMux I__16561 (
            .O(N__75837),
            .I(N__75833));
    InMux I__16560 (
            .O(N__75836),
            .I(N__75830));
    LocalMux I__16559 (
            .O(N__75833),
            .I(N__75827));
    LocalMux I__16558 (
            .O(N__75830),
            .I(N__75819));
    Span4Mux_h I__16557 (
            .O(N__75827),
            .I(N__75819));
    InMux I__16556 (
            .O(N__75826),
            .I(N__75816));
    InMux I__16555 (
            .O(N__75825),
            .I(N__75813));
    InMux I__16554 (
            .O(N__75824),
            .I(N__75810));
    Span4Mux_v I__16553 (
            .O(N__75819),
            .I(N__75807));
    LocalMux I__16552 (
            .O(N__75816),
            .I(N__75804));
    LocalMux I__16551 (
            .O(N__75813),
            .I(encoder0_position_6));
    LocalMux I__16550 (
            .O(N__75810),
            .I(encoder0_position_6));
    Odrv4 I__16549 (
            .O(N__75807),
            .I(encoder0_position_6));
    Odrv4 I__16548 (
            .O(N__75804),
            .I(encoder0_position_6));
    CascadeMux I__16547 (
            .O(N__75795),
            .I(N__75787));
    CascadeMux I__16546 (
            .O(N__75794),
            .I(N__75784));
    CascadeMux I__16545 (
            .O(N__75793),
            .I(N__75781));
    CascadeMux I__16544 (
            .O(N__75792),
            .I(N__75778));
    CascadeMux I__16543 (
            .O(N__75791),
            .I(N__75775));
    CascadeMux I__16542 (
            .O(N__75790),
            .I(N__75772));
    InMux I__16541 (
            .O(N__75787),
            .I(N__75767));
    InMux I__16540 (
            .O(N__75784),
            .I(N__75767));
    InMux I__16539 (
            .O(N__75781),
            .I(N__75758));
    InMux I__16538 (
            .O(N__75778),
            .I(N__75758));
    InMux I__16537 (
            .O(N__75775),
            .I(N__75758));
    InMux I__16536 (
            .O(N__75772),
            .I(N__75758));
    LocalMux I__16535 (
            .O(N__75767),
            .I(\quad_counter1.n36134 ));
    LocalMux I__16534 (
            .O(N__75758),
            .I(\quad_counter1.n36134 ));
    InMux I__16533 (
            .O(N__75753),
            .I(N__75750));
    LocalMux I__16532 (
            .O(N__75750),
            .I(\quad_counter1.n12 ));
    CascadeMux I__16531 (
            .O(N__75747),
            .I(N__75741));
    CascadeMux I__16530 (
            .O(N__75746),
            .I(N__75738));
    CascadeMux I__16529 (
            .O(N__75745),
            .I(N__75732));
    CascadeMux I__16528 (
            .O(N__75744),
            .I(N__75729));
    InMux I__16527 (
            .O(N__75741),
            .I(N__75724));
    InMux I__16526 (
            .O(N__75738),
            .I(N__75724));
    CascadeMux I__16525 (
            .O(N__75737),
            .I(N__75721));
    CascadeMux I__16524 (
            .O(N__75736),
            .I(N__75718));
    CascadeMux I__16523 (
            .O(N__75735),
            .I(N__75715));
    InMux I__16522 (
            .O(N__75732),
            .I(N__75709));
    InMux I__16521 (
            .O(N__75729),
            .I(N__75709));
    LocalMux I__16520 (
            .O(N__75724),
            .I(N__75706));
    InMux I__16519 (
            .O(N__75721),
            .I(N__75697));
    InMux I__16518 (
            .O(N__75718),
            .I(N__75697));
    InMux I__16517 (
            .O(N__75715),
            .I(N__75697));
    InMux I__16516 (
            .O(N__75714),
            .I(N__75697));
    LocalMux I__16515 (
            .O(N__75709),
            .I(\quad_counter1.n2441 ));
    Odrv4 I__16514 (
            .O(N__75706),
            .I(\quad_counter1.n2441 ));
    LocalMux I__16513 (
            .O(N__75697),
            .I(\quad_counter1.n2441 ));
    InMux I__16512 (
            .O(N__75690),
            .I(N__75687));
    LocalMux I__16511 (
            .O(N__75687),
            .I(n34871));
    InMux I__16510 (
            .O(N__75684),
            .I(N__75678));
    InMux I__16509 (
            .O(N__75683),
            .I(N__75678));
    LocalMux I__16508 (
            .O(N__75678),
            .I(count_prev_0_adj_4815));
    CascadeMux I__16507 (
            .O(N__75675),
            .I(n34871_cascade_));
    CascadeMux I__16506 (
            .O(N__75672),
            .I(\quad_counter1.n18_cascade_ ));
    InMux I__16505 (
            .O(N__75669),
            .I(\quad_counter1.n30513 ));
    InMux I__16504 (
            .O(N__75666),
            .I(\quad_counter1.n30514 ));
    InMux I__16503 (
            .O(N__75663),
            .I(\quad_counter1.n30515 ));
    InMux I__16502 (
            .O(N__75660),
            .I(\quad_counter1.n30516 ));
    InMux I__16501 (
            .O(N__75657),
            .I(bfn_21_10_0_));
    InMux I__16500 (
            .O(N__75654),
            .I(\quad_counter1.n30518 ));
    InMux I__16499 (
            .O(N__75651),
            .I(\quad_counter1.n30519 ));
    InMux I__16498 (
            .O(N__75648),
            .I(\quad_counter1.n30520 ));
    InMux I__16497 (
            .O(N__75645),
            .I(\quad_counter1.n30521 ));
    CascadeMux I__16496 (
            .O(N__75642),
            .I(\quad_counter1.n14_cascade_ ));
    CascadeMux I__16495 (
            .O(N__75639),
            .I(\quad_counter1.n28273_cascade_ ));
    CascadeMux I__16494 (
            .O(N__75636),
            .I(\quad_counter1.n10_adj_4450_cascade_ ));
    InMux I__16493 (
            .O(N__75633),
            .I(N__75630));
    LocalMux I__16492 (
            .O(N__75630),
            .I(\quad_counter1.n9_adj_4451 ));
    InMux I__16491 (
            .O(N__75627),
            .I(bfn_21_9_0_));
    InMux I__16490 (
            .O(N__75624),
            .I(\quad_counter1.n30510 ));
    InMux I__16489 (
            .O(N__75621),
            .I(\quad_counter1.n30511 ));
    InMux I__16488 (
            .O(N__75618),
            .I(\quad_counter1.n30512 ));
    InMux I__16487 (
            .O(N__75615),
            .I(N__75610));
    InMux I__16486 (
            .O(N__75614),
            .I(N__75607));
    InMux I__16485 (
            .O(N__75613),
            .I(N__75604));
    LocalMux I__16484 (
            .O(N__75610),
            .I(\quad_counter1.n2712 ));
    LocalMux I__16483 (
            .O(N__75607),
            .I(\quad_counter1.n2712 ));
    LocalMux I__16482 (
            .O(N__75604),
            .I(\quad_counter1.n2712 ));
    InMux I__16481 (
            .O(N__75597),
            .I(\quad_counter1.n30541 ));
    InMux I__16480 (
            .O(N__75594),
            .I(bfn_21_6_0_));
    InMux I__16479 (
            .O(N__75591),
            .I(\quad_counter1.n30543 ));
    InMux I__16478 (
            .O(N__75588),
            .I(\quad_counter1.n30544 ));
    InMux I__16477 (
            .O(N__75585),
            .I(\quad_counter1.n30545 ));
    InMux I__16476 (
            .O(N__75582),
            .I(\quad_counter1.n30546 ));
    InMux I__16475 (
            .O(N__75579),
            .I(\quad_counter1.n30547 ));
    InMux I__16474 (
            .O(N__75576),
            .I(\quad_counter1.n30548 ));
    CascadeMux I__16473 (
            .O(N__75573),
            .I(\quad_counter1.n10_adj_4468_cascade_ ));
    CascadeMux I__16472 (
            .O(N__75570),
            .I(N__75562));
    CascadeMux I__16471 (
            .O(N__75569),
            .I(N__75559));
    CascadeMux I__16470 (
            .O(N__75568),
            .I(N__75556));
    CascadeMux I__16469 (
            .O(N__75567),
            .I(N__75553));
    CascadeMux I__16468 (
            .O(N__75566),
            .I(N__75550));
    CascadeMux I__16467 (
            .O(N__75565),
            .I(N__75547));
    InMux I__16466 (
            .O(N__75562),
            .I(N__75542));
    InMux I__16465 (
            .O(N__75559),
            .I(N__75542));
    InMux I__16464 (
            .O(N__75556),
            .I(N__75533));
    InMux I__16463 (
            .O(N__75553),
            .I(N__75533));
    InMux I__16462 (
            .O(N__75550),
            .I(N__75533));
    InMux I__16461 (
            .O(N__75547),
            .I(N__75533));
    LocalMux I__16460 (
            .O(N__75542),
            .I(\quad_counter1.n36130 ));
    LocalMux I__16459 (
            .O(N__75533),
            .I(\quad_counter1.n36130 ));
    CascadeMux I__16458 (
            .O(N__75528),
            .I(N__75523));
    InMux I__16457 (
            .O(N__75527),
            .I(N__75520));
    InMux I__16456 (
            .O(N__75526),
            .I(N__75517));
    InMux I__16455 (
            .O(N__75523),
            .I(N__75514));
    LocalMux I__16454 (
            .O(N__75520),
            .I(\quad_counter1.n2719 ));
    LocalMux I__16453 (
            .O(N__75517),
            .I(\quad_counter1.n2719 ));
    LocalMux I__16452 (
            .O(N__75514),
            .I(\quad_counter1.n2719 ));
    InMux I__16451 (
            .O(N__75507),
            .I(bfn_21_5_0_));
    InMux I__16450 (
            .O(N__75504),
            .I(N__75500));
    InMux I__16449 (
            .O(N__75503),
            .I(N__75496));
    LocalMux I__16448 (
            .O(N__75500),
            .I(N__75493));
    InMux I__16447 (
            .O(N__75499),
            .I(N__75490));
    LocalMux I__16446 (
            .O(N__75496),
            .I(\quad_counter1.n2718 ));
    Odrv4 I__16445 (
            .O(N__75493),
            .I(\quad_counter1.n2718 ));
    LocalMux I__16444 (
            .O(N__75490),
            .I(\quad_counter1.n2718 ));
    InMux I__16443 (
            .O(N__75483),
            .I(\quad_counter1.n30535 ));
    InMux I__16442 (
            .O(N__75480),
            .I(N__75475));
    InMux I__16441 (
            .O(N__75479),
            .I(N__75472));
    InMux I__16440 (
            .O(N__75478),
            .I(N__75469));
    LocalMux I__16439 (
            .O(N__75475),
            .I(\quad_counter1.n2717 ));
    LocalMux I__16438 (
            .O(N__75472),
            .I(\quad_counter1.n2717 ));
    LocalMux I__16437 (
            .O(N__75469),
            .I(\quad_counter1.n2717 ));
    InMux I__16436 (
            .O(N__75462),
            .I(\quad_counter1.n30536 ));
    InMux I__16435 (
            .O(N__75459),
            .I(N__75454));
    InMux I__16434 (
            .O(N__75458),
            .I(N__75451));
    InMux I__16433 (
            .O(N__75457),
            .I(N__75448));
    LocalMux I__16432 (
            .O(N__75454),
            .I(\quad_counter1.n2716 ));
    LocalMux I__16431 (
            .O(N__75451),
            .I(\quad_counter1.n2716 ));
    LocalMux I__16430 (
            .O(N__75448),
            .I(\quad_counter1.n2716 ));
    InMux I__16429 (
            .O(N__75441),
            .I(\quad_counter1.n30537 ));
    InMux I__16428 (
            .O(N__75438),
            .I(N__75433));
    InMux I__16427 (
            .O(N__75437),
            .I(N__75430));
    InMux I__16426 (
            .O(N__75436),
            .I(N__75427));
    LocalMux I__16425 (
            .O(N__75433),
            .I(\quad_counter1.n2715 ));
    LocalMux I__16424 (
            .O(N__75430),
            .I(\quad_counter1.n2715 ));
    LocalMux I__16423 (
            .O(N__75427),
            .I(\quad_counter1.n2715 ));
    InMux I__16422 (
            .O(N__75420),
            .I(\quad_counter1.n30538 ));
    InMux I__16421 (
            .O(N__75417),
            .I(N__75412));
    InMux I__16420 (
            .O(N__75416),
            .I(N__75409));
    InMux I__16419 (
            .O(N__75415),
            .I(N__75406));
    LocalMux I__16418 (
            .O(N__75412),
            .I(\quad_counter1.n2714 ));
    LocalMux I__16417 (
            .O(N__75409),
            .I(\quad_counter1.n2714 ));
    LocalMux I__16416 (
            .O(N__75406),
            .I(\quad_counter1.n2714 ));
    InMux I__16415 (
            .O(N__75399),
            .I(\quad_counter1.n30539 ));
    InMux I__16414 (
            .O(N__75396),
            .I(\quad_counter1.n30540 ));
    CascadeMux I__16413 (
            .O(N__75393),
            .I(N__75388));
    InMux I__16412 (
            .O(N__75392),
            .I(N__75385));
    InMux I__16411 (
            .O(N__75391),
            .I(N__75380));
    InMux I__16410 (
            .O(N__75388),
            .I(N__75380));
    LocalMux I__16409 (
            .O(N__75385),
            .I(N__75377));
    LocalMux I__16408 (
            .O(N__75380),
            .I(\c0.data_in_frame_24_7 ));
    Odrv12 I__16407 (
            .O(N__75377),
            .I(\c0.data_in_frame_24_7 ));
    InMux I__16406 (
            .O(N__75372),
            .I(N__75366));
    InMux I__16405 (
            .O(N__75371),
            .I(N__75355));
    InMux I__16404 (
            .O(N__75370),
            .I(N__75352));
    InMux I__16403 (
            .O(N__75369),
            .I(N__75348));
    LocalMux I__16402 (
            .O(N__75366),
            .I(N__75345));
    InMux I__16401 (
            .O(N__75365),
            .I(N__75340));
    InMux I__16400 (
            .O(N__75364),
            .I(N__75336));
    InMux I__16399 (
            .O(N__75363),
            .I(N__75330));
    InMux I__16398 (
            .O(N__75362),
            .I(N__75330));
    InMux I__16397 (
            .O(N__75361),
            .I(N__75327));
    InMux I__16396 (
            .O(N__75360),
            .I(N__75321));
    InMux I__16395 (
            .O(N__75359),
            .I(N__75311));
    InMux I__16394 (
            .O(N__75358),
            .I(N__75311));
    LocalMux I__16393 (
            .O(N__75355),
            .I(N__75306));
    LocalMux I__16392 (
            .O(N__75352),
            .I(N__75306));
    InMux I__16391 (
            .O(N__75351),
            .I(N__75303));
    LocalMux I__16390 (
            .O(N__75348),
            .I(N__75300));
    Span4Mux_h I__16389 (
            .O(N__75345),
            .I(N__75297));
    CascadeMux I__16388 (
            .O(N__75344),
            .I(N__75293));
    InMux I__16387 (
            .O(N__75343),
            .I(N__75290));
    LocalMux I__16386 (
            .O(N__75340),
            .I(N__75286));
    InMux I__16385 (
            .O(N__75339),
            .I(N__75283));
    LocalMux I__16384 (
            .O(N__75336),
            .I(N__75280));
    InMux I__16383 (
            .O(N__75335),
            .I(N__75277));
    LocalMux I__16382 (
            .O(N__75330),
            .I(N__75274));
    LocalMux I__16381 (
            .O(N__75327),
            .I(N__75271));
    InMux I__16380 (
            .O(N__75326),
            .I(N__75266));
    InMux I__16379 (
            .O(N__75325),
            .I(N__75263));
    InMux I__16378 (
            .O(N__75324),
            .I(N__75260));
    LocalMux I__16377 (
            .O(N__75321),
            .I(N__75257));
    InMux I__16376 (
            .O(N__75320),
            .I(N__75254));
    InMux I__16375 (
            .O(N__75319),
            .I(N__75249));
    InMux I__16374 (
            .O(N__75318),
            .I(N__75249));
    InMux I__16373 (
            .O(N__75317),
            .I(N__75244));
    InMux I__16372 (
            .O(N__75316),
            .I(N__75244));
    LocalMux I__16371 (
            .O(N__75311),
            .I(N__75241));
    Span4Mux_h I__16370 (
            .O(N__75306),
            .I(N__75238));
    LocalMux I__16369 (
            .O(N__75303),
            .I(N__75231));
    Span4Mux_h I__16368 (
            .O(N__75300),
            .I(N__75231));
    Span4Mux_v I__16367 (
            .O(N__75297),
            .I(N__75231));
    InMux I__16366 (
            .O(N__75296),
            .I(N__75224));
    InMux I__16365 (
            .O(N__75293),
            .I(N__75224));
    LocalMux I__16364 (
            .O(N__75290),
            .I(N__75221));
    InMux I__16363 (
            .O(N__75289),
            .I(N__75218));
    Span4Mux_v I__16362 (
            .O(N__75286),
            .I(N__75213));
    LocalMux I__16361 (
            .O(N__75283),
            .I(N__75213));
    Span4Mux_h I__16360 (
            .O(N__75280),
            .I(N__75210));
    LocalMux I__16359 (
            .O(N__75277),
            .I(N__75203));
    Span4Mux_h I__16358 (
            .O(N__75274),
            .I(N__75203));
    Span4Mux_v I__16357 (
            .O(N__75271),
            .I(N__75203));
    InMux I__16356 (
            .O(N__75270),
            .I(N__75197));
    InMux I__16355 (
            .O(N__75269),
            .I(N__75197));
    LocalMux I__16354 (
            .O(N__75266),
            .I(N__75194));
    LocalMux I__16353 (
            .O(N__75263),
            .I(N__75191));
    LocalMux I__16352 (
            .O(N__75260),
            .I(N__75186));
    Span4Mux_h I__16351 (
            .O(N__75257),
            .I(N__75186));
    LocalMux I__16350 (
            .O(N__75254),
            .I(N__75173));
    LocalMux I__16349 (
            .O(N__75249),
            .I(N__75173));
    LocalMux I__16348 (
            .O(N__75244),
            .I(N__75173));
    Span4Mux_v I__16347 (
            .O(N__75241),
            .I(N__75173));
    Span4Mux_h I__16346 (
            .O(N__75238),
            .I(N__75173));
    Span4Mux_h I__16345 (
            .O(N__75231),
            .I(N__75173));
    InMux I__16344 (
            .O(N__75230),
            .I(N__75170));
    InMux I__16343 (
            .O(N__75229),
            .I(N__75167));
    LocalMux I__16342 (
            .O(N__75224),
            .I(N__75164));
    Span4Mux_h I__16341 (
            .O(N__75221),
            .I(N__75161));
    LocalMux I__16340 (
            .O(N__75218),
            .I(N__75156));
    Span4Mux_h I__16339 (
            .O(N__75213),
            .I(N__75156));
    Span4Mux_h I__16338 (
            .O(N__75210),
            .I(N__75151));
    Span4Mux_h I__16337 (
            .O(N__75203),
            .I(N__75151));
    InMux I__16336 (
            .O(N__75202),
            .I(N__75148));
    LocalMux I__16335 (
            .O(N__75197),
            .I(N__75145));
    Span4Mux_h I__16334 (
            .O(N__75194),
            .I(N__75136));
    Span4Mux_v I__16333 (
            .O(N__75191),
            .I(N__75136));
    Span4Mux_h I__16332 (
            .O(N__75186),
            .I(N__75136));
    Span4Mux_v I__16331 (
            .O(N__75173),
            .I(N__75136));
    LocalMux I__16330 (
            .O(N__75170),
            .I(N__75125));
    LocalMux I__16329 (
            .O(N__75167),
            .I(N__75125));
    Span4Mux_h I__16328 (
            .O(N__75164),
            .I(N__75125));
    Span4Mux_h I__16327 (
            .O(N__75161),
            .I(N__75125));
    Span4Mux_v I__16326 (
            .O(N__75156),
            .I(N__75125));
    Span4Mux_v I__16325 (
            .O(N__75151),
            .I(N__75122));
    LocalMux I__16324 (
            .O(N__75148),
            .I(rx_data_1));
    Odrv4 I__16323 (
            .O(N__75145),
            .I(rx_data_1));
    Odrv4 I__16322 (
            .O(N__75136),
            .I(rx_data_1));
    Odrv4 I__16321 (
            .O(N__75125),
            .I(rx_data_1));
    Odrv4 I__16320 (
            .O(N__75122),
            .I(rx_data_1));
    CascadeMux I__16319 (
            .O(N__75111),
            .I(N__75107));
    InMux I__16318 (
            .O(N__75110),
            .I(N__75103));
    InMux I__16317 (
            .O(N__75107),
            .I(N__75098));
    InMux I__16316 (
            .O(N__75106),
            .I(N__75098));
    LocalMux I__16315 (
            .O(N__75103),
            .I(\c0.data_in_frame_25_1 ));
    LocalMux I__16314 (
            .O(N__75098),
            .I(\c0.data_in_frame_25_1 ));
    InMux I__16313 (
            .O(N__75093),
            .I(N__75090));
    LocalMux I__16312 (
            .O(N__75090),
            .I(N__75080));
    InMux I__16311 (
            .O(N__75089),
            .I(N__75076));
    InMux I__16310 (
            .O(N__75088),
            .I(N__75073));
    InMux I__16309 (
            .O(N__75087),
            .I(N__75067));
    InMux I__16308 (
            .O(N__75086),
            .I(N__75067));
    InMux I__16307 (
            .O(N__75085),
            .I(N__75063));
    InMux I__16306 (
            .O(N__75084),
            .I(N__75058));
    InMux I__16305 (
            .O(N__75083),
            .I(N__75055));
    Span4Mux_v I__16304 (
            .O(N__75080),
            .I(N__75045));
    InMux I__16303 (
            .O(N__75079),
            .I(N__75042));
    LocalMux I__16302 (
            .O(N__75076),
            .I(N__75039));
    LocalMux I__16301 (
            .O(N__75073),
            .I(N__75036));
    InMux I__16300 (
            .O(N__75072),
            .I(N__75033));
    LocalMux I__16299 (
            .O(N__75067),
            .I(N__75030));
    InMux I__16298 (
            .O(N__75066),
            .I(N__75027));
    LocalMux I__16297 (
            .O(N__75063),
            .I(N__75024));
    InMux I__16296 (
            .O(N__75062),
            .I(N__75021));
    InMux I__16295 (
            .O(N__75061),
            .I(N__75018));
    LocalMux I__16294 (
            .O(N__75058),
            .I(N__75015));
    LocalMux I__16293 (
            .O(N__75055),
            .I(N__75012));
    InMux I__16292 (
            .O(N__75054),
            .I(N__75005));
    InMux I__16291 (
            .O(N__75053),
            .I(N__75002));
    InMux I__16290 (
            .O(N__75052),
            .I(N__74999));
    InMux I__16289 (
            .O(N__75051),
            .I(N__74996));
    InMux I__16288 (
            .O(N__75050),
            .I(N__74993));
    InMux I__16287 (
            .O(N__75049),
            .I(N__74987));
    InMux I__16286 (
            .O(N__75048),
            .I(N__74987));
    Span4Mux_v I__16285 (
            .O(N__75045),
            .I(N__74982));
    LocalMux I__16284 (
            .O(N__75042),
            .I(N__74982));
    Span4Mux_v I__16283 (
            .O(N__75039),
            .I(N__74975));
    Span4Mux_v I__16282 (
            .O(N__75036),
            .I(N__74975));
    LocalMux I__16281 (
            .O(N__75033),
            .I(N__74975));
    Span4Mux_v I__16280 (
            .O(N__75030),
            .I(N__74972));
    LocalMux I__16279 (
            .O(N__75027),
            .I(N__74965));
    Span4Mux_h I__16278 (
            .O(N__75024),
            .I(N__74965));
    LocalMux I__16277 (
            .O(N__75021),
            .I(N__74965));
    LocalMux I__16276 (
            .O(N__75018),
            .I(N__74962));
    Span4Mux_h I__16275 (
            .O(N__75015),
            .I(N__74959));
    Span4Mux_v I__16274 (
            .O(N__75012),
            .I(N__74956));
    InMux I__16273 (
            .O(N__75011),
            .I(N__74953));
    InMux I__16272 (
            .O(N__75010),
            .I(N__74950));
    InMux I__16271 (
            .O(N__75009),
            .I(N__74943));
    InMux I__16270 (
            .O(N__75008),
            .I(N__74940));
    LocalMux I__16269 (
            .O(N__75005),
            .I(N__74937));
    LocalMux I__16268 (
            .O(N__75002),
            .I(N__74934));
    LocalMux I__16267 (
            .O(N__74999),
            .I(N__74931));
    LocalMux I__16266 (
            .O(N__74996),
            .I(N__74928));
    LocalMux I__16265 (
            .O(N__74993),
            .I(N__74925));
    InMux I__16264 (
            .O(N__74992),
            .I(N__74922));
    LocalMux I__16263 (
            .O(N__74987),
            .I(N__74917));
    Span4Mux_v I__16262 (
            .O(N__74982),
            .I(N__74917));
    Span4Mux_v I__16261 (
            .O(N__74975),
            .I(N__74912));
    Span4Mux_h I__16260 (
            .O(N__74972),
            .I(N__74912));
    Sp12to4 I__16259 (
            .O(N__74965),
            .I(N__74909));
    Sp12to4 I__16258 (
            .O(N__74962),
            .I(N__74904));
    Sp12to4 I__16257 (
            .O(N__74959),
            .I(N__74904));
    Span4Mux_h I__16256 (
            .O(N__74956),
            .I(N__74901));
    LocalMux I__16255 (
            .O(N__74953),
            .I(N__74896));
    LocalMux I__16254 (
            .O(N__74950),
            .I(N__74896));
    InMux I__16253 (
            .O(N__74949),
            .I(N__74890));
    InMux I__16252 (
            .O(N__74948),
            .I(N__74887));
    InMux I__16251 (
            .O(N__74947),
            .I(N__74882));
    InMux I__16250 (
            .O(N__74946),
            .I(N__74882));
    LocalMux I__16249 (
            .O(N__74943),
            .I(N__74877));
    LocalMux I__16248 (
            .O(N__74940),
            .I(N__74877));
    Span4Mux_v I__16247 (
            .O(N__74937),
            .I(N__74874));
    Span4Mux_v I__16246 (
            .O(N__74934),
            .I(N__74871));
    Span4Mux_v I__16245 (
            .O(N__74931),
            .I(N__74864));
    Span4Mux_v I__16244 (
            .O(N__74928),
            .I(N__74864));
    Span4Mux_v I__16243 (
            .O(N__74925),
            .I(N__74864));
    LocalMux I__16242 (
            .O(N__74922),
            .I(N__74855));
    Sp12to4 I__16241 (
            .O(N__74917),
            .I(N__74855));
    Sp12to4 I__16240 (
            .O(N__74912),
            .I(N__74855));
    Span12Mux_s5_v I__16239 (
            .O(N__74909),
            .I(N__74855));
    Span12Mux_v I__16238 (
            .O(N__74904),
            .I(N__74848));
    Sp12to4 I__16237 (
            .O(N__74901),
            .I(N__74848));
    Span12Mux_s11_v I__16236 (
            .O(N__74896),
            .I(N__74848));
    InMux I__16235 (
            .O(N__74895),
            .I(N__74843));
    InMux I__16234 (
            .O(N__74894),
            .I(N__74843));
    InMux I__16233 (
            .O(N__74893),
            .I(N__74840));
    LocalMux I__16232 (
            .O(N__74890),
            .I(N__74825));
    LocalMux I__16231 (
            .O(N__74887),
            .I(N__74825));
    LocalMux I__16230 (
            .O(N__74882),
            .I(N__74825));
    Span12Mux_s11_v I__16229 (
            .O(N__74877),
            .I(N__74825));
    Sp12to4 I__16228 (
            .O(N__74874),
            .I(N__74825));
    Sp12to4 I__16227 (
            .O(N__74871),
            .I(N__74825));
    Sp12to4 I__16226 (
            .O(N__74864),
            .I(N__74825));
    Span12Mux_h I__16225 (
            .O(N__74855),
            .I(N__74822));
    Span12Mux_h I__16224 (
            .O(N__74848),
            .I(N__74819));
    LocalMux I__16223 (
            .O(N__74843),
            .I(rx_data_5));
    LocalMux I__16222 (
            .O(N__74840),
            .I(rx_data_5));
    Odrv12 I__16221 (
            .O(N__74825),
            .I(rx_data_5));
    Odrv12 I__16220 (
            .O(N__74822),
            .I(rx_data_5));
    Odrv12 I__16219 (
            .O(N__74819),
            .I(rx_data_5));
    InMux I__16218 (
            .O(N__74808),
            .I(N__74803));
    InMux I__16217 (
            .O(N__74807),
            .I(N__74800));
    CascadeMux I__16216 (
            .O(N__74806),
            .I(N__74797));
    LocalMux I__16215 (
            .O(N__74803),
            .I(N__74794));
    LocalMux I__16214 (
            .O(N__74800),
            .I(N__74791));
    InMux I__16213 (
            .O(N__74797),
            .I(N__74787));
    Span4Mux_v I__16212 (
            .O(N__74794),
            .I(N__74782));
    Span4Mux_h I__16211 (
            .O(N__74791),
            .I(N__74782));
    InMux I__16210 (
            .O(N__74790),
            .I(N__74779));
    LocalMux I__16209 (
            .O(N__74787),
            .I(N__74776));
    Span4Mux_h I__16208 (
            .O(N__74782),
            .I(N__74771));
    LocalMux I__16207 (
            .O(N__74779),
            .I(N__74771));
    Span4Mux_h I__16206 (
            .O(N__74776),
            .I(N__74768));
    Span4Mux_v I__16205 (
            .O(N__74771),
            .I(N__74765));
    Odrv4 I__16204 (
            .O(N__74768),
            .I(\c0.n35211 ));
    Odrv4 I__16203 (
            .O(N__74765),
            .I(\c0.n35211 ));
    InMux I__16202 (
            .O(N__74760),
            .I(N__74756));
    CascadeMux I__16201 (
            .O(N__74759),
            .I(N__74753));
    LocalMux I__16200 (
            .O(N__74756),
            .I(N__74749));
    InMux I__16199 (
            .O(N__74753),
            .I(N__74744));
    InMux I__16198 (
            .O(N__74752),
            .I(N__74744));
    Span4Mux_h I__16197 (
            .O(N__74749),
            .I(N__74741));
    LocalMux I__16196 (
            .O(N__74744),
            .I(\c0.data_in_frame_24_5 ));
    Odrv4 I__16195 (
            .O(N__74741),
            .I(\c0.data_in_frame_24_5 ));
    InMux I__16194 (
            .O(N__74736),
            .I(N__74733));
    LocalMux I__16193 (
            .O(N__74733),
            .I(\c0.n33988 ));
    CascadeMux I__16192 (
            .O(N__74730),
            .I(\c0.n33930_cascade_ ));
    InMux I__16191 (
            .O(N__74727),
            .I(N__74722));
    InMux I__16190 (
            .O(N__74726),
            .I(N__74719));
    InMux I__16189 (
            .O(N__74725),
            .I(N__74716));
    LocalMux I__16188 (
            .O(N__74722),
            .I(N__74709));
    LocalMux I__16187 (
            .O(N__74719),
            .I(N__74709));
    LocalMux I__16186 (
            .O(N__74716),
            .I(N__74706));
    InMux I__16185 (
            .O(N__74715),
            .I(N__74703));
    CascadeMux I__16184 (
            .O(N__74714),
            .I(N__74700));
    Span4Mux_v I__16183 (
            .O(N__74709),
            .I(N__74693));
    Span4Mux_v I__16182 (
            .O(N__74706),
            .I(N__74693));
    LocalMux I__16181 (
            .O(N__74703),
            .I(N__74693));
    InMux I__16180 (
            .O(N__74700),
            .I(N__74690));
    Span4Mux_h I__16179 (
            .O(N__74693),
            .I(N__74687));
    LocalMux I__16178 (
            .O(N__74690),
            .I(N__74684));
    Span4Mux_h I__16177 (
            .O(N__74687),
            .I(N__74681));
    Span4Mux_h I__16176 (
            .O(N__74684),
            .I(N__74678));
    Odrv4 I__16175 (
            .O(N__74681),
            .I(\c0.n32341 ));
    Odrv4 I__16174 (
            .O(N__74678),
            .I(\c0.n32341 ));
    InMux I__16173 (
            .O(N__74673),
            .I(N__74670));
    LocalMux I__16172 (
            .O(N__74670),
            .I(\c0.n10_adj_4674 ));
    InMux I__16171 (
            .O(N__74667),
            .I(N__74663));
    InMux I__16170 (
            .O(N__74666),
            .I(N__74660));
    LocalMux I__16169 (
            .O(N__74663),
            .I(N__74654));
    LocalMux I__16168 (
            .O(N__74660),
            .I(N__74654));
    InMux I__16167 (
            .O(N__74659),
            .I(N__74651));
    Odrv4 I__16166 (
            .O(N__74654),
            .I(\quad_counter1.n2811 ));
    LocalMux I__16165 (
            .O(N__74651),
            .I(\quad_counter1.n2811 ));
    InMux I__16164 (
            .O(N__74646),
            .I(N__74642));
    InMux I__16163 (
            .O(N__74645),
            .I(N__74639));
    LocalMux I__16162 (
            .O(N__74642),
            .I(N__74633));
    LocalMux I__16161 (
            .O(N__74639),
            .I(N__74633));
    InMux I__16160 (
            .O(N__74638),
            .I(N__74630));
    Odrv4 I__16159 (
            .O(N__74633),
            .I(\quad_counter1.n2807 ));
    LocalMux I__16158 (
            .O(N__74630),
            .I(\quad_counter1.n2807 ));
    InMux I__16157 (
            .O(N__74625),
            .I(N__74620));
    InMux I__16156 (
            .O(N__74624),
            .I(N__74617));
    CascadeMux I__16155 (
            .O(N__74623),
            .I(N__74614));
    LocalMux I__16154 (
            .O(N__74620),
            .I(N__74609));
    LocalMux I__16153 (
            .O(N__74617),
            .I(N__74609));
    InMux I__16152 (
            .O(N__74614),
            .I(N__74606));
    Odrv4 I__16151 (
            .O(N__74609),
            .I(\quad_counter1.n2810 ));
    LocalMux I__16150 (
            .O(N__74606),
            .I(\quad_counter1.n2810 ));
    InMux I__16149 (
            .O(N__74601),
            .I(N__74598));
    LocalMux I__16148 (
            .O(N__74598),
            .I(N__74594));
    InMux I__16147 (
            .O(N__74597),
            .I(N__74591));
    Span4Mux_h I__16146 (
            .O(N__74594),
            .I(N__74587));
    LocalMux I__16145 (
            .O(N__74591),
            .I(N__74584));
    InMux I__16144 (
            .O(N__74590),
            .I(N__74581));
    Odrv4 I__16143 (
            .O(N__74587),
            .I(\quad_counter1.n2813 ));
    Odrv4 I__16142 (
            .O(N__74584),
            .I(\quad_counter1.n2813 ));
    LocalMux I__16141 (
            .O(N__74581),
            .I(\quad_counter1.n2813 ));
    InMux I__16140 (
            .O(N__74574),
            .I(N__74571));
    LocalMux I__16139 (
            .O(N__74571),
            .I(\quad_counter1.n18_adj_4457 ));
    CascadeMux I__16138 (
            .O(N__74568),
            .I(\quad_counter1.n28269_cascade_ ));
    InMux I__16137 (
            .O(N__74565),
            .I(N__74561));
    InMux I__16136 (
            .O(N__74564),
            .I(N__74558));
    LocalMux I__16135 (
            .O(N__74561),
            .I(N__74555));
    LocalMux I__16134 (
            .O(N__74558),
            .I(\c0.n33948 ));
    Odrv4 I__16133 (
            .O(N__74555),
            .I(\c0.n33948 ));
    InMux I__16132 (
            .O(N__74550),
            .I(N__74544));
    InMux I__16131 (
            .O(N__74549),
            .I(N__74544));
    LocalMux I__16130 (
            .O(N__74544),
            .I(N__74540));
    InMux I__16129 (
            .O(N__74543),
            .I(N__74537));
    Span4Mux_h I__16128 (
            .O(N__74540),
            .I(N__74534));
    LocalMux I__16127 (
            .O(N__74537),
            .I(N__74531));
    Span4Mux_h I__16126 (
            .O(N__74534),
            .I(N__74528));
    Odrv12 I__16125 (
            .O(N__74531),
            .I(\c0.n33467 ));
    Odrv4 I__16124 (
            .O(N__74528),
            .I(\c0.n33467 ));
    CascadeMux I__16123 (
            .O(N__74523),
            .I(N__74519));
    InMux I__16122 (
            .O(N__74522),
            .I(N__74516));
    InMux I__16121 (
            .O(N__74519),
            .I(N__74512));
    LocalMux I__16120 (
            .O(N__74516),
            .I(N__74509));
    InMux I__16119 (
            .O(N__74515),
            .I(N__74506));
    LocalMux I__16118 (
            .O(N__74512),
            .I(\c0.data_in_frame_27_3 ));
    Odrv12 I__16117 (
            .O(N__74509),
            .I(\c0.data_in_frame_27_3 ));
    LocalMux I__16116 (
            .O(N__74506),
            .I(\c0.data_in_frame_27_3 ));
    CascadeMux I__16115 (
            .O(N__74499),
            .I(N__74496));
    InMux I__16114 (
            .O(N__74496),
            .I(N__74493));
    LocalMux I__16113 (
            .O(N__74493),
            .I(N__74489));
    InMux I__16112 (
            .O(N__74492),
            .I(N__74486));
    Span4Mux_h I__16111 (
            .O(N__74489),
            .I(N__74483));
    LocalMux I__16110 (
            .O(N__74486),
            .I(N__74480));
    Odrv4 I__16109 (
            .O(N__74483),
            .I(\c0.n33678 ));
    Odrv4 I__16108 (
            .O(N__74480),
            .I(\c0.n33678 ));
    CascadeMux I__16107 (
            .O(N__74475),
            .I(N__74471));
    InMux I__16106 (
            .O(N__74474),
            .I(N__74468));
    InMux I__16105 (
            .O(N__74471),
            .I(N__74465));
    LocalMux I__16104 (
            .O(N__74468),
            .I(N__74462));
    LocalMux I__16103 (
            .O(N__74465),
            .I(\c0.data_in_frame_29_5 ));
    Odrv4 I__16102 (
            .O(N__74462),
            .I(\c0.data_in_frame_29_5 ));
    InMux I__16101 (
            .O(N__74457),
            .I(N__74450));
    CascadeMux I__16100 (
            .O(N__74456),
            .I(N__74446));
    CascadeMux I__16099 (
            .O(N__74455),
            .I(N__74442));
    InMux I__16098 (
            .O(N__74454),
            .I(N__74436));
    InMux I__16097 (
            .O(N__74453),
            .I(N__74436));
    LocalMux I__16096 (
            .O(N__74450),
            .I(N__74433));
    InMux I__16095 (
            .O(N__74449),
            .I(N__74428));
    InMux I__16094 (
            .O(N__74446),
            .I(N__74428));
    InMux I__16093 (
            .O(N__74445),
            .I(N__74425));
    InMux I__16092 (
            .O(N__74442),
            .I(N__74420));
    InMux I__16091 (
            .O(N__74441),
            .I(N__74420));
    LocalMux I__16090 (
            .O(N__74436),
            .I(N__74417));
    Span4Mux_v I__16089 (
            .O(N__74433),
            .I(N__74414));
    LocalMux I__16088 (
            .O(N__74428),
            .I(N__74411));
    LocalMux I__16087 (
            .O(N__74425),
            .I(N__74408));
    LocalMux I__16086 (
            .O(N__74420),
            .I(N__74403));
    Span4Mux_v I__16085 (
            .O(N__74417),
            .I(N__74403));
    Span4Mux_v I__16084 (
            .O(N__74414),
            .I(N__74400));
    Span4Mux_v I__16083 (
            .O(N__74411),
            .I(N__74397));
    Span4Mux_v I__16082 (
            .O(N__74408),
            .I(N__74394));
    Span4Mux_v I__16081 (
            .O(N__74403),
            .I(N__74391));
    Span4Mux_h I__16080 (
            .O(N__74400),
            .I(N__74387));
    Span4Mux_v I__16079 (
            .O(N__74397),
            .I(N__74380));
    Span4Mux_v I__16078 (
            .O(N__74394),
            .I(N__74380));
    Span4Mux_h I__16077 (
            .O(N__74391),
            .I(N__74380));
    InMux I__16076 (
            .O(N__74390),
            .I(N__74377));
    Odrv4 I__16075 (
            .O(N__74387),
            .I(\c0.n12_adj_4518 ));
    Odrv4 I__16074 (
            .O(N__74380),
            .I(\c0.n12_adj_4518 ));
    LocalMux I__16073 (
            .O(N__74377),
            .I(\c0.n12_adj_4518 ));
    CascadeMux I__16072 (
            .O(N__74370),
            .I(N__74367));
    InMux I__16071 (
            .O(N__74367),
            .I(N__74363));
    InMux I__16070 (
            .O(N__74366),
            .I(N__74360));
    LocalMux I__16069 (
            .O(N__74363),
            .I(\c0.data_in_frame_29_3 ));
    LocalMux I__16068 (
            .O(N__74360),
            .I(\c0.data_in_frame_29_3 ));
    InMux I__16067 (
            .O(N__74355),
            .I(N__74351));
    InMux I__16066 (
            .O(N__74354),
            .I(N__74348));
    LocalMux I__16065 (
            .O(N__74351),
            .I(N__74342));
    LocalMux I__16064 (
            .O(N__74348),
            .I(N__74337));
    InMux I__16063 (
            .O(N__74347),
            .I(N__74330));
    InMux I__16062 (
            .O(N__74346),
            .I(N__74330));
    InMux I__16061 (
            .O(N__74345),
            .I(N__74330));
    Span4Mux_v I__16060 (
            .O(N__74342),
            .I(N__74327));
    InMux I__16059 (
            .O(N__74341),
            .I(N__74322));
    InMux I__16058 (
            .O(N__74340),
            .I(N__74322));
    Span4Mux_h I__16057 (
            .O(N__74337),
            .I(N__74319));
    LocalMux I__16056 (
            .O(N__74330),
            .I(N__74316));
    Span4Mux_h I__16055 (
            .O(N__74327),
            .I(N__74310));
    LocalMux I__16054 (
            .O(N__74322),
            .I(N__74310));
    Span4Mux_h I__16053 (
            .O(N__74319),
            .I(N__74307));
    Span4Mux_v I__16052 (
            .O(N__74316),
            .I(N__74304));
    InMux I__16051 (
            .O(N__74315),
            .I(N__74301));
    Odrv4 I__16050 (
            .O(N__74310),
            .I(\c0.n18971 ));
    Odrv4 I__16049 (
            .O(N__74307),
            .I(\c0.n18971 ));
    Odrv4 I__16048 (
            .O(N__74304),
            .I(\c0.n18971 ));
    LocalMux I__16047 (
            .O(N__74301),
            .I(\c0.n18971 ));
    CascadeMux I__16046 (
            .O(N__74292),
            .I(N__74287));
    CascadeMux I__16045 (
            .O(N__74291),
            .I(N__74283));
    InMux I__16044 (
            .O(N__74290),
            .I(N__74280));
    InMux I__16043 (
            .O(N__74287),
            .I(N__74274));
    InMux I__16042 (
            .O(N__74286),
            .I(N__74274));
    InMux I__16041 (
            .O(N__74283),
            .I(N__74270));
    LocalMux I__16040 (
            .O(N__74280),
            .I(N__74267));
    CascadeMux I__16039 (
            .O(N__74279),
            .I(N__74264));
    LocalMux I__16038 (
            .O(N__74274),
            .I(N__74260));
    InMux I__16037 (
            .O(N__74273),
            .I(N__74257));
    LocalMux I__16036 (
            .O(N__74270),
            .I(N__74252));
    Span4Mux_v I__16035 (
            .O(N__74267),
            .I(N__74252));
    InMux I__16034 (
            .O(N__74264),
            .I(N__74247));
    InMux I__16033 (
            .O(N__74263),
            .I(N__74247));
    Span4Mux_v I__16032 (
            .O(N__74260),
            .I(N__74237));
    LocalMux I__16031 (
            .O(N__74257),
            .I(N__74237));
    Span4Mux_h I__16030 (
            .O(N__74252),
            .I(N__74237));
    LocalMux I__16029 (
            .O(N__74247),
            .I(N__74237));
    InMux I__16028 (
            .O(N__74246),
            .I(N__74234));
    Span4Mux_h I__16027 (
            .O(N__74237),
            .I(N__74231));
    LocalMux I__16026 (
            .O(N__74234),
            .I(\c0.n33551 ));
    Odrv4 I__16025 (
            .O(N__74231),
            .I(\c0.n33551 ));
    InMux I__16024 (
            .O(N__74226),
            .I(N__74222));
    CascadeMux I__16023 (
            .O(N__74225),
            .I(N__74219));
    LocalMux I__16022 (
            .O(N__74222),
            .I(N__74215));
    InMux I__16021 (
            .O(N__74219),
            .I(N__74212));
    InMux I__16020 (
            .O(N__74218),
            .I(N__74209));
    Span4Mux_h I__16019 (
            .O(N__74215),
            .I(N__74204));
    LocalMux I__16018 (
            .O(N__74212),
            .I(N__74204));
    LocalMux I__16017 (
            .O(N__74209),
            .I(N__74201));
    Span4Mux_h I__16016 (
            .O(N__74204),
            .I(N__74198));
    Span4Mux_h I__16015 (
            .O(N__74201),
            .I(N__74195));
    Span4Mux_h I__16014 (
            .O(N__74198),
            .I(N__74192));
    Odrv4 I__16013 (
            .O(N__74195),
            .I(\c0.n32433 ));
    Odrv4 I__16012 (
            .O(N__74192),
            .I(\c0.n32433 ));
    InMux I__16011 (
            .O(N__74187),
            .I(N__74184));
    LocalMux I__16010 (
            .O(N__74184),
            .I(N__74181));
    Span4Mux_h I__16009 (
            .O(N__74181),
            .I(N__74178));
    Odrv4 I__16008 (
            .O(N__74178),
            .I(\c0.n33762 ));
    InMux I__16007 (
            .O(N__74175),
            .I(N__74168));
    InMux I__16006 (
            .O(N__74174),
            .I(N__74168));
    InMux I__16005 (
            .O(N__74173),
            .I(N__74165));
    LocalMux I__16004 (
            .O(N__74168),
            .I(N__74162));
    LocalMux I__16003 (
            .O(N__74165),
            .I(\c0.data_in_frame_25_0 ));
    Odrv4 I__16002 (
            .O(N__74162),
            .I(\c0.data_in_frame_25_0 ));
    InMux I__16001 (
            .O(N__74157),
            .I(N__74153));
    InMux I__16000 (
            .O(N__74156),
            .I(N__74148));
    LocalMux I__15999 (
            .O(N__74153),
            .I(N__74145));
    InMux I__15998 (
            .O(N__74152),
            .I(N__74142));
    InMux I__15997 (
            .O(N__74151),
            .I(N__74139));
    LocalMux I__15996 (
            .O(N__74148),
            .I(N__74136));
    Odrv4 I__15995 (
            .O(N__74145),
            .I(\c0.n32259 ));
    LocalMux I__15994 (
            .O(N__74142),
            .I(\c0.n32259 ));
    LocalMux I__15993 (
            .O(N__74139),
            .I(\c0.n32259 ));
    Odrv12 I__15992 (
            .O(N__74136),
            .I(\c0.n32259 ));
    InMux I__15991 (
            .O(N__74127),
            .I(N__74124));
    LocalMux I__15990 (
            .O(N__74124),
            .I(N__74120));
    CascadeMux I__15989 (
            .O(N__74123),
            .I(N__74116));
    Span4Mux_v I__15988 (
            .O(N__74120),
            .I(N__74113));
    CascadeMux I__15987 (
            .O(N__74119),
            .I(N__74110));
    InMux I__15986 (
            .O(N__74116),
            .I(N__74107));
    Span4Mux_h I__15985 (
            .O(N__74113),
            .I(N__74104));
    InMux I__15984 (
            .O(N__74110),
            .I(N__74101));
    LocalMux I__15983 (
            .O(N__74107),
            .I(\c0.data_in_frame_22_6 ));
    Odrv4 I__15982 (
            .O(N__74104),
            .I(\c0.data_in_frame_22_6 ));
    LocalMux I__15981 (
            .O(N__74101),
            .I(\c0.data_in_frame_22_6 ));
    InMux I__15980 (
            .O(N__74094),
            .I(N__74089));
    InMux I__15979 (
            .O(N__74093),
            .I(N__74086));
    InMux I__15978 (
            .O(N__74092),
            .I(N__74083));
    LocalMux I__15977 (
            .O(N__74089),
            .I(N__74080));
    LocalMux I__15976 (
            .O(N__74086),
            .I(N__74077));
    LocalMux I__15975 (
            .O(N__74083),
            .I(N__74074));
    Span4Mux_v I__15974 (
            .O(N__74080),
            .I(N__74069));
    Span4Mux_v I__15973 (
            .O(N__74077),
            .I(N__74069));
    Span4Mux_v I__15972 (
            .O(N__74074),
            .I(N__74066));
    Odrv4 I__15971 (
            .O(N__74069),
            .I(\c0.n32320 ));
    Odrv4 I__15970 (
            .O(N__74066),
            .I(\c0.n32320 ));
    InMux I__15969 (
            .O(N__74061),
            .I(N__74057));
    InMux I__15968 (
            .O(N__74060),
            .I(N__74054));
    LocalMux I__15967 (
            .O(N__74057),
            .I(N__74051));
    LocalMux I__15966 (
            .O(N__74054),
            .I(N__74046));
    Span4Mux_h I__15965 (
            .O(N__74051),
            .I(N__74046));
    Odrv4 I__15964 (
            .O(N__74046),
            .I(\c0.n33563 ));
    CascadeMux I__15963 (
            .O(N__74043),
            .I(N__74039));
    InMux I__15962 (
            .O(N__74042),
            .I(N__74035));
    InMux I__15961 (
            .O(N__74039),
            .I(N__74030));
    InMux I__15960 (
            .O(N__74038),
            .I(N__74030));
    LocalMux I__15959 (
            .O(N__74035),
            .I(\c0.data_in_frame_25_2 ));
    LocalMux I__15958 (
            .O(N__74030),
            .I(\c0.data_in_frame_25_2 ));
    CascadeMux I__15957 (
            .O(N__74025),
            .I(\c0.n33988_cascade_ ));
    CascadeMux I__15956 (
            .O(N__74022),
            .I(N__74019));
    InMux I__15955 (
            .O(N__74019),
            .I(N__74013));
    InMux I__15954 (
            .O(N__74018),
            .I(N__74013));
    LocalMux I__15953 (
            .O(N__74013),
            .I(N__74010));
    Span4Mux_v I__15952 (
            .O(N__74010),
            .I(N__74007));
    Odrv4 I__15951 (
            .O(N__74007),
            .I(\c0.n33536 ));
    InMux I__15950 (
            .O(N__74004),
            .I(N__74001));
    LocalMux I__15949 (
            .O(N__74001),
            .I(N__73997));
    CascadeMux I__15948 (
            .O(N__74000),
            .I(N__73994));
    Span4Mux_v I__15947 (
            .O(N__73997),
            .I(N__73991));
    InMux I__15946 (
            .O(N__73994),
            .I(N__73988));
    Span4Mux_h I__15945 (
            .O(N__73991),
            .I(N__73985));
    LocalMux I__15944 (
            .O(N__73988),
            .I(\c0.data_in_frame_28_2 ));
    Odrv4 I__15943 (
            .O(N__73985),
            .I(\c0.data_in_frame_28_2 ));
    CascadeMux I__15942 (
            .O(N__73980),
            .I(N__73974));
    InMux I__15941 (
            .O(N__73979),
            .I(N__73967));
    InMux I__15940 (
            .O(N__73978),
            .I(N__73967));
    InMux I__15939 (
            .O(N__73977),
            .I(N__73967));
    InMux I__15938 (
            .O(N__73974),
            .I(N__73964));
    LocalMux I__15937 (
            .O(N__73967),
            .I(N__73961));
    LocalMux I__15936 (
            .O(N__73964),
            .I(N__73958));
    Span4Mux_h I__15935 (
            .O(N__73961),
            .I(N__73955));
    Odrv4 I__15934 (
            .O(N__73958),
            .I(\c0.data_in_frame_27_5 ));
    Odrv4 I__15933 (
            .O(N__73955),
            .I(\c0.data_in_frame_27_5 ));
    CascadeMux I__15932 (
            .O(N__73950),
            .I(N__73943));
    CascadeMux I__15931 (
            .O(N__73949),
            .I(N__73938));
    CascadeMux I__15930 (
            .O(N__73948),
            .I(N__73931));
    CascadeMux I__15929 (
            .O(N__73947),
            .I(N__73923));
    InMux I__15928 (
            .O(N__73946),
            .I(N__73915));
    InMux I__15927 (
            .O(N__73943),
            .I(N__73915));
    InMux I__15926 (
            .O(N__73942),
            .I(N__73911));
    InMux I__15925 (
            .O(N__73941),
            .I(N__73903));
    InMux I__15924 (
            .O(N__73938),
            .I(N__73898));
    InMux I__15923 (
            .O(N__73937),
            .I(N__73898));
    InMux I__15922 (
            .O(N__73936),
            .I(N__73893));
    InMux I__15921 (
            .O(N__73935),
            .I(N__73893));
    InMux I__15920 (
            .O(N__73934),
            .I(N__73890));
    InMux I__15919 (
            .O(N__73931),
            .I(N__73887));
    InMux I__15918 (
            .O(N__73930),
            .I(N__73884));
    CascadeMux I__15917 (
            .O(N__73929),
            .I(N__73881));
    InMux I__15916 (
            .O(N__73928),
            .I(N__73875));
    InMux I__15915 (
            .O(N__73927),
            .I(N__73872));
    InMux I__15914 (
            .O(N__73926),
            .I(N__73869));
    InMux I__15913 (
            .O(N__73923),
            .I(N__73864));
    InMux I__15912 (
            .O(N__73922),
            .I(N__73864));
    CascadeMux I__15911 (
            .O(N__73921),
            .I(N__73861));
    InMux I__15910 (
            .O(N__73920),
            .I(N__73858));
    LocalMux I__15909 (
            .O(N__73915),
            .I(N__73855));
    InMux I__15908 (
            .O(N__73914),
            .I(N__73852));
    LocalMux I__15907 (
            .O(N__73911),
            .I(N__73849));
    CascadeMux I__15906 (
            .O(N__73910),
            .I(N__73844));
    InMux I__15905 (
            .O(N__73909),
            .I(N__73841));
    InMux I__15904 (
            .O(N__73908),
            .I(N__73834));
    InMux I__15903 (
            .O(N__73907),
            .I(N__73834));
    InMux I__15902 (
            .O(N__73906),
            .I(N__73834));
    LocalMux I__15901 (
            .O(N__73903),
            .I(N__73829));
    LocalMux I__15900 (
            .O(N__73898),
            .I(N__73829));
    LocalMux I__15899 (
            .O(N__73893),
            .I(N__73826));
    LocalMux I__15898 (
            .O(N__73890),
            .I(N__73823));
    LocalMux I__15897 (
            .O(N__73887),
            .I(N__73818));
    LocalMux I__15896 (
            .O(N__73884),
            .I(N__73818));
    InMux I__15895 (
            .O(N__73881),
            .I(N__73808));
    InMux I__15894 (
            .O(N__73880),
            .I(N__73808));
    InMux I__15893 (
            .O(N__73879),
            .I(N__73808));
    InMux I__15892 (
            .O(N__73878),
            .I(N__73808));
    LocalMux I__15891 (
            .O(N__73875),
            .I(N__73805));
    LocalMux I__15890 (
            .O(N__73872),
            .I(N__73802));
    LocalMux I__15889 (
            .O(N__73869),
            .I(N__73799));
    LocalMux I__15888 (
            .O(N__73864),
            .I(N__73796));
    InMux I__15887 (
            .O(N__73861),
            .I(N__73793));
    LocalMux I__15886 (
            .O(N__73858),
            .I(N__73788));
    Span4Mux_v I__15885 (
            .O(N__73855),
            .I(N__73788));
    LocalMux I__15884 (
            .O(N__73852),
            .I(N__73785));
    Span4Mux_h I__15883 (
            .O(N__73849),
            .I(N__73782));
    InMux I__15882 (
            .O(N__73848),
            .I(N__73778));
    InMux I__15881 (
            .O(N__73847),
            .I(N__73773));
    InMux I__15880 (
            .O(N__73844),
            .I(N__73773));
    LocalMux I__15879 (
            .O(N__73841),
            .I(N__73768));
    LocalMux I__15878 (
            .O(N__73834),
            .I(N__73768));
    Span4Mux_v I__15877 (
            .O(N__73829),
            .I(N__73765));
    Span4Mux_v I__15876 (
            .O(N__73826),
            .I(N__73760));
    Span4Mux_v I__15875 (
            .O(N__73823),
            .I(N__73760));
    Span4Mux_v I__15874 (
            .O(N__73818),
            .I(N__73757));
    InMux I__15873 (
            .O(N__73817),
            .I(N__73754));
    LocalMux I__15872 (
            .O(N__73808),
            .I(N__73747));
    Span4Mux_v I__15871 (
            .O(N__73805),
            .I(N__73747));
    Span4Mux_v I__15870 (
            .O(N__73802),
            .I(N__73747));
    Span4Mux_v I__15869 (
            .O(N__73799),
            .I(N__73742));
    Span4Mux_h I__15868 (
            .O(N__73796),
            .I(N__73742));
    LocalMux I__15867 (
            .O(N__73793),
            .I(N__73737));
    Span4Mux_h I__15866 (
            .O(N__73788),
            .I(N__73737));
    Span4Mux_h I__15865 (
            .O(N__73785),
            .I(N__73732));
    Span4Mux_h I__15864 (
            .O(N__73782),
            .I(N__73732));
    InMux I__15863 (
            .O(N__73781),
            .I(N__73729));
    LocalMux I__15862 (
            .O(N__73778),
            .I(N__73726));
    LocalMux I__15861 (
            .O(N__73773),
            .I(N__73723));
    Span4Mux_v I__15860 (
            .O(N__73768),
            .I(N__73714));
    Span4Mux_v I__15859 (
            .O(N__73765),
            .I(N__73714));
    Span4Mux_h I__15858 (
            .O(N__73760),
            .I(N__73714));
    Span4Mux_h I__15857 (
            .O(N__73757),
            .I(N__73714));
    LocalMux I__15856 (
            .O(N__73754),
            .I(N__73707));
    Span4Mux_v I__15855 (
            .O(N__73747),
            .I(N__73707));
    Span4Mux_h I__15854 (
            .O(N__73742),
            .I(N__73707));
    Span4Mux_v I__15853 (
            .O(N__73737),
            .I(N__73702));
    Span4Mux_h I__15852 (
            .O(N__73732),
            .I(N__73702));
    LocalMux I__15851 (
            .O(N__73729),
            .I(\c0.n9_adj_4631 ));
    Odrv4 I__15850 (
            .O(N__73726),
            .I(\c0.n9_adj_4631 ));
    Odrv12 I__15849 (
            .O(N__73723),
            .I(\c0.n9_adj_4631 ));
    Odrv4 I__15848 (
            .O(N__73714),
            .I(\c0.n9_adj_4631 ));
    Odrv4 I__15847 (
            .O(N__73707),
            .I(\c0.n9_adj_4631 ));
    Odrv4 I__15846 (
            .O(N__73702),
            .I(\c0.n9_adj_4631 ));
    InMux I__15845 (
            .O(N__73689),
            .I(N__73685));
    InMux I__15844 (
            .O(N__73688),
            .I(N__73682));
    LocalMux I__15843 (
            .O(N__73685),
            .I(N__73679));
    LocalMux I__15842 (
            .O(N__73682),
            .I(\c0.data_in_frame_28_0 ));
    Odrv4 I__15841 (
            .O(N__73679),
            .I(\c0.data_in_frame_28_0 ));
    CascadeMux I__15840 (
            .O(N__73674),
            .I(N__73668));
    InMux I__15839 (
            .O(N__73673),
            .I(N__73665));
    InMux I__15838 (
            .O(N__73672),
            .I(N__73662));
    InMux I__15837 (
            .O(N__73671),
            .I(N__73659));
    InMux I__15836 (
            .O(N__73668),
            .I(N__73656));
    LocalMux I__15835 (
            .O(N__73665),
            .I(N__73652));
    LocalMux I__15834 (
            .O(N__73662),
            .I(N__73647));
    LocalMux I__15833 (
            .O(N__73659),
            .I(N__73647));
    LocalMux I__15832 (
            .O(N__73656),
            .I(N__73644));
    InMux I__15831 (
            .O(N__73655),
            .I(N__73641));
    Span4Mux_v I__15830 (
            .O(N__73652),
            .I(N__73626));
    Span4Mux_v I__15829 (
            .O(N__73647),
            .I(N__73626));
    Span4Mux_v I__15828 (
            .O(N__73644),
            .I(N__73626));
    LocalMux I__15827 (
            .O(N__73641),
            .I(N__73618));
    InMux I__15826 (
            .O(N__73640),
            .I(N__73613));
    InMux I__15825 (
            .O(N__73639),
            .I(N__73606));
    InMux I__15824 (
            .O(N__73638),
            .I(N__73606));
    InMux I__15823 (
            .O(N__73637),
            .I(N__73606));
    InMux I__15822 (
            .O(N__73636),
            .I(N__73601));
    InMux I__15821 (
            .O(N__73635),
            .I(N__73601));
    InMux I__15820 (
            .O(N__73634),
            .I(N__73598));
    CascadeMux I__15819 (
            .O(N__73633),
            .I(N__73590));
    Span4Mux_h I__15818 (
            .O(N__73626),
            .I(N__73587));
    InMux I__15817 (
            .O(N__73625),
            .I(N__73584));
    InMux I__15816 (
            .O(N__73624),
            .I(N__73581));
    InMux I__15815 (
            .O(N__73623),
            .I(N__73578));
    InMux I__15814 (
            .O(N__73622),
            .I(N__73574));
    InMux I__15813 (
            .O(N__73621),
            .I(N__73571));
    Span4Mux_h I__15812 (
            .O(N__73618),
            .I(N__73568));
    InMux I__15811 (
            .O(N__73617),
            .I(N__73565));
    InMux I__15810 (
            .O(N__73616),
            .I(N__73562));
    LocalMux I__15809 (
            .O(N__73613),
            .I(N__73559));
    LocalMux I__15808 (
            .O(N__73606),
            .I(N__73556));
    LocalMux I__15807 (
            .O(N__73601),
            .I(N__73551));
    LocalMux I__15806 (
            .O(N__73598),
            .I(N__73551));
    InMux I__15805 (
            .O(N__73597),
            .I(N__73546));
    InMux I__15804 (
            .O(N__73596),
            .I(N__73546));
    InMux I__15803 (
            .O(N__73595),
            .I(N__73540));
    InMux I__15802 (
            .O(N__73594),
            .I(N__73540));
    InMux I__15801 (
            .O(N__73593),
            .I(N__73535));
    InMux I__15800 (
            .O(N__73590),
            .I(N__73535));
    Span4Mux_h I__15799 (
            .O(N__73587),
            .I(N__73528));
    LocalMux I__15798 (
            .O(N__73584),
            .I(N__73528));
    LocalMux I__15797 (
            .O(N__73581),
            .I(N__73528));
    LocalMux I__15796 (
            .O(N__73578),
            .I(N__73525));
    InMux I__15795 (
            .O(N__73577),
            .I(N__73519));
    LocalMux I__15794 (
            .O(N__73574),
            .I(N__73515));
    LocalMux I__15793 (
            .O(N__73571),
            .I(N__73508));
    Span4Mux_h I__15792 (
            .O(N__73568),
            .I(N__73508));
    LocalMux I__15791 (
            .O(N__73565),
            .I(N__73508));
    LocalMux I__15790 (
            .O(N__73562),
            .I(N__73501));
    Span4Mux_h I__15789 (
            .O(N__73559),
            .I(N__73501));
    Span4Mux_v I__15788 (
            .O(N__73556),
            .I(N__73501));
    Span4Mux_v I__15787 (
            .O(N__73551),
            .I(N__73498));
    LocalMux I__15786 (
            .O(N__73546),
            .I(N__73495));
    InMux I__15785 (
            .O(N__73545),
            .I(N__73492));
    LocalMux I__15784 (
            .O(N__73540),
            .I(N__73487));
    LocalMux I__15783 (
            .O(N__73535),
            .I(N__73487));
    Span4Mux_v I__15782 (
            .O(N__73528),
            .I(N__73484));
    Span4Mux_v I__15781 (
            .O(N__73525),
            .I(N__73481));
    InMux I__15780 (
            .O(N__73524),
            .I(N__73477));
    InMux I__15779 (
            .O(N__73523),
            .I(N__73474));
    InMux I__15778 (
            .O(N__73522),
            .I(N__73471));
    LocalMux I__15777 (
            .O(N__73519),
            .I(N__73468));
    InMux I__15776 (
            .O(N__73518),
            .I(N__73465));
    Sp12to4 I__15775 (
            .O(N__73515),
            .I(N__73460));
    Sp12to4 I__15774 (
            .O(N__73508),
            .I(N__73460));
    Span4Mux_v I__15773 (
            .O(N__73501),
            .I(N__73455));
    Span4Mux_v I__15772 (
            .O(N__73498),
            .I(N__73455));
    Span4Mux_v I__15771 (
            .O(N__73495),
            .I(N__73452));
    LocalMux I__15770 (
            .O(N__73492),
            .I(N__73449));
    Span4Mux_v I__15769 (
            .O(N__73487),
            .I(N__73442));
    Span4Mux_h I__15768 (
            .O(N__73484),
            .I(N__73442));
    Span4Mux_h I__15767 (
            .O(N__73481),
            .I(N__73442));
    InMux I__15766 (
            .O(N__73480),
            .I(N__73439));
    LocalMux I__15765 (
            .O(N__73477),
            .I(N__73434));
    LocalMux I__15764 (
            .O(N__73474),
            .I(N__73434));
    LocalMux I__15763 (
            .O(N__73471),
            .I(N__73429));
    Span12Mux_h I__15762 (
            .O(N__73468),
            .I(N__73429));
    LocalMux I__15761 (
            .O(N__73465),
            .I(N__73420));
    Span12Mux_v I__15760 (
            .O(N__73460),
            .I(N__73420));
    Sp12to4 I__15759 (
            .O(N__73455),
            .I(N__73420));
    Sp12to4 I__15758 (
            .O(N__73452),
            .I(N__73420));
    Span4Mux_v I__15757 (
            .O(N__73449),
            .I(N__73415));
    Span4Mux_h I__15756 (
            .O(N__73442),
            .I(N__73415));
    LocalMux I__15755 (
            .O(N__73439),
            .I(rx_data_6));
    Odrv4 I__15754 (
            .O(N__73434),
            .I(rx_data_6));
    Odrv12 I__15753 (
            .O(N__73429),
            .I(rx_data_6));
    Odrv12 I__15752 (
            .O(N__73420),
            .I(rx_data_6));
    Odrv4 I__15751 (
            .O(N__73415),
            .I(rx_data_6));
    InMux I__15750 (
            .O(N__73404),
            .I(N__73400));
    InMux I__15749 (
            .O(N__73403),
            .I(N__73396));
    LocalMux I__15748 (
            .O(N__73400),
            .I(N__73393));
    InMux I__15747 (
            .O(N__73399),
            .I(N__73390));
    LocalMux I__15746 (
            .O(N__73396),
            .I(N__73387));
    Span4Mux_h I__15745 (
            .O(N__73393),
            .I(N__73382));
    LocalMux I__15744 (
            .O(N__73390),
            .I(N__73382));
    Span4Mux_h I__15743 (
            .O(N__73387),
            .I(N__73379));
    Span4Mux_h I__15742 (
            .O(N__73382),
            .I(N__73376));
    Odrv4 I__15741 (
            .O(N__73379),
            .I(\c0.n33539 ));
    Odrv4 I__15740 (
            .O(N__73376),
            .I(\c0.n33539 ));
    InMux I__15739 (
            .O(N__73371),
            .I(N__73368));
    LocalMux I__15738 (
            .O(N__73368),
            .I(N__73364));
    InMux I__15737 (
            .O(N__73367),
            .I(N__73361));
    Span4Mux_v I__15736 (
            .O(N__73364),
            .I(N__73358));
    LocalMux I__15735 (
            .O(N__73361),
            .I(\c0.n33933 ));
    Odrv4 I__15734 (
            .O(N__73358),
            .I(\c0.n33933 ));
    CascadeMux I__15733 (
            .O(N__73353),
            .I(N__73348));
    InMux I__15732 (
            .O(N__73352),
            .I(N__73344));
    InMux I__15731 (
            .O(N__73351),
            .I(N__73341));
    InMux I__15730 (
            .O(N__73348),
            .I(N__73338));
    InMux I__15729 (
            .O(N__73347),
            .I(N__73335));
    LocalMux I__15728 (
            .O(N__73344),
            .I(\c0.data_in_frame_27_1 ));
    LocalMux I__15727 (
            .O(N__73341),
            .I(\c0.data_in_frame_27_1 ));
    LocalMux I__15726 (
            .O(N__73338),
            .I(\c0.data_in_frame_27_1 ));
    LocalMux I__15725 (
            .O(N__73335),
            .I(\c0.data_in_frame_27_1 ));
    CascadeMux I__15724 (
            .O(N__73326),
            .I(N__73323));
    InMux I__15723 (
            .O(N__73323),
            .I(N__73318));
    InMux I__15722 (
            .O(N__73322),
            .I(N__73313));
    InMux I__15721 (
            .O(N__73321),
            .I(N__73313));
    LocalMux I__15720 (
            .O(N__73318),
            .I(N__73307));
    LocalMux I__15719 (
            .O(N__73313),
            .I(N__73307));
    InMux I__15718 (
            .O(N__73312),
            .I(N__73304));
    Odrv12 I__15717 (
            .O(N__73307),
            .I(\c0.data_in_frame_21_1 ));
    LocalMux I__15716 (
            .O(N__73304),
            .I(\c0.data_in_frame_21_1 ));
    InMux I__15715 (
            .O(N__73299),
            .I(N__73293));
    InMux I__15714 (
            .O(N__73298),
            .I(N__73293));
    LocalMux I__15713 (
            .O(N__73293),
            .I(N__73288));
    CascadeMux I__15712 (
            .O(N__73292),
            .I(N__73285));
    CascadeMux I__15711 (
            .O(N__73291),
            .I(N__73282));
    Span4Mux_v I__15710 (
            .O(N__73288),
            .I(N__73279));
    InMux I__15709 (
            .O(N__73285),
            .I(N__73274));
    InMux I__15708 (
            .O(N__73282),
            .I(N__73274));
    Odrv4 I__15707 (
            .O(N__73279),
            .I(\c0.data_in_frame_21_2 ));
    LocalMux I__15706 (
            .O(N__73274),
            .I(\c0.data_in_frame_21_2 ));
    InMux I__15705 (
            .O(N__73269),
            .I(N__73265));
    InMux I__15704 (
            .O(N__73268),
            .I(N__73262));
    LocalMux I__15703 (
            .O(N__73265),
            .I(\c0.data_in_frame_29_2 ));
    LocalMux I__15702 (
            .O(N__73262),
            .I(\c0.data_in_frame_29_2 ));
    CascadeMux I__15701 (
            .O(N__73257),
            .I(N__73253));
    CascadeMux I__15700 (
            .O(N__73256),
            .I(N__73250));
    InMux I__15699 (
            .O(N__73253),
            .I(N__73247));
    InMux I__15698 (
            .O(N__73250),
            .I(N__73244));
    LocalMux I__15697 (
            .O(N__73247),
            .I(N__73241));
    LocalMux I__15696 (
            .O(N__73244),
            .I(\c0.data_in_frame_29_1 ));
    Odrv4 I__15695 (
            .O(N__73241),
            .I(\c0.data_in_frame_29_1 ));
    CascadeMux I__15694 (
            .O(N__73236),
            .I(N__73233));
    InMux I__15693 (
            .O(N__73233),
            .I(N__73228));
    InMux I__15692 (
            .O(N__73232),
            .I(N__73225));
    InMux I__15691 (
            .O(N__73231),
            .I(N__73222));
    LocalMux I__15690 (
            .O(N__73228),
            .I(N__73218));
    LocalMux I__15689 (
            .O(N__73225),
            .I(N__73215));
    LocalMux I__15688 (
            .O(N__73222),
            .I(N__73212));
    InMux I__15687 (
            .O(N__73221),
            .I(N__73208));
    Span12Mux_h I__15686 (
            .O(N__73218),
            .I(N__73205));
    Span4Mux_h I__15685 (
            .O(N__73215),
            .I(N__73202));
    Span4Mux_v I__15684 (
            .O(N__73212),
            .I(N__73199));
    InMux I__15683 (
            .O(N__73211),
            .I(N__73196));
    LocalMux I__15682 (
            .O(N__73208),
            .I(encoder0_position_8));
    Odrv12 I__15681 (
            .O(N__73205),
            .I(encoder0_position_8));
    Odrv4 I__15680 (
            .O(N__73202),
            .I(encoder0_position_8));
    Odrv4 I__15679 (
            .O(N__73199),
            .I(encoder0_position_8));
    LocalMux I__15678 (
            .O(N__73196),
            .I(encoder0_position_8));
    InMux I__15677 (
            .O(N__73185),
            .I(N__73182));
    LocalMux I__15676 (
            .O(N__73182),
            .I(N__73179));
    Span4Mux_h I__15675 (
            .O(N__73179),
            .I(N__73176));
    Odrv4 I__15674 (
            .O(N__73176),
            .I(n2341));
    CascadeMux I__15673 (
            .O(N__73173),
            .I(N__73170));
    InMux I__15672 (
            .O(N__73170),
            .I(N__73166));
    CascadeMux I__15671 (
            .O(N__73169),
            .I(N__73163));
    LocalMux I__15670 (
            .O(N__73166),
            .I(N__73159));
    InMux I__15669 (
            .O(N__73163),
            .I(N__73156));
    InMux I__15668 (
            .O(N__73162),
            .I(N__73153));
    Span12Mux_h I__15667 (
            .O(N__73159),
            .I(N__73148));
    LocalMux I__15666 (
            .O(N__73156),
            .I(N__73148));
    LocalMux I__15665 (
            .O(N__73153),
            .I(\c0.data_in_frame_26_3 ));
    Odrv12 I__15664 (
            .O(N__73148),
            .I(\c0.data_in_frame_26_3 ));
    CascadeMux I__15663 (
            .O(N__73143),
            .I(N__73140));
    InMux I__15662 (
            .O(N__73140),
            .I(N__73137));
    LocalMux I__15661 (
            .O(N__73137),
            .I(N__73134));
    Span4Mux_v I__15660 (
            .O(N__73134),
            .I(N__73128));
    InMux I__15659 (
            .O(N__73133),
            .I(N__73123));
    InMux I__15658 (
            .O(N__73132),
            .I(N__73123));
    InMux I__15657 (
            .O(N__73131),
            .I(N__73120));
    Span4Mux_h I__15656 (
            .O(N__73128),
            .I(N__73115));
    LocalMux I__15655 (
            .O(N__73123),
            .I(N__73115));
    LocalMux I__15654 (
            .O(N__73120),
            .I(\c0.data_in_frame_25_3 ));
    Odrv4 I__15653 (
            .O(N__73115),
            .I(\c0.data_in_frame_25_3 ));
    InMux I__15652 (
            .O(N__73110),
            .I(N__73107));
    LocalMux I__15651 (
            .O(N__73107),
            .I(N__73104));
    Span4Mux_h I__15650 (
            .O(N__73104),
            .I(N__73101));
    Odrv4 I__15649 (
            .O(N__73101),
            .I(n2320));
    CascadeMux I__15648 (
            .O(N__73098),
            .I(N__73094));
    CascadeMux I__15647 (
            .O(N__73097),
            .I(N__73091));
    InMux I__15646 (
            .O(N__73094),
            .I(N__73087));
    InMux I__15645 (
            .O(N__73091),
            .I(N__73084));
    CascadeMux I__15644 (
            .O(N__73090),
            .I(N__73081));
    LocalMux I__15643 (
            .O(N__73087),
            .I(N__73076));
    LocalMux I__15642 (
            .O(N__73084),
            .I(N__73073));
    InMux I__15641 (
            .O(N__73081),
            .I(N__73070));
    InMux I__15640 (
            .O(N__73080),
            .I(N__73067));
    InMux I__15639 (
            .O(N__73079),
            .I(N__73064));
    Span4Mux_h I__15638 (
            .O(N__73076),
            .I(N__73055));
    Span4Mux_h I__15637 (
            .O(N__73073),
            .I(N__73055));
    LocalMux I__15636 (
            .O(N__73070),
            .I(N__73055));
    LocalMux I__15635 (
            .O(N__73067),
            .I(N__73055));
    LocalMux I__15634 (
            .O(N__73064),
            .I(encoder0_position_25));
    Odrv4 I__15633 (
            .O(N__73055),
            .I(encoder0_position_25));
    InMux I__15632 (
            .O(N__73050),
            .I(N__73047));
    LocalMux I__15631 (
            .O(N__73047),
            .I(N__73042));
    CascadeMux I__15630 (
            .O(N__73046),
            .I(N__73033));
    CascadeMux I__15629 (
            .O(N__73045),
            .I(N__73003));
    Span4Mux_v I__15628 (
            .O(N__73042),
            .I(N__73000));
    InMux I__15627 (
            .O(N__73041),
            .I(N__72995));
    InMux I__15626 (
            .O(N__73040),
            .I(N__72995));
    InMux I__15625 (
            .O(N__73039),
            .I(N__72992));
    InMux I__15624 (
            .O(N__73038),
            .I(N__72987));
    InMux I__15623 (
            .O(N__73037),
            .I(N__72987));
    InMux I__15622 (
            .O(N__73036),
            .I(N__72979));
    InMux I__15621 (
            .O(N__73033),
            .I(N__72976));
    InMux I__15620 (
            .O(N__73032),
            .I(N__72972));
    InMux I__15619 (
            .O(N__73031),
            .I(N__72969));
    InMux I__15618 (
            .O(N__73030),
            .I(N__72964));
    InMux I__15617 (
            .O(N__73029),
            .I(N__72964));
    InMux I__15616 (
            .O(N__73028),
            .I(N__72961));
    InMux I__15615 (
            .O(N__73027),
            .I(N__72958));
    InMux I__15614 (
            .O(N__73026),
            .I(N__72955));
    InMux I__15613 (
            .O(N__73025),
            .I(N__72944));
    InMux I__15612 (
            .O(N__73024),
            .I(N__72944));
    InMux I__15611 (
            .O(N__73023),
            .I(N__72944));
    InMux I__15610 (
            .O(N__73022),
            .I(N__72944));
    InMux I__15609 (
            .O(N__73021),
            .I(N__72944));
    InMux I__15608 (
            .O(N__73020),
            .I(N__72937));
    InMux I__15607 (
            .O(N__73019),
            .I(N__72937));
    InMux I__15606 (
            .O(N__73018),
            .I(N__72937));
    InMux I__15605 (
            .O(N__73017),
            .I(N__72926));
    InMux I__15604 (
            .O(N__73016),
            .I(N__72926));
    InMux I__15603 (
            .O(N__73015),
            .I(N__72926));
    InMux I__15602 (
            .O(N__73014),
            .I(N__72926));
    InMux I__15601 (
            .O(N__73013),
            .I(N__72926));
    InMux I__15600 (
            .O(N__73012),
            .I(N__72913));
    InMux I__15599 (
            .O(N__73011),
            .I(N__72913));
    InMux I__15598 (
            .O(N__73010),
            .I(N__72913));
    InMux I__15597 (
            .O(N__73009),
            .I(N__72913));
    InMux I__15596 (
            .O(N__73008),
            .I(N__72913));
    InMux I__15595 (
            .O(N__73007),
            .I(N__72910));
    CascadeMux I__15594 (
            .O(N__73006),
            .I(N__72907));
    InMux I__15593 (
            .O(N__73003),
            .I(N__72904));
    Span4Mux_h I__15592 (
            .O(N__73000),
            .I(N__72897));
    LocalMux I__15591 (
            .O(N__72995),
            .I(N__72897));
    LocalMux I__15590 (
            .O(N__72992),
            .I(N__72892));
    LocalMux I__15589 (
            .O(N__72987),
            .I(N__72892));
    InMux I__15588 (
            .O(N__72986),
            .I(N__72889));
    InMux I__15587 (
            .O(N__72985),
            .I(N__72886));
    InMux I__15586 (
            .O(N__72984),
            .I(N__72881));
    InMux I__15585 (
            .O(N__72983),
            .I(N__72881));
    InMux I__15584 (
            .O(N__72982),
            .I(N__72876));
    LocalMux I__15583 (
            .O(N__72979),
            .I(N__72871));
    LocalMux I__15582 (
            .O(N__72976),
            .I(N__72871));
    InMux I__15581 (
            .O(N__72975),
            .I(N__72863));
    LocalMux I__15580 (
            .O(N__72972),
            .I(N__72860));
    LocalMux I__15579 (
            .O(N__72969),
            .I(N__72851));
    LocalMux I__15578 (
            .O(N__72964),
            .I(N__72851));
    LocalMux I__15577 (
            .O(N__72961),
            .I(N__72851));
    LocalMux I__15576 (
            .O(N__72958),
            .I(N__72851));
    LocalMux I__15575 (
            .O(N__72955),
            .I(N__72842));
    LocalMux I__15574 (
            .O(N__72944),
            .I(N__72842));
    LocalMux I__15573 (
            .O(N__72937),
            .I(N__72842));
    LocalMux I__15572 (
            .O(N__72926),
            .I(N__72842));
    InMux I__15571 (
            .O(N__72925),
            .I(N__72837));
    InMux I__15570 (
            .O(N__72924),
            .I(N__72837));
    LocalMux I__15569 (
            .O(N__72913),
            .I(N__72834));
    LocalMux I__15568 (
            .O(N__72910),
            .I(N__72831));
    InMux I__15567 (
            .O(N__72907),
            .I(N__72828));
    LocalMux I__15566 (
            .O(N__72904),
            .I(N__72825));
    InMux I__15565 (
            .O(N__72903),
            .I(N__72820));
    InMux I__15564 (
            .O(N__72902),
            .I(N__72820));
    Span4Mux_v I__15563 (
            .O(N__72897),
            .I(N__72817));
    Span4Mux_v I__15562 (
            .O(N__72892),
            .I(N__72812));
    LocalMux I__15561 (
            .O(N__72889),
            .I(N__72812));
    LocalMux I__15560 (
            .O(N__72886),
            .I(N__72807));
    LocalMux I__15559 (
            .O(N__72881),
            .I(N__72807));
    CascadeMux I__15558 (
            .O(N__72880),
            .I(N__72804));
    CascadeMux I__15557 (
            .O(N__72879),
            .I(N__72800));
    LocalMux I__15556 (
            .O(N__72876),
            .I(N__72796));
    Span4Mux_v I__15555 (
            .O(N__72871),
            .I(N__72793));
    InMux I__15554 (
            .O(N__72870),
            .I(N__72790));
    InMux I__15553 (
            .O(N__72869),
            .I(N__72785));
    InMux I__15552 (
            .O(N__72868),
            .I(N__72785));
    InMux I__15551 (
            .O(N__72867),
            .I(N__72780));
    InMux I__15550 (
            .O(N__72866),
            .I(N__72780));
    LocalMux I__15549 (
            .O(N__72863),
            .I(N__72771));
    Span4Mux_v I__15548 (
            .O(N__72860),
            .I(N__72771));
    Span4Mux_v I__15547 (
            .O(N__72851),
            .I(N__72771));
    Span4Mux_v I__15546 (
            .O(N__72842),
            .I(N__72771));
    LocalMux I__15545 (
            .O(N__72837),
            .I(N__72766));
    Span4Mux_v I__15544 (
            .O(N__72834),
            .I(N__72766));
    Span4Mux_v I__15543 (
            .O(N__72831),
            .I(N__72763));
    LocalMux I__15542 (
            .O(N__72828),
            .I(N__72750));
    Span4Mux_h I__15541 (
            .O(N__72825),
            .I(N__72750));
    LocalMux I__15540 (
            .O(N__72820),
            .I(N__72750));
    Span4Mux_h I__15539 (
            .O(N__72817),
            .I(N__72750));
    Span4Mux_h I__15538 (
            .O(N__72812),
            .I(N__72750));
    Span4Mux_v I__15537 (
            .O(N__72807),
            .I(N__72750));
    InMux I__15536 (
            .O(N__72804),
            .I(N__72745));
    InMux I__15535 (
            .O(N__72803),
            .I(N__72745));
    InMux I__15534 (
            .O(N__72800),
            .I(N__72740));
    InMux I__15533 (
            .O(N__72799),
            .I(N__72740));
    Span4Mux_h I__15532 (
            .O(N__72796),
            .I(N__72735));
    Span4Mux_h I__15531 (
            .O(N__72793),
            .I(N__72735));
    LocalMux I__15530 (
            .O(N__72790),
            .I(N__72726));
    LocalMux I__15529 (
            .O(N__72785),
            .I(N__72726));
    LocalMux I__15528 (
            .O(N__72780),
            .I(N__72726));
    Span4Mux_h I__15527 (
            .O(N__72771),
            .I(N__72726));
    Span4Mux_v I__15526 (
            .O(N__72766),
            .I(N__72719));
    Span4Mux_v I__15525 (
            .O(N__72763),
            .I(N__72719));
    Span4Mux_v I__15524 (
            .O(N__72750),
            .I(N__72719));
    LocalMux I__15523 (
            .O(N__72745),
            .I(\c0.n33233 ));
    LocalMux I__15522 (
            .O(N__72740),
            .I(\c0.n33233 ));
    Odrv4 I__15521 (
            .O(N__72735),
            .I(\c0.n33233 ));
    Odrv4 I__15520 (
            .O(N__72726),
            .I(\c0.n33233 ));
    Odrv4 I__15519 (
            .O(N__72719),
            .I(\c0.n33233 ));
    InMux I__15518 (
            .O(N__72708),
            .I(N__72705));
    LocalMux I__15517 (
            .O(N__72705),
            .I(N__72701));
    InMux I__15516 (
            .O(N__72704),
            .I(N__72697));
    Span4Mux_v I__15515 (
            .O(N__72701),
            .I(N__72694));
    InMux I__15514 (
            .O(N__72700),
            .I(N__72691));
    LocalMux I__15513 (
            .O(N__72697),
            .I(\c0.data_in_frame_22_3 ));
    Odrv4 I__15512 (
            .O(N__72694),
            .I(\c0.data_in_frame_22_3 ));
    LocalMux I__15511 (
            .O(N__72691),
            .I(\c0.data_in_frame_22_3 ));
    InMux I__15510 (
            .O(N__72684),
            .I(N__72681));
    LocalMux I__15509 (
            .O(N__72681),
            .I(N__72678));
    Span4Mux_h I__15508 (
            .O(N__72678),
            .I(N__72675));
    Odrv4 I__15507 (
            .O(N__72675),
            .I(n2328));
    CascadeMux I__15506 (
            .O(N__72672),
            .I(N__72669));
    InMux I__15505 (
            .O(N__72669),
            .I(N__72666));
    LocalMux I__15504 (
            .O(N__72666),
            .I(\c0.n10_adj_4547 ));
    InMux I__15503 (
            .O(N__72663),
            .I(N__72655));
    InMux I__15502 (
            .O(N__72662),
            .I(N__72655));
    CascadeMux I__15501 (
            .O(N__72661),
            .I(N__72652));
    InMux I__15500 (
            .O(N__72660),
            .I(N__72647));
    LocalMux I__15499 (
            .O(N__72655),
            .I(N__72644));
    InMux I__15498 (
            .O(N__72652),
            .I(N__72641));
    InMux I__15497 (
            .O(N__72651),
            .I(N__72636));
    InMux I__15496 (
            .O(N__72650),
            .I(N__72636));
    LocalMux I__15495 (
            .O(N__72647),
            .I(N__72631));
    Span4Mux_v I__15494 (
            .O(N__72644),
            .I(N__72631));
    LocalMux I__15493 (
            .O(N__72641),
            .I(control_mode_6));
    LocalMux I__15492 (
            .O(N__72636),
            .I(control_mode_6));
    Odrv4 I__15491 (
            .O(N__72631),
            .I(control_mode_6));
    InMux I__15490 (
            .O(N__72624),
            .I(N__72618));
    InMux I__15489 (
            .O(N__72623),
            .I(N__72618));
    LocalMux I__15488 (
            .O(N__72618),
            .I(N__72615));
    Odrv4 I__15487 (
            .O(N__72615),
            .I(\c0.n33414 ));
    InMux I__15486 (
            .O(N__72612),
            .I(N__72609));
    LocalMux I__15485 (
            .O(N__72609),
            .I(N__72606));
    Span4Mux_v I__15484 (
            .O(N__72606),
            .I(N__72603));
    Odrv4 I__15483 (
            .O(N__72603),
            .I(n2322));
    CascadeMux I__15482 (
            .O(N__72600),
            .I(N__72597));
    InMux I__15481 (
            .O(N__72597),
            .I(N__72593));
    CascadeMux I__15480 (
            .O(N__72596),
            .I(N__72590));
    LocalMux I__15479 (
            .O(N__72593),
            .I(N__72585));
    InMux I__15478 (
            .O(N__72590),
            .I(N__72582));
    InMux I__15477 (
            .O(N__72589),
            .I(N__72579));
    CascadeMux I__15476 (
            .O(N__72588),
            .I(N__72576));
    Span4Mux_v I__15475 (
            .O(N__72585),
            .I(N__72572));
    LocalMux I__15474 (
            .O(N__72582),
            .I(N__72569));
    LocalMux I__15473 (
            .O(N__72579),
            .I(N__72566));
    InMux I__15472 (
            .O(N__72576),
            .I(N__72563));
    InMux I__15471 (
            .O(N__72575),
            .I(N__72560));
    Span4Mux_h I__15470 (
            .O(N__72572),
            .I(N__72557));
    Span4Mux_h I__15469 (
            .O(N__72569),
            .I(N__72550));
    Span4Mux_v I__15468 (
            .O(N__72566),
            .I(N__72550));
    LocalMux I__15467 (
            .O(N__72563),
            .I(N__72550));
    LocalMux I__15466 (
            .O(N__72560),
            .I(encoder0_position_23));
    Odrv4 I__15465 (
            .O(N__72557),
            .I(encoder0_position_23));
    Odrv4 I__15464 (
            .O(N__72550),
            .I(encoder0_position_23));
    InMux I__15463 (
            .O(N__72543),
            .I(N__72540));
    LocalMux I__15462 (
            .O(N__72540),
            .I(N__72537));
    Span4Mux_v I__15461 (
            .O(N__72537),
            .I(N__72534));
    Odrv4 I__15460 (
            .O(N__72534),
            .I(n2336));
    InMux I__15459 (
            .O(N__72531),
            .I(N__72528));
    LocalMux I__15458 (
            .O(N__72528),
            .I(N__72525));
    Odrv4 I__15457 (
            .O(N__72525),
            .I(n2329));
    InMux I__15456 (
            .O(N__72522),
            .I(N__72516));
    InMux I__15455 (
            .O(N__72521),
            .I(N__72516));
    LocalMux I__15454 (
            .O(N__72516),
            .I(N__72512));
    CascadeMux I__15453 (
            .O(N__72515),
            .I(N__72509));
    Span4Mux_h I__15452 (
            .O(N__72512),
            .I(N__72506));
    InMux I__15451 (
            .O(N__72509),
            .I(N__72503));
    Span4Mux_h I__15450 (
            .O(N__72506),
            .I(N__72500));
    LocalMux I__15449 (
            .O(N__72503),
            .I(\c0.data_in_frame_22_4 ));
    Odrv4 I__15448 (
            .O(N__72500),
            .I(\c0.data_in_frame_22_4 ));
    CascadeMux I__15447 (
            .O(N__72495),
            .I(\c0.data_out_frame_29__7__N_738_cascade_ ));
    InMux I__15446 (
            .O(N__72492),
            .I(N__72489));
    LocalMux I__15445 (
            .O(N__72489),
            .I(\c0.n33389 ));
    InMux I__15444 (
            .O(N__72486),
            .I(N__72483));
    LocalMux I__15443 (
            .O(N__72483),
            .I(\c0.n22 ));
    CascadeMux I__15442 (
            .O(N__72480),
            .I(\c0.n33579_cascade_ ));
    InMux I__15441 (
            .O(N__72477),
            .I(N__72474));
    LocalMux I__15440 (
            .O(N__72474),
            .I(N__72471));
    Odrv12 I__15439 (
            .O(N__72471),
            .I(n2343));
    CascadeMux I__15438 (
            .O(N__72468),
            .I(N__72465));
    InMux I__15437 (
            .O(N__72465),
            .I(N__72461));
    InMux I__15436 (
            .O(N__72464),
            .I(N__72457));
    LocalMux I__15435 (
            .O(N__72461),
            .I(N__72451));
    InMux I__15434 (
            .O(N__72460),
            .I(N__72448));
    LocalMux I__15433 (
            .O(N__72457),
            .I(N__72445));
    InMux I__15432 (
            .O(N__72456),
            .I(N__72438));
    InMux I__15431 (
            .O(N__72455),
            .I(N__72438));
    InMux I__15430 (
            .O(N__72454),
            .I(N__72438));
    Odrv12 I__15429 (
            .O(N__72451),
            .I(control_mode_7));
    LocalMux I__15428 (
            .O(N__72448),
            .I(control_mode_7));
    Odrv4 I__15427 (
            .O(N__72445),
            .I(control_mode_7));
    LocalMux I__15426 (
            .O(N__72438),
            .I(control_mode_7));
    InMux I__15425 (
            .O(N__72429),
            .I(N__72426));
    LocalMux I__15424 (
            .O(N__72426),
            .I(N__72422));
    InMux I__15423 (
            .O(N__72425),
            .I(N__72419));
    Span4Mux_h I__15422 (
            .O(N__72422),
            .I(N__72412));
    LocalMux I__15421 (
            .O(N__72419),
            .I(N__72409));
    InMux I__15420 (
            .O(N__72418),
            .I(N__72406));
    InMux I__15419 (
            .O(N__72417),
            .I(N__72401));
    InMux I__15418 (
            .O(N__72416),
            .I(N__72401));
    InMux I__15417 (
            .O(N__72415),
            .I(N__72398));
    Span4Mux_h I__15416 (
            .O(N__72412),
            .I(N__72393));
    Span4Mux_h I__15415 (
            .O(N__72409),
            .I(N__72393));
    LocalMux I__15414 (
            .O(N__72406),
            .I(N__72388));
    LocalMux I__15413 (
            .O(N__72401),
            .I(N__72388));
    LocalMux I__15412 (
            .O(N__72398),
            .I(data_in_frame_1_5));
    Odrv4 I__15411 (
            .O(N__72393),
            .I(data_in_frame_1_5));
    Odrv4 I__15410 (
            .O(N__72388),
            .I(data_in_frame_1_5));
    InMux I__15409 (
            .O(N__72381),
            .I(N__72376));
    InMux I__15408 (
            .O(N__72380),
            .I(N__72373));
    InMux I__15407 (
            .O(N__72379),
            .I(N__72370));
    LocalMux I__15406 (
            .O(N__72376),
            .I(N__72367));
    LocalMux I__15405 (
            .O(N__72373),
            .I(N__72363));
    LocalMux I__15404 (
            .O(N__72370),
            .I(N__72359));
    Span12Mux_h I__15403 (
            .O(N__72367),
            .I(N__72356));
    InMux I__15402 (
            .O(N__72366),
            .I(N__72353));
    Span4Mux_h I__15401 (
            .O(N__72363),
            .I(N__72350));
    InMux I__15400 (
            .O(N__72362),
            .I(N__72347));
    Span4Mux_v I__15399 (
            .O(N__72359),
            .I(N__72344));
    Odrv12 I__15398 (
            .O(N__72356),
            .I(encoder0_position_10));
    LocalMux I__15397 (
            .O(N__72353),
            .I(encoder0_position_10));
    Odrv4 I__15396 (
            .O(N__72350),
            .I(encoder0_position_10));
    LocalMux I__15395 (
            .O(N__72347),
            .I(encoder0_position_10));
    Odrv4 I__15394 (
            .O(N__72344),
            .I(encoder0_position_10));
    CascadeMux I__15393 (
            .O(N__72333),
            .I(\c0.n33493_cascade_ ));
    InMux I__15392 (
            .O(N__72330),
            .I(N__72326));
    InMux I__15391 (
            .O(N__72329),
            .I(N__72323));
    LocalMux I__15390 (
            .O(N__72326),
            .I(N__72318));
    LocalMux I__15389 (
            .O(N__72323),
            .I(N__72318));
    Odrv4 I__15388 (
            .O(N__72318),
            .I(\c0.n33749 ));
    CascadeMux I__15387 (
            .O(N__72315),
            .I(N__72312));
    InMux I__15386 (
            .O(N__72312),
            .I(N__72309));
    LocalMux I__15385 (
            .O(N__72309),
            .I(N__72305));
    InMux I__15384 (
            .O(N__72308),
            .I(N__72299));
    Span4Mux_v I__15383 (
            .O(N__72305),
            .I(N__72296));
    InMux I__15382 (
            .O(N__72304),
            .I(N__72293));
    InMux I__15381 (
            .O(N__72303),
            .I(N__72288));
    InMux I__15380 (
            .O(N__72302),
            .I(N__72288));
    LocalMux I__15379 (
            .O(N__72299),
            .I(control_mode_1));
    Odrv4 I__15378 (
            .O(N__72296),
            .I(control_mode_1));
    LocalMux I__15377 (
            .O(N__72293),
            .I(control_mode_1));
    LocalMux I__15376 (
            .O(N__72288),
            .I(control_mode_1));
    InMux I__15375 (
            .O(N__72279),
            .I(N__72275));
    InMux I__15374 (
            .O(N__72278),
            .I(N__72270));
    LocalMux I__15373 (
            .O(N__72275),
            .I(N__72267));
    InMux I__15372 (
            .O(N__72274),
            .I(N__72264));
    InMux I__15371 (
            .O(N__72273),
            .I(N__72261));
    LocalMux I__15370 (
            .O(N__72270),
            .I(N__72253));
    Span4Mux_v I__15369 (
            .O(N__72267),
            .I(N__72253));
    LocalMux I__15368 (
            .O(N__72264),
            .I(N__72253));
    LocalMux I__15367 (
            .O(N__72261),
            .I(N__72250));
    InMux I__15366 (
            .O(N__72260),
            .I(N__72247));
    Span4Mux_h I__15365 (
            .O(N__72253),
            .I(N__72244));
    Odrv12 I__15364 (
            .O(N__72250),
            .I(encoder1_position_26));
    LocalMux I__15363 (
            .O(N__72247),
            .I(encoder1_position_26));
    Odrv4 I__15362 (
            .O(N__72244),
            .I(encoder1_position_26));
    CascadeMux I__15361 (
            .O(N__72237),
            .I(\c0.n33432_cascade_ ));
    InMux I__15360 (
            .O(N__72234),
            .I(N__72231));
    LocalMux I__15359 (
            .O(N__72231),
            .I(N__72228));
    Span4Mux_h I__15358 (
            .O(N__72228),
            .I(N__72225));
    Odrv4 I__15357 (
            .O(N__72225),
            .I(n2248));
    InMux I__15356 (
            .O(N__72222),
            .I(N__72218));
    InMux I__15355 (
            .O(N__72221),
            .I(N__72215));
    LocalMux I__15354 (
            .O(N__72218),
            .I(N__72212));
    LocalMux I__15353 (
            .O(N__72215),
            .I(data_out_frame_6_1));
    Odrv12 I__15352 (
            .O(N__72212),
            .I(data_out_frame_6_1));
    CascadeMux I__15351 (
            .O(N__72207),
            .I(N__72204));
    InMux I__15350 (
            .O(N__72204),
            .I(N__72198));
    InMux I__15349 (
            .O(N__72203),
            .I(N__72194));
    InMux I__15348 (
            .O(N__72202),
            .I(N__72189));
    InMux I__15347 (
            .O(N__72201),
            .I(N__72189));
    LocalMux I__15346 (
            .O(N__72198),
            .I(N__72185));
    InMux I__15345 (
            .O(N__72197),
            .I(N__72182));
    LocalMux I__15344 (
            .O(N__72194),
            .I(N__72177));
    LocalMux I__15343 (
            .O(N__72189),
            .I(N__72177));
    InMux I__15342 (
            .O(N__72188),
            .I(N__72174));
    Span4Mux_h I__15341 (
            .O(N__72185),
            .I(N__72171));
    LocalMux I__15340 (
            .O(N__72182),
            .I(N__72166));
    Span4Mux_v I__15339 (
            .O(N__72177),
            .I(N__72166));
    LocalMux I__15338 (
            .O(N__72174),
            .I(control_mode_2));
    Odrv4 I__15337 (
            .O(N__72171),
            .I(control_mode_2));
    Odrv4 I__15336 (
            .O(N__72166),
            .I(control_mode_2));
    InMux I__15335 (
            .O(N__72159),
            .I(N__72155));
    CascadeMux I__15334 (
            .O(N__72158),
            .I(N__72149));
    LocalMux I__15333 (
            .O(N__72155),
            .I(N__72145));
    InMux I__15332 (
            .O(N__72154),
            .I(N__72138));
    InMux I__15331 (
            .O(N__72153),
            .I(N__72138));
    InMux I__15330 (
            .O(N__72152),
            .I(N__72138));
    InMux I__15329 (
            .O(N__72149),
            .I(N__72135));
    InMux I__15328 (
            .O(N__72148),
            .I(N__72132));
    Span4Mux_h I__15327 (
            .O(N__72145),
            .I(N__72129));
    LocalMux I__15326 (
            .O(N__72138),
            .I(N__72126));
    LocalMux I__15325 (
            .O(N__72135),
            .I(control_mode_3));
    LocalMux I__15324 (
            .O(N__72132),
            .I(control_mode_3));
    Odrv4 I__15323 (
            .O(N__72129),
            .I(control_mode_3));
    Odrv12 I__15322 (
            .O(N__72126),
            .I(control_mode_3));
    CascadeMux I__15321 (
            .O(N__72117),
            .I(\c0.n30_cascade_ ));
    InMux I__15320 (
            .O(N__72114),
            .I(N__72111));
    LocalMux I__15319 (
            .O(N__72111),
            .I(\c0.n39_adj_4567 ));
    InMux I__15318 (
            .O(N__72108),
            .I(N__72105));
    LocalMux I__15317 (
            .O(N__72105),
            .I(\c0.n45_adj_4572 ));
    CascadeMux I__15316 (
            .O(N__72102),
            .I(\c0.n33314_cascade_ ));
    InMux I__15315 (
            .O(N__72099),
            .I(N__72095));
    InMux I__15314 (
            .O(N__72098),
            .I(N__72092));
    LocalMux I__15313 (
            .O(N__72095),
            .I(N__72087));
    LocalMux I__15312 (
            .O(N__72092),
            .I(N__72087));
    Span4Mux_h I__15311 (
            .O(N__72087),
            .I(N__72084));
    Odrv4 I__15310 (
            .O(N__72084),
            .I(\c0.n18124 ));
    CascadeMux I__15309 (
            .O(N__72081),
            .I(\c0.n24_cascade_ ));
    CascadeMux I__15308 (
            .O(N__72078),
            .I(N__72074));
    CascadeMux I__15307 (
            .O(N__72077),
            .I(N__72070));
    InMux I__15306 (
            .O(N__72074),
            .I(N__72066));
    InMux I__15305 (
            .O(N__72073),
            .I(N__72063));
    InMux I__15304 (
            .O(N__72070),
            .I(N__72059));
    InMux I__15303 (
            .O(N__72069),
            .I(N__72056));
    LocalMux I__15302 (
            .O(N__72066),
            .I(N__72053));
    LocalMux I__15301 (
            .O(N__72063),
            .I(N__72050));
    InMux I__15300 (
            .O(N__72062),
            .I(N__72047));
    LocalMux I__15299 (
            .O(N__72059),
            .I(N__72043));
    LocalMux I__15298 (
            .O(N__72056),
            .I(N__72040));
    Span4Mux_v I__15297 (
            .O(N__72053),
            .I(N__72033));
    Span4Mux_h I__15296 (
            .O(N__72050),
            .I(N__72033));
    LocalMux I__15295 (
            .O(N__72047),
            .I(N__72033));
    InMux I__15294 (
            .O(N__72046),
            .I(N__72030));
    Span12Mux_v I__15293 (
            .O(N__72043),
            .I(N__72027));
    Span4Mux_h I__15292 (
            .O(N__72040),
            .I(N__72022));
    Span4Mux_h I__15291 (
            .O(N__72033),
            .I(N__72022));
    LocalMux I__15290 (
            .O(N__72030),
            .I(encoder0_position_19));
    Odrv12 I__15289 (
            .O(N__72027),
            .I(encoder0_position_19));
    Odrv4 I__15288 (
            .O(N__72022),
            .I(encoder0_position_19));
    InMux I__15287 (
            .O(N__72015),
            .I(N__72012));
    LocalMux I__15286 (
            .O(N__72012),
            .I(\c0.n18 ));
    InMux I__15285 (
            .O(N__72009),
            .I(N__72005));
    CascadeMux I__15284 (
            .O(N__72008),
            .I(N__71998));
    LocalMux I__15283 (
            .O(N__72005),
            .I(N__71995));
    CascadeMux I__15282 (
            .O(N__72004),
            .I(N__71992));
    InMux I__15281 (
            .O(N__72003),
            .I(N__71989));
    InMux I__15280 (
            .O(N__72002),
            .I(N__71984));
    InMux I__15279 (
            .O(N__72001),
            .I(N__71984));
    InMux I__15278 (
            .O(N__71998),
            .I(N__71980));
    Span4Mux_h I__15277 (
            .O(N__71995),
            .I(N__71977));
    InMux I__15276 (
            .O(N__71992),
            .I(N__71974));
    LocalMux I__15275 (
            .O(N__71989),
            .I(N__71971));
    LocalMux I__15274 (
            .O(N__71984),
            .I(N__71968));
    InMux I__15273 (
            .O(N__71983),
            .I(N__71965));
    LocalMux I__15272 (
            .O(N__71980),
            .I(N__71960));
    Span4Mux_v I__15271 (
            .O(N__71977),
            .I(N__71960));
    LocalMux I__15270 (
            .O(N__71974),
            .I(N__71955));
    Span4Mux_h I__15269 (
            .O(N__71971),
            .I(N__71955));
    Span4Mux_h I__15268 (
            .O(N__71968),
            .I(N__71952));
    LocalMux I__15267 (
            .O(N__71965),
            .I(encoder0_position_20));
    Odrv4 I__15266 (
            .O(N__71960),
            .I(encoder0_position_20));
    Odrv4 I__15265 (
            .O(N__71955),
            .I(encoder0_position_20));
    Odrv4 I__15264 (
            .O(N__71952),
            .I(encoder0_position_20));
    InMux I__15263 (
            .O(N__71943),
            .I(N__71940));
    LocalMux I__15262 (
            .O(N__71940),
            .I(\c0.n33765 ));
    CascadeMux I__15261 (
            .O(N__71937),
            .I(\c0.n33765_cascade_ ));
    InMux I__15260 (
            .O(N__71934),
            .I(N__71931));
    LocalMux I__15259 (
            .O(N__71931),
            .I(\c0.n26_adj_4559 ));
    InMux I__15258 (
            .O(N__71928),
            .I(N__71925));
    LocalMux I__15257 (
            .O(N__71925),
            .I(N__71922));
    Odrv4 I__15256 (
            .O(N__71922),
            .I(\c0.n33493 ));
    InMux I__15255 (
            .O(N__71919),
            .I(N__71915));
    InMux I__15254 (
            .O(N__71918),
            .I(N__71912));
    LocalMux I__15253 (
            .O(N__71915),
            .I(N__71909));
    LocalMux I__15252 (
            .O(N__71912),
            .I(N__71904));
    Span4Mux_v I__15251 (
            .O(N__71909),
            .I(N__71904));
    Odrv4 I__15250 (
            .O(N__71904),
            .I(data_out_frame_7_7));
    InMux I__15249 (
            .O(N__71901),
            .I(N__71898));
    LocalMux I__15248 (
            .O(N__71898),
            .I(N__71895));
    Odrv12 I__15247 (
            .O(N__71895),
            .I(\c0.n5_adj_4653 ));
    InMux I__15246 (
            .O(N__71892),
            .I(N__71886));
    InMux I__15245 (
            .O(N__71891),
            .I(N__71883));
    InMux I__15244 (
            .O(N__71890),
            .I(N__71880));
    InMux I__15243 (
            .O(N__71889),
            .I(N__71877));
    LocalMux I__15242 (
            .O(N__71886),
            .I(N__71872));
    LocalMux I__15241 (
            .O(N__71883),
            .I(N__71872));
    LocalMux I__15240 (
            .O(N__71880),
            .I(N__71868));
    LocalMux I__15239 (
            .O(N__71877),
            .I(N__71863));
    Span4Mux_h I__15238 (
            .O(N__71872),
            .I(N__71863));
    InMux I__15237 (
            .O(N__71871),
            .I(N__71860));
    Odrv4 I__15236 (
            .O(N__71868),
            .I(encoder1_position_22));
    Odrv4 I__15235 (
            .O(N__71863),
            .I(encoder1_position_22));
    LocalMux I__15234 (
            .O(N__71860),
            .I(encoder1_position_22));
    InMux I__15233 (
            .O(N__71853),
            .I(N__71849));
    InMux I__15232 (
            .O(N__71852),
            .I(N__71846));
    LocalMux I__15231 (
            .O(N__71849),
            .I(data_out_frame_5_7));
    LocalMux I__15230 (
            .O(N__71846),
            .I(data_out_frame_5_7));
    InMux I__15229 (
            .O(N__71841),
            .I(N__71837));
    InMux I__15228 (
            .O(N__71840),
            .I(N__71834));
    LocalMux I__15227 (
            .O(N__71837),
            .I(data_out_frame_5_1));
    LocalMux I__15226 (
            .O(N__71834),
            .I(data_out_frame_5_1));
    InMux I__15225 (
            .O(N__71829),
            .I(N__71826));
    LocalMux I__15224 (
            .O(N__71826),
            .I(N__71823));
    Span4Mux_h I__15223 (
            .O(N__71823),
            .I(N__71820));
    Odrv4 I__15222 (
            .O(N__71820),
            .I(\c0.n36090 ));
    InMux I__15221 (
            .O(N__71817),
            .I(N__71811));
    InMux I__15220 (
            .O(N__71816),
            .I(N__71811));
    LocalMux I__15219 (
            .O(N__71811),
            .I(data_out_frame_6_7));
    CascadeMux I__15218 (
            .O(N__71808),
            .I(N__71805));
    InMux I__15217 (
            .O(N__71805),
            .I(N__71801));
    CascadeMux I__15216 (
            .O(N__71804),
            .I(N__71797));
    LocalMux I__15215 (
            .O(N__71801),
            .I(N__71794));
    InMux I__15214 (
            .O(N__71800),
            .I(N__71791));
    InMux I__15213 (
            .O(N__71797),
            .I(N__71787));
    Span4Mux_h I__15212 (
            .O(N__71794),
            .I(N__71782));
    LocalMux I__15211 (
            .O(N__71791),
            .I(N__71782));
    InMux I__15210 (
            .O(N__71790),
            .I(N__71779));
    LocalMux I__15209 (
            .O(N__71787),
            .I(N__71774));
    Span4Mux_v I__15208 (
            .O(N__71782),
            .I(N__71774));
    LocalMux I__15207 (
            .O(N__71779),
            .I(encoder0_position_1));
    Odrv4 I__15206 (
            .O(N__71774),
            .I(encoder0_position_1));
    CascadeMux I__15205 (
            .O(N__71769),
            .I(\c0.n33503_cascade_ ));
    InMux I__15204 (
            .O(N__71766),
            .I(N__71763));
    LocalMux I__15203 (
            .O(N__71763),
            .I(\c0.n47 ));
    CascadeMux I__15202 (
            .O(N__71760),
            .I(\c0.n41_adj_4571_cascade_ ));
    InMux I__15201 (
            .O(N__71757),
            .I(N__71753));
    InMux I__15200 (
            .O(N__71756),
            .I(N__71750));
    LocalMux I__15199 (
            .O(N__71753),
            .I(data_out_frame_10_5));
    LocalMux I__15198 (
            .O(N__71750),
            .I(data_out_frame_10_5));
    CascadeMux I__15197 (
            .O(N__71745),
            .I(\c0.n36016_cascade_ ));
    CascadeMux I__15196 (
            .O(N__71742),
            .I(\c0.n35827_cascade_ ));
    InMux I__15195 (
            .O(N__71739),
            .I(N__71736));
    LocalMux I__15194 (
            .O(N__71736),
            .I(N__71733));
    Span4Mux_h I__15193 (
            .O(N__71733),
            .I(N__71730));
    Odrv4 I__15192 (
            .O(N__71730),
            .I(n35829));
    InMux I__15191 (
            .O(N__71727),
            .I(N__71724));
    LocalMux I__15190 (
            .O(N__71724),
            .I(N__71721));
    Odrv4 I__15189 (
            .O(N__71721),
            .I(n2271));
    InMux I__15188 (
            .O(N__71718),
            .I(N__71714));
    InMux I__15187 (
            .O(N__71717),
            .I(N__71711));
    LocalMux I__15186 (
            .O(N__71714),
            .I(N__71708));
    LocalMux I__15185 (
            .O(N__71711),
            .I(data_out_frame_5_0));
    Odrv4 I__15184 (
            .O(N__71708),
            .I(data_out_frame_5_0));
    InMux I__15183 (
            .O(N__71703),
            .I(N__71700));
    LocalMux I__15182 (
            .O(N__71700),
            .I(N__71697));
    Odrv4 I__15181 (
            .O(N__71697),
            .I(n2259));
    InMux I__15180 (
            .O(N__71694),
            .I(N__71691));
    LocalMux I__15179 (
            .O(N__71691),
            .I(N__71685));
    InMux I__15178 (
            .O(N__71690),
            .I(N__71682));
    InMux I__15177 (
            .O(N__71689),
            .I(N__71677));
    InMux I__15176 (
            .O(N__71688),
            .I(N__71677));
    Span4Mux_v I__15175 (
            .O(N__71685),
            .I(N__71673));
    LocalMux I__15174 (
            .O(N__71682),
            .I(N__71670));
    LocalMux I__15173 (
            .O(N__71677),
            .I(N__71667));
    InMux I__15172 (
            .O(N__71676),
            .I(N__71663));
    Span4Mux_h I__15171 (
            .O(N__71673),
            .I(N__71655));
    Span4Mux_v I__15170 (
            .O(N__71670),
            .I(N__71655));
    Span4Mux_v I__15169 (
            .O(N__71667),
            .I(N__71655));
    InMux I__15168 (
            .O(N__71666),
            .I(N__71652));
    LocalMux I__15167 (
            .O(N__71663),
            .I(N__71648));
    InMux I__15166 (
            .O(N__71662),
            .I(N__71645));
    Span4Mux_h I__15165 (
            .O(N__71655),
            .I(N__71640));
    LocalMux I__15164 (
            .O(N__71652),
            .I(N__71640));
    InMux I__15163 (
            .O(N__71651),
            .I(N__71637));
    Span4Mux_h I__15162 (
            .O(N__71648),
            .I(N__71634));
    LocalMux I__15161 (
            .O(N__71645),
            .I(N__71631));
    Span4Mux_h I__15160 (
            .O(N__71640),
            .I(N__71628));
    LocalMux I__15159 (
            .O(N__71637),
            .I(N__71625));
    Odrv4 I__15158 (
            .O(N__71634),
            .I(n14821));
    Odrv12 I__15157 (
            .O(N__71631),
            .I(n14821));
    Odrv4 I__15156 (
            .O(N__71628),
            .I(n14821));
    Odrv12 I__15155 (
            .O(N__71625),
            .I(n14821));
    InMux I__15154 (
            .O(N__71616),
            .I(N__71613));
    LocalMux I__15153 (
            .O(N__71613),
            .I(N__71610));
    Span4Mux_v I__15152 (
            .O(N__71610),
            .I(N__71606));
    InMux I__15151 (
            .O(N__71609),
            .I(N__71603));
    Sp12to4 I__15150 (
            .O(N__71606),
            .I(N__71600));
    LocalMux I__15149 (
            .O(N__71603),
            .I(r_Tx_Data_5));
    Odrv12 I__15148 (
            .O(N__71600),
            .I(r_Tx_Data_5));
    InMux I__15147 (
            .O(N__71595),
            .I(N__71592));
    LocalMux I__15146 (
            .O(N__71592),
            .I(N__71589));
    Odrv4 I__15145 (
            .O(N__71589),
            .I(\quad_counter1.n35603 ));
    InMux I__15144 (
            .O(N__71586),
            .I(N__71583));
    LocalMux I__15143 (
            .O(N__71583),
            .I(N__71580));
    Span4Mux_h I__15142 (
            .O(N__71580),
            .I(N__71577));
    Span4Mux_v I__15141 (
            .O(N__71577),
            .I(N__71574));
    Odrv4 I__15140 (
            .O(N__71574),
            .I(\c0.n35824 ));
    CascadeMux I__15139 (
            .O(N__71571),
            .I(\c0.n26_adj_4625_cascade_ ));
    CascadeMux I__15138 (
            .O(N__71568),
            .I(N__71565));
    InMux I__15137 (
            .O(N__71565),
            .I(N__71562));
    LocalMux I__15136 (
            .O(N__71562),
            .I(N__71559));
    Sp12to4 I__15135 (
            .O(N__71559),
            .I(N__71556));
    Span12Mux_v I__15134 (
            .O(N__71556),
            .I(N__71553));
    Odrv12 I__15133 (
            .O(N__71553),
            .I(n35826));
    InMux I__15132 (
            .O(N__71550),
            .I(N__71547));
    LocalMux I__15131 (
            .O(N__71547),
            .I(N__71544));
    Odrv4 I__15130 (
            .O(N__71544),
            .I(n2274));
    CascadeMux I__15129 (
            .O(N__71541),
            .I(N__71538));
    InMux I__15128 (
            .O(N__71538),
            .I(N__71532));
    InMux I__15127 (
            .O(N__71537),
            .I(N__71532));
    LocalMux I__15126 (
            .O(N__71532),
            .I(data_out_frame_7_1));
    CascadeMux I__15125 (
            .O(N__71529),
            .I(\c0.n5_adj_4505_cascade_ ));
    CascadeMux I__15124 (
            .O(N__71526),
            .I(\c0.n35830_cascade_ ));
    CascadeMux I__15123 (
            .O(N__71523),
            .I(N__71520));
    InMux I__15122 (
            .O(N__71520),
            .I(N__71517));
    LocalMux I__15121 (
            .O(N__71517),
            .I(N__71514));
    Span4Mux_h I__15120 (
            .O(N__71514),
            .I(N__71511));
    Span4Mux_h I__15119 (
            .O(N__71511),
            .I(N__71508));
    Odrv4 I__15118 (
            .O(N__71508),
            .I(n35832));
    InMux I__15117 (
            .O(N__71505),
            .I(N__71485));
    InMux I__15116 (
            .O(N__71504),
            .I(N__71482));
    InMux I__15115 (
            .O(N__71503),
            .I(N__71479));
    InMux I__15114 (
            .O(N__71502),
            .I(N__71476));
    InMux I__15113 (
            .O(N__71501),
            .I(N__71469));
    InMux I__15112 (
            .O(N__71500),
            .I(N__71466));
    InMux I__15111 (
            .O(N__71499),
            .I(N__71463));
    InMux I__15110 (
            .O(N__71498),
            .I(N__71460));
    InMux I__15109 (
            .O(N__71497),
            .I(N__71457));
    InMux I__15108 (
            .O(N__71496),
            .I(N__71454));
    InMux I__15107 (
            .O(N__71495),
            .I(N__71451));
    InMux I__15106 (
            .O(N__71494),
            .I(N__71448));
    InMux I__15105 (
            .O(N__71493),
            .I(N__71441));
    InMux I__15104 (
            .O(N__71492),
            .I(N__71438));
    InMux I__15103 (
            .O(N__71491),
            .I(N__71435));
    InMux I__15102 (
            .O(N__71490),
            .I(N__71432));
    InMux I__15101 (
            .O(N__71489),
            .I(N__71429));
    InMux I__15100 (
            .O(N__71488),
            .I(N__71426));
    LocalMux I__15099 (
            .O(N__71485),
            .I(N__71417));
    LocalMux I__15098 (
            .O(N__71482),
            .I(N__71417));
    LocalMux I__15097 (
            .O(N__71479),
            .I(N__71417));
    LocalMux I__15096 (
            .O(N__71476),
            .I(N__71417));
    InMux I__15095 (
            .O(N__71475),
            .I(N__71414));
    InMux I__15094 (
            .O(N__71474),
            .I(N__71411));
    InMux I__15093 (
            .O(N__71473),
            .I(N__71407));
    InMux I__15092 (
            .O(N__71472),
            .I(N__71404));
    LocalMux I__15091 (
            .O(N__71469),
            .I(N__71401));
    LocalMux I__15090 (
            .O(N__71466),
            .I(N__71394));
    LocalMux I__15089 (
            .O(N__71463),
            .I(N__71394));
    LocalMux I__15088 (
            .O(N__71460),
            .I(N__71394));
    LocalMux I__15087 (
            .O(N__71457),
            .I(N__71385));
    LocalMux I__15086 (
            .O(N__71454),
            .I(N__71385));
    LocalMux I__15085 (
            .O(N__71451),
            .I(N__71385));
    LocalMux I__15084 (
            .O(N__71448),
            .I(N__71385));
    InMux I__15083 (
            .O(N__71447),
            .I(N__71382));
    InMux I__15082 (
            .O(N__71446),
            .I(N__71379));
    InMux I__15081 (
            .O(N__71445),
            .I(N__71376));
    InMux I__15080 (
            .O(N__71444),
            .I(N__71373));
    LocalMux I__15079 (
            .O(N__71441),
            .I(N__71368));
    LocalMux I__15078 (
            .O(N__71438),
            .I(N__71368));
    LocalMux I__15077 (
            .O(N__71435),
            .I(N__71363));
    LocalMux I__15076 (
            .O(N__71432),
            .I(N__71363));
    LocalMux I__15075 (
            .O(N__71429),
            .I(N__71356));
    LocalMux I__15074 (
            .O(N__71426),
            .I(N__71356));
    Span4Mux_v I__15073 (
            .O(N__71417),
            .I(N__71356));
    LocalMux I__15072 (
            .O(N__71414),
            .I(N__71351));
    LocalMux I__15071 (
            .O(N__71411),
            .I(N__71351));
    InMux I__15070 (
            .O(N__71410),
            .I(N__71348));
    LocalMux I__15069 (
            .O(N__71407),
            .I(N__71337));
    LocalMux I__15068 (
            .O(N__71404),
            .I(N__71337));
    Span4Mux_v I__15067 (
            .O(N__71401),
            .I(N__71337));
    Span4Mux_v I__15066 (
            .O(N__71394),
            .I(N__71337));
    Span4Mux_v I__15065 (
            .O(N__71385),
            .I(N__71337));
    LocalMux I__15064 (
            .O(N__71382),
            .I(N__71332));
    LocalMux I__15063 (
            .O(N__71379),
            .I(N__71332));
    LocalMux I__15062 (
            .O(N__71376),
            .I(N__71323));
    LocalMux I__15061 (
            .O(N__71373),
            .I(N__71323));
    Span4Mux_v I__15060 (
            .O(N__71368),
            .I(N__71323));
    Span4Mux_v I__15059 (
            .O(N__71363),
            .I(N__71323));
    Span4Mux_v I__15058 (
            .O(N__71356),
            .I(N__71317));
    Span4Mux_v I__15057 (
            .O(N__71351),
            .I(N__71317));
    LocalMux I__15056 (
            .O(N__71348),
            .I(N__71313));
    Sp12to4 I__15055 (
            .O(N__71337),
            .I(N__71310));
    Span4Mux_v I__15054 (
            .O(N__71332),
            .I(N__71305));
    Span4Mux_h I__15053 (
            .O(N__71323),
            .I(N__71305));
    InMux I__15052 (
            .O(N__71322),
            .I(N__71302));
    Span4Mux_h I__15051 (
            .O(N__71317),
            .I(N__71299));
    InMux I__15050 (
            .O(N__71316),
            .I(N__71296));
    Span12Mux_h I__15049 (
            .O(N__71313),
            .I(N__71293));
    Span12Mux_s8_h I__15048 (
            .O(N__71310),
            .I(N__71290));
    Span4Mux_h I__15047 (
            .O(N__71305),
            .I(N__71287));
    LocalMux I__15046 (
            .O(N__71302),
            .I(N__71282));
    Span4Mux_h I__15045 (
            .O(N__71299),
            .I(N__71282));
    LocalMux I__15044 (
            .O(N__71296),
            .I(\c0.n4_adj_4623 ));
    Odrv12 I__15043 (
            .O(N__71293),
            .I(\c0.n4_adj_4623 ));
    Odrv12 I__15042 (
            .O(N__71290),
            .I(\c0.n4_adj_4623 ));
    Odrv4 I__15041 (
            .O(N__71287),
            .I(\c0.n4_adj_4623 ));
    Odrv4 I__15040 (
            .O(N__71282),
            .I(\c0.n4_adj_4623 ));
    CascadeMux I__15039 (
            .O(N__71271),
            .I(N__71267));
    InMux I__15038 (
            .O(N__71270),
            .I(N__71264));
    InMux I__15037 (
            .O(N__71267),
            .I(N__71259));
    LocalMux I__15036 (
            .O(N__71264),
            .I(N__71256));
    InMux I__15035 (
            .O(N__71263),
            .I(N__71251));
    InMux I__15034 (
            .O(N__71262),
            .I(N__71251));
    LocalMux I__15033 (
            .O(N__71259),
            .I(N__71248));
    Span4Mux_v I__15032 (
            .O(N__71256),
            .I(N__71245));
    LocalMux I__15031 (
            .O(N__71251),
            .I(N__71242));
    Span4Mux_v I__15030 (
            .O(N__71248),
            .I(N__71239));
    Span4Mux_h I__15029 (
            .O(N__71245),
            .I(N__71234));
    Span4Mux_v I__15028 (
            .O(N__71242),
            .I(N__71234));
    Span4Mux_h I__15027 (
            .O(N__71239),
            .I(N__71230));
    Span4Mux_h I__15026 (
            .O(N__71234),
            .I(N__71227));
    InMux I__15025 (
            .O(N__71233),
            .I(N__71224));
    Span4Mux_h I__15024 (
            .O(N__71230),
            .I(N__71221));
    Span4Mux_h I__15023 (
            .O(N__71227),
            .I(N__71218));
    LocalMux I__15022 (
            .O(N__71224),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__15021 (
            .O(N__71221),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__15020 (
            .O(N__71218),
            .I(\c0.FRAME_MATCHER_state_3 ));
    SRMux I__15019 (
            .O(N__71211),
            .I(N__71208));
    LocalMux I__15018 (
            .O(N__71208),
            .I(N__71205));
    Sp12to4 I__15017 (
            .O(N__71205),
            .I(N__71202));
    Span12Mux_v I__15016 (
            .O(N__71202),
            .I(N__71199));
    Odrv12 I__15015 (
            .O(N__71199),
            .I(\c0.n32750 ));
    InMux I__15014 (
            .O(N__71196),
            .I(N__71193));
    LocalMux I__15013 (
            .O(N__71193),
            .I(\quad_counter1.n8 ));
    InMux I__15012 (
            .O(N__71190),
            .I(N__71187));
    LocalMux I__15011 (
            .O(N__71187),
            .I(\quad_counter1.n8_adj_4444 ));
    CascadeMux I__15010 (
            .O(N__71184),
            .I(\quad_counter1.n35309_cascade_ ));
    CascadeMux I__15009 (
            .O(N__71181),
            .I(N__71178));
    InMux I__15008 (
            .O(N__71178),
            .I(N__71175));
    LocalMux I__15007 (
            .O(N__71175),
            .I(\quad_counter1.n7 ));
    InMux I__15006 (
            .O(N__71172),
            .I(N__71169));
    LocalMux I__15005 (
            .O(N__71169),
            .I(N__71166));
    Odrv4 I__15004 (
            .O(N__71166),
            .I(n10_adj_4821));
    CascadeMux I__15003 (
            .O(N__71163),
            .I(N__71160));
    InMux I__15002 (
            .O(N__71160),
            .I(N__71156));
    CascadeMux I__15001 (
            .O(N__71159),
            .I(N__71151));
    LocalMux I__15000 (
            .O(N__71156),
            .I(N__71148));
    CascadeMux I__14999 (
            .O(N__71155),
            .I(N__71143));
    InMux I__14998 (
            .O(N__71154),
            .I(N__71140));
    InMux I__14997 (
            .O(N__71151),
            .I(N__71137));
    Span4Mux_v I__14996 (
            .O(N__71148),
            .I(N__71134));
    CascadeMux I__14995 (
            .O(N__71147),
            .I(N__71131));
    CascadeMux I__14994 (
            .O(N__71146),
            .I(N__71128));
    InMux I__14993 (
            .O(N__71143),
            .I(N__71125));
    LocalMux I__14992 (
            .O(N__71140),
            .I(N__71121));
    LocalMux I__14991 (
            .O(N__71137),
            .I(N__71118));
    Span4Mux_h I__14990 (
            .O(N__71134),
            .I(N__71115));
    InMux I__14989 (
            .O(N__71131),
            .I(N__71109));
    InMux I__14988 (
            .O(N__71128),
            .I(N__71106));
    LocalMux I__14987 (
            .O(N__71125),
            .I(N__71103));
    InMux I__14986 (
            .O(N__71124),
            .I(N__71100));
    Span4Mux_h I__14985 (
            .O(N__71121),
            .I(N__71097));
    Span4Mux_h I__14984 (
            .O(N__71118),
            .I(N__71092));
    Span4Mux_h I__14983 (
            .O(N__71115),
            .I(N__71092));
    InMux I__14982 (
            .O(N__71114),
            .I(N__71085));
    InMux I__14981 (
            .O(N__71113),
            .I(N__71085));
    InMux I__14980 (
            .O(N__71112),
            .I(N__71085));
    LocalMux I__14979 (
            .O(N__71109),
            .I(byte_transmit_counter_5));
    LocalMux I__14978 (
            .O(N__71106),
            .I(byte_transmit_counter_5));
    Odrv12 I__14977 (
            .O(N__71103),
            .I(byte_transmit_counter_5));
    LocalMux I__14976 (
            .O(N__71100),
            .I(byte_transmit_counter_5));
    Odrv4 I__14975 (
            .O(N__71097),
            .I(byte_transmit_counter_5));
    Odrv4 I__14974 (
            .O(N__71092),
            .I(byte_transmit_counter_5));
    LocalMux I__14973 (
            .O(N__71085),
            .I(byte_transmit_counter_5));
    InMux I__14972 (
            .O(N__71070),
            .I(N__71066));
    InMux I__14971 (
            .O(N__71069),
            .I(N__71063));
    LocalMux I__14970 (
            .O(N__71066),
            .I(N__71057));
    LocalMux I__14969 (
            .O(N__71063),
            .I(N__71057));
    InMux I__14968 (
            .O(N__71062),
            .I(N__71054));
    Odrv4 I__14967 (
            .O(N__71057),
            .I(\quad_counter1.n3105 ));
    LocalMux I__14966 (
            .O(N__71054),
            .I(\quad_counter1.n3105 ));
    InMux I__14965 (
            .O(N__71049),
            .I(N__71045));
    InMux I__14964 (
            .O(N__71048),
            .I(N__71042));
    LocalMux I__14963 (
            .O(N__71045),
            .I(N__71036));
    LocalMux I__14962 (
            .O(N__71042),
            .I(N__71036));
    CascadeMux I__14961 (
            .O(N__71041),
            .I(N__71033));
    Span4Mux_v I__14960 (
            .O(N__71036),
            .I(N__71030));
    InMux I__14959 (
            .O(N__71033),
            .I(N__71027));
    Odrv4 I__14958 (
            .O(N__71030),
            .I(\quad_counter1.n3204 ));
    LocalMux I__14957 (
            .O(N__71027),
            .I(\quad_counter1.n3204 ));
    InMux I__14956 (
            .O(N__71022),
            .I(\quad_counter1.n30629 ));
    InMux I__14955 (
            .O(N__71019),
            .I(N__71016));
    LocalMux I__14954 (
            .O(N__71016),
            .I(N__71012));
    InMux I__14953 (
            .O(N__71015),
            .I(N__71009));
    Span4Mux_h I__14952 (
            .O(N__71012),
            .I(N__71004));
    LocalMux I__14951 (
            .O(N__71009),
            .I(N__71004));
    Span4Mux_v I__14950 (
            .O(N__71004),
            .I(N__71000));
    InMux I__14949 (
            .O(N__71003),
            .I(N__70997));
    Odrv4 I__14948 (
            .O(N__71000),
            .I(\quad_counter1.n3104 ));
    LocalMux I__14947 (
            .O(N__70997),
            .I(\quad_counter1.n3104 ));
    InMux I__14946 (
            .O(N__70992),
            .I(N__70988));
    InMux I__14945 (
            .O(N__70991),
            .I(N__70985));
    LocalMux I__14944 (
            .O(N__70988),
            .I(N__70980));
    LocalMux I__14943 (
            .O(N__70985),
            .I(N__70980));
    Span4Mux_v I__14942 (
            .O(N__70980),
            .I(N__70976));
    InMux I__14941 (
            .O(N__70979),
            .I(N__70973));
    Odrv4 I__14940 (
            .O(N__70976),
            .I(\quad_counter1.n3203 ));
    LocalMux I__14939 (
            .O(N__70973),
            .I(\quad_counter1.n3203 ));
    InMux I__14938 (
            .O(N__70968),
            .I(bfn_20_10_0_));
    InMux I__14937 (
            .O(N__70965),
            .I(N__70962));
    LocalMux I__14936 (
            .O(N__70962),
            .I(N__70958));
    InMux I__14935 (
            .O(N__70961),
            .I(N__70955));
    Span4Mux_v I__14934 (
            .O(N__70958),
            .I(N__70952));
    LocalMux I__14933 (
            .O(N__70955),
            .I(N__70949));
    Span4Mux_h I__14932 (
            .O(N__70952),
            .I(N__70943));
    Span4Mux_v I__14931 (
            .O(N__70949),
            .I(N__70943));
    InMux I__14930 (
            .O(N__70948),
            .I(N__70940));
    Odrv4 I__14929 (
            .O(N__70943),
            .I(\quad_counter1.n3103 ));
    LocalMux I__14928 (
            .O(N__70940),
            .I(\quad_counter1.n3103 ));
    InMux I__14927 (
            .O(N__70935),
            .I(N__70930));
    InMux I__14926 (
            .O(N__70934),
            .I(N__70925));
    InMux I__14925 (
            .O(N__70933),
            .I(N__70925));
    LocalMux I__14924 (
            .O(N__70930),
            .I(N__70920));
    LocalMux I__14923 (
            .O(N__70925),
            .I(N__70920));
    Span4Mux_v I__14922 (
            .O(N__70920),
            .I(N__70917));
    Odrv4 I__14921 (
            .O(N__70917),
            .I(\quad_counter1.n3202 ));
    InMux I__14920 (
            .O(N__70914),
            .I(\quad_counter1.n30631 ));
    InMux I__14919 (
            .O(N__70911),
            .I(N__70907));
    InMux I__14918 (
            .O(N__70910),
            .I(N__70904));
    LocalMux I__14917 (
            .O(N__70907),
            .I(N__70898));
    LocalMux I__14916 (
            .O(N__70904),
            .I(N__70898));
    InMux I__14915 (
            .O(N__70903),
            .I(N__70895));
    Span4Mux_v I__14914 (
            .O(N__70898),
            .I(N__70892));
    LocalMux I__14913 (
            .O(N__70895),
            .I(N__70889));
    Odrv4 I__14912 (
            .O(N__70892),
            .I(\quad_counter1.n3102 ));
    Odrv4 I__14911 (
            .O(N__70889),
            .I(\quad_counter1.n3102 ));
    InMux I__14910 (
            .O(N__70884),
            .I(N__70880));
    InMux I__14909 (
            .O(N__70883),
            .I(N__70877));
    LocalMux I__14908 (
            .O(N__70880),
            .I(N__70872));
    LocalMux I__14907 (
            .O(N__70877),
            .I(N__70872));
    Span4Mux_h I__14906 (
            .O(N__70872),
            .I(N__70868));
    InMux I__14905 (
            .O(N__70871),
            .I(N__70865));
    Odrv4 I__14904 (
            .O(N__70868),
            .I(\quad_counter1.n3201 ));
    LocalMux I__14903 (
            .O(N__70865),
            .I(\quad_counter1.n3201 ));
    InMux I__14902 (
            .O(N__70860),
            .I(\quad_counter1.n30632 ));
    InMux I__14901 (
            .O(N__70857),
            .I(N__70853));
    InMux I__14900 (
            .O(N__70856),
            .I(N__70850));
    LocalMux I__14899 (
            .O(N__70853),
            .I(N__70844));
    LocalMux I__14898 (
            .O(N__70850),
            .I(N__70844));
    InMux I__14897 (
            .O(N__70849),
            .I(N__70841));
    Odrv4 I__14896 (
            .O(N__70844),
            .I(\quad_counter1.n3101 ));
    LocalMux I__14895 (
            .O(N__70841),
            .I(\quad_counter1.n3101 ));
    CascadeMux I__14894 (
            .O(N__70836),
            .I(N__70830));
    CascadeMux I__14893 (
            .O(N__70835),
            .I(N__70827));
    CascadeMux I__14892 (
            .O(N__70834),
            .I(N__70824));
    CascadeMux I__14891 (
            .O(N__70833),
            .I(N__70821));
    InMux I__14890 (
            .O(N__70830),
            .I(N__70808));
    InMux I__14889 (
            .O(N__70827),
            .I(N__70808));
    InMux I__14888 (
            .O(N__70824),
            .I(N__70803));
    InMux I__14887 (
            .O(N__70821),
            .I(N__70803));
    CascadeMux I__14886 (
            .O(N__70820),
            .I(N__70800));
    CascadeMux I__14885 (
            .O(N__70819),
            .I(N__70797));
    CascadeMux I__14884 (
            .O(N__70818),
            .I(N__70794));
    CascadeMux I__14883 (
            .O(N__70817),
            .I(N__70791));
    CascadeMux I__14882 (
            .O(N__70816),
            .I(N__70788));
    CascadeMux I__14881 (
            .O(N__70815),
            .I(N__70785));
    CascadeMux I__14880 (
            .O(N__70814),
            .I(N__70782));
    CascadeMux I__14879 (
            .O(N__70813),
            .I(N__70779));
    LocalMux I__14878 (
            .O(N__70808),
            .I(N__70772));
    LocalMux I__14877 (
            .O(N__70803),
            .I(N__70772));
    InMux I__14876 (
            .O(N__70800),
            .I(N__70763));
    InMux I__14875 (
            .O(N__70797),
            .I(N__70763));
    InMux I__14874 (
            .O(N__70794),
            .I(N__70763));
    InMux I__14873 (
            .O(N__70791),
            .I(N__70763));
    InMux I__14872 (
            .O(N__70788),
            .I(N__70754));
    InMux I__14871 (
            .O(N__70785),
            .I(N__70754));
    InMux I__14870 (
            .O(N__70782),
            .I(N__70754));
    InMux I__14869 (
            .O(N__70779),
            .I(N__70754));
    CascadeMux I__14868 (
            .O(N__70778),
            .I(N__70751));
    CascadeMux I__14867 (
            .O(N__70777),
            .I(N__70748));
    Sp12to4 I__14866 (
            .O(N__70772),
            .I(N__70741));
    LocalMux I__14865 (
            .O(N__70763),
            .I(N__70741));
    LocalMux I__14864 (
            .O(N__70754),
            .I(N__70741));
    InMux I__14863 (
            .O(N__70751),
            .I(N__70736));
    InMux I__14862 (
            .O(N__70748),
            .I(N__70736));
    Odrv12 I__14861 (
            .O(N__70741),
            .I(\quad_counter1.n3134 ));
    LocalMux I__14860 (
            .O(N__70736),
            .I(\quad_counter1.n3134 ));
    InMux I__14859 (
            .O(N__70731),
            .I(\quad_counter1.n30633 ));
    InMux I__14858 (
            .O(N__70728),
            .I(N__70724));
    InMux I__14857 (
            .O(N__70727),
            .I(N__70721));
    LocalMux I__14856 (
            .O(N__70724),
            .I(N__70716));
    LocalMux I__14855 (
            .O(N__70721),
            .I(N__70716));
    Span4Mux_v I__14854 (
            .O(N__70716),
            .I(N__70712));
    InMux I__14853 (
            .O(N__70715),
            .I(N__70709));
    Odrv4 I__14852 (
            .O(N__70712),
            .I(\quad_counter1.n3200 ));
    LocalMux I__14851 (
            .O(N__70709),
            .I(\quad_counter1.n3200 ));
    CascadeMux I__14850 (
            .O(N__70704),
            .I(N__70701));
    InMux I__14849 (
            .O(N__70701),
            .I(N__70698));
    LocalMux I__14848 (
            .O(N__70698),
            .I(N__70693));
    InMux I__14847 (
            .O(N__70697),
            .I(N__70690));
    InMux I__14846 (
            .O(N__70696),
            .I(N__70687));
    Span12Mux_h I__14845 (
            .O(N__70693),
            .I(N__70684));
    LocalMux I__14844 (
            .O(N__70690),
            .I(\quad_counter0.n3117 ));
    LocalMux I__14843 (
            .O(N__70687),
            .I(\quad_counter0.n3117 ));
    Odrv12 I__14842 (
            .O(N__70684),
            .I(\quad_counter0.n3117 ));
    InMux I__14841 (
            .O(N__70677),
            .I(N__70674));
    LocalMux I__14840 (
            .O(N__70674),
            .I(N__70671));
    Span4Mux_h I__14839 (
            .O(N__70671),
            .I(N__70668));
    Span4Mux_h I__14838 (
            .O(N__70668),
            .I(N__70663));
    InMux I__14837 (
            .O(N__70667),
            .I(N__70660));
    InMux I__14836 (
            .O(N__70666),
            .I(N__70657));
    Span4Mux_h I__14835 (
            .O(N__70663),
            .I(N__70654));
    LocalMux I__14834 (
            .O(N__70660),
            .I(\quad_counter0.n3114 ));
    LocalMux I__14833 (
            .O(N__70657),
            .I(\quad_counter0.n3114 ));
    Odrv4 I__14832 (
            .O(N__70654),
            .I(\quad_counter0.n3114 ));
    InMux I__14831 (
            .O(N__70647),
            .I(N__70644));
    LocalMux I__14830 (
            .O(N__70644),
            .I(N__70641));
    Span4Mux_h I__14829 (
            .O(N__70641),
            .I(N__70638));
    Span4Mux_h I__14828 (
            .O(N__70638),
            .I(N__70635));
    Span4Mux_h I__14827 (
            .O(N__70635),
            .I(N__70632));
    Odrv4 I__14826 (
            .O(N__70632),
            .I(\quad_counter0.n8 ));
    CascadeMux I__14825 (
            .O(N__70629),
            .I(N__70624));
    InMux I__14824 (
            .O(N__70628),
            .I(N__70621));
    InMux I__14823 (
            .O(N__70627),
            .I(N__70618));
    InMux I__14822 (
            .O(N__70624),
            .I(N__70615));
    LocalMux I__14821 (
            .O(N__70621),
            .I(N__70610));
    LocalMux I__14820 (
            .O(N__70618),
            .I(N__70610));
    LocalMux I__14819 (
            .O(N__70615),
            .I(N__70607));
    Odrv12 I__14818 (
            .O(N__70610),
            .I(\quad_counter0.n2417 ));
    Odrv4 I__14817 (
            .O(N__70607),
            .I(\quad_counter0.n2417 ));
    InMux I__14816 (
            .O(N__70602),
            .I(N__70598));
    InMux I__14815 (
            .O(N__70601),
            .I(N__70595));
    LocalMux I__14814 (
            .O(N__70598),
            .I(N__70589));
    LocalMux I__14813 (
            .O(N__70595),
            .I(N__70589));
    InMux I__14812 (
            .O(N__70594),
            .I(N__70586));
    Span4Mux_v I__14811 (
            .O(N__70589),
            .I(N__70581));
    LocalMux I__14810 (
            .O(N__70586),
            .I(N__70581));
    Odrv4 I__14809 (
            .O(N__70581),
            .I(\quad_counter0.n2414 ));
    InMux I__14808 (
            .O(N__70578),
            .I(N__70575));
    LocalMux I__14807 (
            .O(N__70575),
            .I(N__70572));
    Span4Mux_h I__14806 (
            .O(N__70572),
            .I(N__70569));
    Span4Mux_h I__14805 (
            .O(N__70569),
            .I(N__70566));
    Odrv4 I__14804 (
            .O(N__70566),
            .I(\quad_counter0.n8_adj_4394 ));
    InMux I__14803 (
            .O(N__70563),
            .I(\quad_counter1.n30621 ));
    InMux I__14802 (
            .O(N__70560),
            .I(N__70556));
    InMux I__14801 (
            .O(N__70559),
            .I(N__70553));
    LocalMux I__14800 (
            .O(N__70556),
            .I(N__70547));
    LocalMux I__14799 (
            .O(N__70553),
            .I(N__70547));
    InMux I__14798 (
            .O(N__70552),
            .I(N__70544));
    Span4Mux_v I__14797 (
            .O(N__70547),
            .I(N__70539));
    LocalMux I__14796 (
            .O(N__70544),
            .I(N__70539));
    Odrv4 I__14795 (
            .O(N__70539),
            .I(\quad_counter1.n3112 ));
    InMux I__14794 (
            .O(N__70536),
            .I(N__70532));
    InMux I__14793 (
            .O(N__70535),
            .I(N__70529));
    LocalMux I__14792 (
            .O(N__70532),
            .I(N__70524));
    LocalMux I__14791 (
            .O(N__70529),
            .I(N__70524));
    Span4Mux_v I__14790 (
            .O(N__70524),
            .I(N__70520));
    InMux I__14789 (
            .O(N__70523),
            .I(N__70517));
    Odrv4 I__14788 (
            .O(N__70520),
            .I(\quad_counter1.n3211 ));
    LocalMux I__14787 (
            .O(N__70517),
            .I(\quad_counter1.n3211 ));
    InMux I__14786 (
            .O(N__70512),
            .I(bfn_20_9_0_));
    InMux I__14785 (
            .O(N__70509),
            .I(N__70505));
    InMux I__14784 (
            .O(N__70508),
            .I(N__70502));
    LocalMux I__14783 (
            .O(N__70505),
            .I(N__70497));
    LocalMux I__14782 (
            .O(N__70502),
            .I(N__70497));
    Span4Mux_v I__14781 (
            .O(N__70497),
            .I(N__70493));
    InMux I__14780 (
            .O(N__70496),
            .I(N__70490));
    Odrv4 I__14779 (
            .O(N__70493),
            .I(\quad_counter1.n3111 ));
    LocalMux I__14778 (
            .O(N__70490),
            .I(\quad_counter1.n3111 ));
    InMux I__14777 (
            .O(N__70485),
            .I(N__70481));
    InMux I__14776 (
            .O(N__70484),
            .I(N__70478));
    LocalMux I__14775 (
            .O(N__70481),
            .I(N__70472));
    LocalMux I__14774 (
            .O(N__70478),
            .I(N__70472));
    CascadeMux I__14773 (
            .O(N__70477),
            .I(N__70469));
    Span4Mux_v I__14772 (
            .O(N__70472),
            .I(N__70466));
    InMux I__14771 (
            .O(N__70469),
            .I(N__70463));
    Odrv4 I__14770 (
            .O(N__70466),
            .I(\quad_counter1.n3210 ));
    LocalMux I__14769 (
            .O(N__70463),
            .I(\quad_counter1.n3210 ));
    InMux I__14768 (
            .O(N__70458),
            .I(\quad_counter1.n30623 ));
    InMux I__14767 (
            .O(N__70455),
            .I(N__70451));
    InMux I__14766 (
            .O(N__70454),
            .I(N__70448));
    LocalMux I__14765 (
            .O(N__70451),
            .I(N__70442));
    LocalMux I__14764 (
            .O(N__70448),
            .I(N__70442));
    CascadeMux I__14763 (
            .O(N__70447),
            .I(N__70439));
    Span4Mux_v I__14762 (
            .O(N__70442),
            .I(N__70436));
    InMux I__14761 (
            .O(N__70439),
            .I(N__70433));
    Odrv4 I__14760 (
            .O(N__70436),
            .I(\quad_counter1.n3110 ));
    LocalMux I__14759 (
            .O(N__70433),
            .I(\quad_counter1.n3110 ));
    InMux I__14758 (
            .O(N__70428),
            .I(N__70425));
    LocalMux I__14757 (
            .O(N__70425),
            .I(N__70421));
    InMux I__14756 (
            .O(N__70424),
            .I(N__70418));
    Span4Mux_h I__14755 (
            .O(N__70421),
            .I(N__70412));
    LocalMux I__14754 (
            .O(N__70418),
            .I(N__70412));
    InMux I__14753 (
            .O(N__70417),
            .I(N__70409));
    Odrv4 I__14752 (
            .O(N__70412),
            .I(\quad_counter1.n3209 ));
    LocalMux I__14751 (
            .O(N__70409),
            .I(\quad_counter1.n3209 ));
    InMux I__14750 (
            .O(N__70404),
            .I(\quad_counter1.n30624 ));
    InMux I__14749 (
            .O(N__70401),
            .I(N__70397));
    InMux I__14748 (
            .O(N__70400),
            .I(N__70394));
    LocalMux I__14747 (
            .O(N__70397),
            .I(N__70388));
    LocalMux I__14746 (
            .O(N__70394),
            .I(N__70388));
    CascadeMux I__14745 (
            .O(N__70393),
            .I(N__70385));
    Span4Mux_v I__14744 (
            .O(N__70388),
            .I(N__70382));
    InMux I__14743 (
            .O(N__70385),
            .I(N__70379));
    Odrv4 I__14742 (
            .O(N__70382),
            .I(\quad_counter1.n3109 ));
    LocalMux I__14741 (
            .O(N__70379),
            .I(\quad_counter1.n3109 ));
    InMux I__14740 (
            .O(N__70374),
            .I(N__70370));
    InMux I__14739 (
            .O(N__70373),
            .I(N__70367));
    LocalMux I__14738 (
            .O(N__70370),
            .I(N__70364));
    LocalMux I__14737 (
            .O(N__70367),
            .I(N__70358));
    Span4Mux_h I__14736 (
            .O(N__70364),
            .I(N__70358));
    InMux I__14735 (
            .O(N__70363),
            .I(N__70355));
    Odrv4 I__14734 (
            .O(N__70358),
            .I(\quad_counter1.n3208 ));
    LocalMux I__14733 (
            .O(N__70355),
            .I(\quad_counter1.n3208 ));
    InMux I__14732 (
            .O(N__70350),
            .I(\quad_counter1.n30625 ));
    InMux I__14731 (
            .O(N__70347),
            .I(N__70343));
    InMux I__14730 (
            .O(N__70346),
            .I(N__70340));
    LocalMux I__14729 (
            .O(N__70343),
            .I(N__70334));
    LocalMux I__14728 (
            .O(N__70340),
            .I(N__70334));
    InMux I__14727 (
            .O(N__70339),
            .I(N__70331));
    Odrv4 I__14726 (
            .O(N__70334),
            .I(\quad_counter1.n3108 ));
    LocalMux I__14725 (
            .O(N__70331),
            .I(\quad_counter1.n3108 ));
    InMux I__14724 (
            .O(N__70326),
            .I(N__70323));
    LocalMux I__14723 (
            .O(N__70323),
            .I(N__70319));
    InMux I__14722 (
            .O(N__70322),
            .I(N__70316));
    Span4Mux_h I__14721 (
            .O(N__70319),
            .I(N__70310));
    LocalMux I__14720 (
            .O(N__70316),
            .I(N__70310));
    InMux I__14719 (
            .O(N__70315),
            .I(N__70307));
    Odrv4 I__14718 (
            .O(N__70310),
            .I(\quad_counter1.n3207 ));
    LocalMux I__14717 (
            .O(N__70307),
            .I(\quad_counter1.n3207 ));
    InMux I__14716 (
            .O(N__70302),
            .I(\quad_counter1.n30626 ));
    InMux I__14715 (
            .O(N__70299),
            .I(N__70295));
    InMux I__14714 (
            .O(N__70298),
            .I(N__70292));
    LocalMux I__14713 (
            .O(N__70295),
            .I(N__70286));
    LocalMux I__14712 (
            .O(N__70292),
            .I(N__70286));
    InMux I__14711 (
            .O(N__70291),
            .I(N__70283));
    Odrv4 I__14710 (
            .O(N__70286),
            .I(\quad_counter1.n3107 ));
    LocalMux I__14709 (
            .O(N__70283),
            .I(\quad_counter1.n3107 ));
    InMux I__14708 (
            .O(N__70278),
            .I(N__70274));
    InMux I__14707 (
            .O(N__70277),
            .I(N__70270));
    LocalMux I__14706 (
            .O(N__70274),
            .I(N__70267));
    CascadeMux I__14705 (
            .O(N__70273),
            .I(N__70264));
    LocalMux I__14704 (
            .O(N__70270),
            .I(N__70259));
    Span4Mux_h I__14703 (
            .O(N__70267),
            .I(N__70259));
    InMux I__14702 (
            .O(N__70264),
            .I(N__70256));
    Odrv4 I__14701 (
            .O(N__70259),
            .I(\quad_counter1.n3206 ));
    LocalMux I__14700 (
            .O(N__70256),
            .I(\quad_counter1.n3206 ));
    InMux I__14699 (
            .O(N__70251),
            .I(\quad_counter1.n30627 ));
    InMux I__14698 (
            .O(N__70248),
            .I(N__70243));
    InMux I__14697 (
            .O(N__70247),
            .I(N__70240));
    CascadeMux I__14696 (
            .O(N__70246),
            .I(N__70237));
    LocalMux I__14695 (
            .O(N__70243),
            .I(N__70232));
    LocalMux I__14694 (
            .O(N__70240),
            .I(N__70232));
    InMux I__14693 (
            .O(N__70237),
            .I(N__70229));
    Odrv4 I__14692 (
            .O(N__70232),
            .I(\quad_counter1.n3106 ));
    LocalMux I__14691 (
            .O(N__70229),
            .I(\quad_counter1.n3106 ));
    InMux I__14690 (
            .O(N__70224),
            .I(N__70220));
    InMux I__14689 (
            .O(N__70223),
            .I(N__70217));
    LocalMux I__14688 (
            .O(N__70220),
            .I(N__70214));
    LocalMux I__14687 (
            .O(N__70217),
            .I(N__70208));
    Span4Mux_h I__14686 (
            .O(N__70214),
            .I(N__70208));
    InMux I__14685 (
            .O(N__70213),
            .I(N__70205));
    Odrv4 I__14684 (
            .O(N__70208),
            .I(\quad_counter1.n3205 ));
    LocalMux I__14683 (
            .O(N__70205),
            .I(\quad_counter1.n3205 ));
    InMux I__14682 (
            .O(N__70200),
            .I(\quad_counter1.n30628 ));
    CascadeMux I__14681 (
            .O(N__70197),
            .I(\quad_counter1.n34587_cascade_ ));
    InMux I__14680 (
            .O(N__70194),
            .I(N__70191));
    LocalMux I__14679 (
            .O(N__70191),
            .I(\quad_counter1.n22_adj_4481 ));
    InMux I__14678 (
            .O(N__70188),
            .I(bfn_20_8_0_));
    InMux I__14677 (
            .O(N__70185),
            .I(N__70182));
    LocalMux I__14676 (
            .O(N__70182),
            .I(N__70178));
    InMux I__14675 (
            .O(N__70181),
            .I(N__70175));
    Span4Mux_v I__14674 (
            .O(N__70178),
            .I(N__70172));
    LocalMux I__14673 (
            .O(N__70175),
            .I(N__70169));
    Span4Mux_h I__14672 (
            .O(N__70172),
            .I(N__70163));
    Span4Mux_v I__14671 (
            .O(N__70169),
            .I(N__70163));
    InMux I__14670 (
            .O(N__70168),
            .I(N__70160));
    Odrv4 I__14669 (
            .O(N__70163),
            .I(\quad_counter1.n3119 ));
    LocalMux I__14668 (
            .O(N__70160),
            .I(\quad_counter1.n3119 ));
    InMux I__14667 (
            .O(N__70155),
            .I(\quad_counter1.n30615 ));
    InMux I__14666 (
            .O(N__70152),
            .I(N__70148));
    InMux I__14665 (
            .O(N__70151),
            .I(N__70145));
    LocalMux I__14664 (
            .O(N__70148),
            .I(N__70139));
    LocalMux I__14663 (
            .O(N__70145),
            .I(N__70139));
    CascadeMux I__14662 (
            .O(N__70144),
            .I(N__70136));
    Span4Mux_v I__14661 (
            .O(N__70139),
            .I(N__70133));
    InMux I__14660 (
            .O(N__70136),
            .I(N__70130));
    Odrv4 I__14659 (
            .O(N__70133),
            .I(\quad_counter1.n3118 ));
    LocalMux I__14658 (
            .O(N__70130),
            .I(\quad_counter1.n3118 ));
    InMux I__14657 (
            .O(N__70125),
            .I(\quad_counter1.n30616 ));
    InMux I__14656 (
            .O(N__70122),
            .I(N__70118));
    InMux I__14655 (
            .O(N__70121),
            .I(N__70115));
    LocalMux I__14654 (
            .O(N__70118),
            .I(N__70109));
    LocalMux I__14653 (
            .O(N__70115),
            .I(N__70109));
    InMux I__14652 (
            .O(N__70114),
            .I(N__70106));
    Span4Mux_h I__14651 (
            .O(N__70109),
            .I(N__70101));
    LocalMux I__14650 (
            .O(N__70106),
            .I(N__70101));
    Odrv4 I__14649 (
            .O(N__70101),
            .I(\quad_counter1.n3117 ));
    InMux I__14648 (
            .O(N__70098),
            .I(N__70094));
    InMux I__14647 (
            .O(N__70097),
            .I(N__70091));
    LocalMux I__14646 (
            .O(N__70094),
            .I(N__70088));
    LocalMux I__14645 (
            .O(N__70091),
            .I(N__70082));
    Span4Mux_h I__14644 (
            .O(N__70088),
            .I(N__70082));
    InMux I__14643 (
            .O(N__70087),
            .I(N__70079));
    Odrv4 I__14642 (
            .O(N__70082),
            .I(\quad_counter1.n3216 ));
    LocalMux I__14641 (
            .O(N__70079),
            .I(\quad_counter1.n3216 ));
    InMux I__14640 (
            .O(N__70074),
            .I(\quad_counter1.n30617 ));
    InMux I__14639 (
            .O(N__70071),
            .I(N__70066));
    InMux I__14638 (
            .O(N__70070),
            .I(N__70063));
    InMux I__14637 (
            .O(N__70069),
            .I(N__70060));
    LocalMux I__14636 (
            .O(N__70066),
            .I(N__70053));
    LocalMux I__14635 (
            .O(N__70063),
            .I(N__70053));
    LocalMux I__14634 (
            .O(N__70060),
            .I(N__70053));
    Odrv4 I__14633 (
            .O(N__70053),
            .I(\quad_counter1.n3116 ));
    InMux I__14632 (
            .O(N__70050),
            .I(N__70046));
    InMux I__14631 (
            .O(N__70049),
            .I(N__70043));
    LocalMux I__14630 (
            .O(N__70046),
            .I(N__70040));
    LocalMux I__14629 (
            .O(N__70043),
            .I(N__70034));
    Span4Mux_h I__14628 (
            .O(N__70040),
            .I(N__70034));
    InMux I__14627 (
            .O(N__70039),
            .I(N__70031));
    Odrv4 I__14626 (
            .O(N__70034),
            .I(\quad_counter1.n3215 ));
    LocalMux I__14625 (
            .O(N__70031),
            .I(\quad_counter1.n3215 ));
    InMux I__14624 (
            .O(N__70026),
            .I(\quad_counter1.n30618 ));
    InMux I__14623 (
            .O(N__70023),
            .I(N__70018));
    InMux I__14622 (
            .O(N__70022),
            .I(N__70015));
    CascadeMux I__14621 (
            .O(N__70021),
            .I(N__70012));
    LocalMux I__14620 (
            .O(N__70018),
            .I(N__70007));
    LocalMux I__14619 (
            .O(N__70015),
            .I(N__70007));
    InMux I__14618 (
            .O(N__70012),
            .I(N__70004));
    Span4Mux_v I__14617 (
            .O(N__70007),
            .I(N__69999));
    LocalMux I__14616 (
            .O(N__70004),
            .I(N__69999));
    Odrv4 I__14615 (
            .O(N__69999),
            .I(\quad_counter1.n3115 ));
    InMux I__14614 (
            .O(N__69996),
            .I(\quad_counter1.n30619 ));
    InMux I__14613 (
            .O(N__69993),
            .I(N__69988));
    InMux I__14612 (
            .O(N__69992),
            .I(N__69985));
    InMux I__14611 (
            .O(N__69991),
            .I(N__69982));
    LocalMux I__14610 (
            .O(N__69988),
            .I(N__69975));
    LocalMux I__14609 (
            .O(N__69985),
            .I(N__69975));
    LocalMux I__14608 (
            .O(N__69982),
            .I(N__69975));
    Odrv4 I__14607 (
            .O(N__69975),
            .I(\quad_counter1.n3114 ));
    CascadeMux I__14606 (
            .O(N__69972),
            .I(N__69964));
    CascadeMux I__14605 (
            .O(N__69971),
            .I(N__69961));
    CascadeMux I__14604 (
            .O(N__69970),
            .I(N__69958));
    CascadeMux I__14603 (
            .O(N__69969),
            .I(N__69955));
    CascadeMux I__14602 (
            .O(N__69968),
            .I(N__69952));
    CascadeMux I__14601 (
            .O(N__69967),
            .I(N__69949));
    InMux I__14600 (
            .O(N__69964),
            .I(N__69944));
    InMux I__14599 (
            .O(N__69961),
            .I(N__69944));
    InMux I__14598 (
            .O(N__69958),
            .I(N__69935));
    InMux I__14597 (
            .O(N__69955),
            .I(N__69935));
    InMux I__14596 (
            .O(N__69952),
            .I(N__69935));
    InMux I__14595 (
            .O(N__69949),
            .I(N__69935));
    LocalMux I__14594 (
            .O(N__69944),
            .I(\quad_counter1.n36152 ));
    LocalMux I__14593 (
            .O(N__69935),
            .I(\quad_counter1.n36152 ));
    InMux I__14592 (
            .O(N__69930),
            .I(N__69926));
    InMux I__14591 (
            .O(N__69929),
            .I(N__69923));
    LocalMux I__14590 (
            .O(N__69926),
            .I(N__69920));
    LocalMux I__14589 (
            .O(N__69923),
            .I(N__69914));
    Span4Mux_h I__14588 (
            .O(N__69920),
            .I(N__69914));
    InMux I__14587 (
            .O(N__69919),
            .I(N__69911));
    Odrv4 I__14586 (
            .O(N__69914),
            .I(\quad_counter1.n3213 ));
    LocalMux I__14585 (
            .O(N__69911),
            .I(\quad_counter1.n3213 ));
    InMux I__14584 (
            .O(N__69906),
            .I(\quad_counter1.n30620 ));
    InMux I__14583 (
            .O(N__69903),
            .I(N__69899));
    InMux I__14582 (
            .O(N__69902),
            .I(N__69896));
    LocalMux I__14581 (
            .O(N__69899),
            .I(N__69890));
    LocalMux I__14580 (
            .O(N__69896),
            .I(N__69890));
    InMux I__14579 (
            .O(N__69895),
            .I(N__69887));
    Span4Mux_v I__14578 (
            .O(N__69890),
            .I(N__69882));
    LocalMux I__14577 (
            .O(N__69887),
            .I(N__69882));
    Span4Mux_h I__14576 (
            .O(N__69882),
            .I(N__69879));
    Odrv4 I__14575 (
            .O(N__69879),
            .I(\quad_counter1.n3113 ));
    InMux I__14574 (
            .O(N__69876),
            .I(N__69872));
    InMux I__14573 (
            .O(N__69875),
            .I(N__69869));
    LocalMux I__14572 (
            .O(N__69872),
            .I(N__69866));
    LocalMux I__14571 (
            .O(N__69869),
            .I(N__69863));
    Span4Mux_v I__14570 (
            .O(N__69866),
            .I(N__69859));
    Span4Mux_v I__14569 (
            .O(N__69863),
            .I(N__69856));
    InMux I__14568 (
            .O(N__69862),
            .I(N__69853));
    Odrv4 I__14567 (
            .O(N__69859),
            .I(\quad_counter1.n3212 ));
    Odrv4 I__14566 (
            .O(N__69856),
            .I(\quad_counter1.n3212 ));
    LocalMux I__14565 (
            .O(N__69853),
            .I(\quad_counter1.n3212 ));
    InMux I__14564 (
            .O(N__69846),
            .I(\quad_counter1.n30559 ));
    InMux I__14563 (
            .O(N__69843),
            .I(\quad_counter1.n30560 ));
    InMux I__14562 (
            .O(N__69840),
            .I(N__69837));
    LocalMux I__14561 (
            .O(N__69837),
            .I(N__69832));
    InMux I__14560 (
            .O(N__69836),
            .I(N__69829));
    InMux I__14559 (
            .O(N__69835),
            .I(N__69826));
    Span4Mux_h I__14558 (
            .O(N__69832),
            .I(N__69823));
    LocalMux I__14557 (
            .O(N__69829),
            .I(N__69818));
    LocalMux I__14556 (
            .O(N__69826),
            .I(N__69818));
    Odrv4 I__14555 (
            .O(N__69823),
            .I(\quad_counter1.n2806 ));
    Odrv4 I__14554 (
            .O(N__69818),
            .I(\quad_counter1.n2806 ));
    InMux I__14553 (
            .O(N__69813),
            .I(\quad_counter1.n30561 ));
    InMux I__14552 (
            .O(N__69810),
            .I(N__69806));
    CascadeMux I__14551 (
            .O(N__69809),
            .I(N__69802));
    LocalMux I__14550 (
            .O(N__69806),
            .I(N__69799));
    InMux I__14549 (
            .O(N__69805),
            .I(N__69796));
    InMux I__14548 (
            .O(N__69802),
            .I(N__69793));
    Span4Mux_s2_v I__14547 (
            .O(N__69799),
            .I(N__69790));
    LocalMux I__14546 (
            .O(N__69796),
            .I(N__69785));
    LocalMux I__14545 (
            .O(N__69793),
            .I(N__69785));
    Odrv4 I__14544 (
            .O(N__69790),
            .I(\quad_counter1.n2805 ));
    Odrv4 I__14543 (
            .O(N__69785),
            .I(\quad_counter1.n2805 ));
    InMux I__14542 (
            .O(N__69780),
            .I(\quad_counter1.n30562 ));
    InMux I__14541 (
            .O(N__69777),
            .I(\quad_counter1.n30563 ));
    InMux I__14540 (
            .O(N__69774),
            .I(N__69769));
    InMux I__14539 (
            .O(N__69773),
            .I(N__69766));
    InMux I__14538 (
            .O(N__69772),
            .I(N__69763));
    LocalMux I__14537 (
            .O(N__69769),
            .I(N__69760));
    LocalMux I__14536 (
            .O(N__69766),
            .I(\quad_counter1.n2804 ));
    LocalMux I__14535 (
            .O(N__69763),
            .I(\quad_counter1.n2804 ));
    Odrv4 I__14534 (
            .O(N__69760),
            .I(\quad_counter1.n2804 ));
    InMux I__14533 (
            .O(N__69753),
            .I(N__69750));
    LocalMux I__14532 (
            .O(N__69750),
            .I(\quad_counter1.n26_adj_4482 ));
    CascadeMux I__14531 (
            .O(N__69747),
            .I(\quad_counter1.n3134_cascade_ ));
    InMux I__14530 (
            .O(N__69744),
            .I(N__69741));
    LocalMux I__14529 (
            .O(N__69741),
            .I(\quad_counter1.n8_adj_4477 ));
    InMux I__14528 (
            .O(N__69738),
            .I(N__69735));
    LocalMux I__14527 (
            .O(N__69735),
            .I(\quad_counter1.n7_adj_4478 ));
    InMux I__14526 (
            .O(N__69732),
            .I(N__69728));
    InMux I__14525 (
            .O(N__69731),
            .I(N__69725));
    LocalMux I__14524 (
            .O(N__69728),
            .I(N__69721));
    LocalMux I__14523 (
            .O(N__69725),
            .I(N__69718));
    InMux I__14522 (
            .O(N__69724),
            .I(N__69715));
    Odrv4 I__14521 (
            .O(N__69721),
            .I(\quad_counter1.n2816 ));
    Odrv4 I__14520 (
            .O(N__69718),
            .I(\quad_counter1.n2816 ));
    LocalMux I__14519 (
            .O(N__69715),
            .I(\quad_counter1.n2816 ));
    InMux I__14518 (
            .O(N__69708),
            .I(\quad_counter1.n30551 ));
    InMux I__14517 (
            .O(N__69705),
            .I(N__69701));
    InMux I__14516 (
            .O(N__69704),
            .I(N__69698));
    LocalMux I__14515 (
            .O(N__69701),
            .I(N__69692));
    LocalMux I__14514 (
            .O(N__69698),
            .I(N__69692));
    InMux I__14513 (
            .O(N__69697),
            .I(N__69689));
    Odrv4 I__14512 (
            .O(N__69692),
            .I(\quad_counter1.n2815 ));
    LocalMux I__14511 (
            .O(N__69689),
            .I(\quad_counter1.n2815 ));
    InMux I__14510 (
            .O(N__69684),
            .I(\quad_counter1.n30552 ));
    InMux I__14509 (
            .O(N__69681),
            .I(N__69678));
    LocalMux I__14508 (
            .O(N__69678),
            .I(N__69674));
    InMux I__14507 (
            .O(N__69677),
            .I(N__69671));
    Span4Mux_s1_v I__14506 (
            .O(N__69674),
            .I(N__69667));
    LocalMux I__14505 (
            .O(N__69671),
            .I(N__69664));
    InMux I__14504 (
            .O(N__69670),
            .I(N__69661));
    Odrv4 I__14503 (
            .O(N__69667),
            .I(\quad_counter1.n2814 ));
    Odrv4 I__14502 (
            .O(N__69664),
            .I(\quad_counter1.n2814 ));
    LocalMux I__14501 (
            .O(N__69661),
            .I(\quad_counter1.n2814 ));
    InMux I__14500 (
            .O(N__69654),
            .I(\quad_counter1.n30553 ));
    InMux I__14499 (
            .O(N__69651),
            .I(\quad_counter1.n30554 ));
    InMux I__14498 (
            .O(N__69648),
            .I(N__69643));
    InMux I__14497 (
            .O(N__69647),
            .I(N__69640));
    InMux I__14496 (
            .O(N__69646),
            .I(N__69637));
    LocalMux I__14495 (
            .O(N__69643),
            .I(\quad_counter1.n2812 ));
    LocalMux I__14494 (
            .O(N__69640),
            .I(\quad_counter1.n2812 ));
    LocalMux I__14493 (
            .O(N__69637),
            .I(\quad_counter1.n2812 ));
    InMux I__14492 (
            .O(N__69630),
            .I(\quad_counter1.n30555 ));
    InMux I__14491 (
            .O(N__69627),
            .I(bfn_20_5_0_));
    InMux I__14490 (
            .O(N__69624),
            .I(\quad_counter1.n30557 ));
    InMux I__14489 (
            .O(N__69621),
            .I(N__69616));
    InMux I__14488 (
            .O(N__69620),
            .I(N__69613));
    InMux I__14487 (
            .O(N__69619),
            .I(N__69610));
    LocalMux I__14486 (
            .O(N__69616),
            .I(N__69607));
    LocalMux I__14485 (
            .O(N__69613),
            .I(N__69602));
    LocalMux I__14484 (
            .O(N__69610),
            .I(N__69602));
    Odrv4 I__14483 (
            .O(N__69607),
            .I(\quad_counter1.n2809 ));
    Odrv4 I__14482 (
            .O(N__69602),
            .I(\quad_counter1.n2809 ));
    InMux I__14481 (
            .O(N__69597),
            .I(\quad_counter1.n30558 ));
    InMux I__14480 (
            .O(N__69594),
            .I(N__69589));
    InMux I__14479 (
            .O(N__69593),
            .I(N__69586));
    InMux I__14478 (
            .O(N__69592),
            .I(N__69583));
    LocalMux I__14477 (
            .O(N__69589),
            .I(N__69580));
    LocalMux I__14476 (
            .O(N__69586),
            .I(N__69575));
    LocalMux I__14475 (
            .O(N__69583),
            .I(N__69575));
    Odrv4 I__14474 (
            .O(N__69580),
            .I(\quad_counter1.n2808 ));
    Odrv4 I__14473 (
            .O(N__69575),
            .I(\quad_counter1.n2808 ));
    CascadeMux I__14472 (
            .O(N__69570),
            .I(N__69562));
    CascadeMux I__14471 (
            .O(N__69569),
            .I(N__69559));
    CascadeMux I__14470 (
            .O(N__69568),
            .I(N__69556));
    CascadeMux I__14469 (
            .O(N__69567),
            .I(N__69553));
    CascadeMux I__14468 (
            .O(N__69566),
            .I(N__69550));
    CascadeMux I__14467 (
            .O(N__69565),
            .I(N__69547));
    InMux I__14466 (
            .O(N__69562),
            .I(N__69542));
    InMux I__14465 (
            .O(N__69559),
            .I(N__69542));
    InMux I__14464 (
            .O(N__69556),
            .I(N__69533));
    InMux I__14463 (
            .O(N__69553),
            .I(N__69533));
    InMux I__14462 (
            .O(N__69550),
            .I(N__69533));
    InMux I__14461 (
            .O(N__69547),
            .I(N__69533));
    LocalMux I__14460 (
            .O(N__69542),
            .I(\quad_counter1.n36131 ));
    LocalMux I__14459 (
            .O(N__69533),
            .I(\quad_counter1.n36131 ));
    CascadeMux I__14458 (
            .O(N__69528),
            .I(\quad_counter1.n19_cascade_ ));
    CascadeMux I__14457 (
            .O(N__69525),
            .I(N__69512));
    CascadeMux I__14456 (
            .O(N__69524),
            .I(N__69509));
    CascadeMux I__14455 (
            .O(N__69523),
            .I(N__69506));
    CascadeMux I__14454 (
            .O(N__69522),
            .I(N__69503));
    CascadeMux I__14453 (
            .O(N__69521),
            .I(N__69500));
    CascadeMux I__14452 (
            .O(N__69520),
            .I(N__69497));
    CascadeMux I__14451 (
            .O(N__69519),
            .I(N__69494));
    CascadeMux I__14450 (
            .O(N__69518),
            .I(N__69491));
    CascadeMux I__14449 (
            .O(N__69517),
            .I(N__69488));
    CascadeMux I__14448 (
            .O(N__69516),
            .I(N__69485));
    CascadeMux I__14447 (
            .O(N__69515),
            .I(N__69482));
    InMux I__14446 (
            .O(N__69512),
            .I(N__69477));
    InMux I__14445 (
            .O(N__69509),
            .I(N__69477));
    InMux I__14444 (
            .O(N__69506),
            .I(N__69473));
    InMux I__14443 (
            .O(N__69503),
            .I(N__69464));
    InMux I__14442 (
            .O(N__69500),
            .I(N__69464));
    InMux I__14441 (
            .O(N__69497),
            .I(N__69464));
    InMux I__14440 (
            .O(N__69494),
            .I(N__69464));
    InMux I__14439 (
            .O(N__69491),
            .I(N__69455));
    InMux I__14438 (
            .O(N__69488),
            .I(N__69455));
    InMux I__14437 (
            .O(N__69485),
            .I(N__69455));
    InMux I__14436 (
            .O(N__69482),
            .I(N__69455));
    LocalMux I__14435 (
            .O(N__69477),
            .I(N__69452));
    InMux I__14434 (
            .O(N__69476),
            .I(N__69449));
    LocalMux I__14433 (
            .O(N__69473),
            .I(\quad_counter1.n2837 ));
    LocalMux I__14432 (
            .O(N__69464),
            .I(\quad_counter1.n2837 ));
    LocalMux I__14431 (
            .O(N__69455),
            .I(\quad_counter1.n2837 ));
    Odrv4 I__14430 (
            .O(N__69452),
            .I(\quad_counter1.n2837 ));
    LocalMux I__14429 (
            .O(N__69449),
            .I(\quad_counter1.n2837 ));
    CascadeMux I__14428 (
            .O(N__69438),
            .I(\quad_counter1.n28267_cascade_ ));
    CascadeMux I__14427 (
            .O(N__69435),
            .I(\quad_counter1.n10_adj_4455_cascade_ ));
    InMux I__14426 (
            .O(N__69432),
            .I(N__69429));
    LocalMux I__14425 (
            .O(N__69429),
            .I(\quad_counter1.n12_adj_4456 ));
    InMux I__14424 (
            .O(N__69426),
            .I(N__69421));
    InMux I__14423 (
            .O(N__69425),
            .I(N__69418));
    CascadeMux I__14422 (
            .O(N__69424),
            .I(N__69415));
    LocalMux I__14421 (
            .O(N__69421),
            .I(N__69410));
    LocalMux I__14420 (
            .O(N__69418),
            .I(N__69410));
    InMux I__14419 (
            .O(N__69415),
            .I(N__69407));
    Odrv4 I__14418 (
            .O(N__69410),
            .I(\quad_counter1.n2819 ));
    LocalMux I__14417 (
            .O(N__69407),
            .I(\quad_counter1.n2819 ));
    InMux I__14416 (
            .O(N__69402),
            .I(bfn_20_4_0_));
    InMux I__14415 (
            .O(N__69399),
            .I(N__69395));
    InMux I__14414 (
            .O(N__69398),
            .I(N__69392));
    LocalMux I__14413 (
            .O(N__69395),
            .I(N__69386));
    LocalMux I__14412 (
            .O(N__69392),
            .I(N__69386));
    InMux I__14411 (
            .O(N__69391),
            .I(N__69383));
    Odrv4 I__14410 (
            .O(N__69386),
            .I(\quad_counter1.n2818 ));
    LocalMux I__14409 (
            .O(N__69383),
            .I(\quad_counter1.n2818 ));
    InMux I__14408 (
            .O(N__69378),
            .I(\quad_counter1.n30549 ));
    InMux I__14407 (
            .O(N__69375),
            .I(N__69371));
    InMux I__14406 (
            .O(N__69374),
            .I(N__69368));
    LocalMux I__14405 (
            .O(N__69371),
            .I(N__69362));
    LocalMux I__14404 (
            .O(N__69368),
            .I(N__69362));
    InMux I__14403 (
            .O(N__69367),
            .I(N__69359));
    Odrv4 I__14402 (
            .O(N__69362),
            .I(\quad_counter1.n2817 ));
    LocalMux I__14401 (
            .O(N__69359),
            .I(\quad_counter1.n2817 ));
    InMux I__14400 (
            .O(N__69354),
            .I(\quad_counter1.n30550 ));
    InMux I__14399 (
            .O(N__69351),
            .I(N__69346));
    InMux I__14398 (
            .O(N__69350),
            .I(N__69343));
    InMux I__14397 (
            .O(N__69349),
            .I(N__69340));
    LocalMux I__14396 (
            .O(N__69346),
            .I(\c0.n31784 ));
    LocalMux I__14395 (
            .O(N__69343),
            .I(\c0.n31784 ));
    LocalMux I__14394 (
            .O(N__69340),
            .I(\c0.n31784 ));
    InMux I__14393 (
            .O(N__69333),
            .I(N__69330));
    LocalMux I__14392 (
            .O(N__69330),
            .I(\c0.n17_adj_4753 ));
    CascadeMux I__14391 (
            .O(N__69327),
            .I(\c0.n4_adj_4751_cascade_ ));
    InMux I__14390 (
            .O(N__69324),
            .I(N__69321));
    LocalMux I__14389 (
            .O(N__69321),
            .I(N__69318));
    Odrv4 I__14388 (
            .O(N__69318),
            .I(\c0.n20_adj_4754 ));
    CascadeMux I__14387 (
            .O(N__69315),
            .I(N__69312));
    InMux I__14386 (
            .O(N__69312),
            .I(N__69306));
    InMux I__14385 (
            .O(N__69311),
            .I(N__69306));
    LocalMux I__14384 (
            .O(N__69306),
            .I(\c0.data_in_frame_29_7 ));
    CascadeMux I__14383 (
            .O(N__69303),
            .I(N__69300));
    InMux I__14382 (
            .O(N__69300),
            .I(N__69296));
    CascadeMux I__14381 (
            .O(N__69299),
            .I(N__69293));
    LocalMux I__14380 (
            .O(N__69296),
            .I(N__69289));
    InMux I__14379 (
            .O(N__69293),
            .I(N__69284));
    InMux I__14378 (
            .O(N__69292),
            .I(N__69284));
    Odrv12 I__14377 (
            .O(N__69289),
            .I(\c0.data_in_frame_27_6 ));
    LocalMux I__14376 (
            .O(N__69284),
            .I(\c0.data_in_frame_27_6 ));
    InMux I__14375 (
            .O(N__69279),
            .I(N__69276));
    LocalMux I__14374 (
            .O(N__69276),
            .I(N__69272));
    InMux I__14373 (
            .O(N__69275),
            .I(N__69269));
    Span4Mux_h I__14372 (
            .O(N__69272),
            .I(N__69264));
    LocalMux I__14371 (
            .O(N__69269),
            .I(N__69264));
    Odrv4 I__14370 (
            .O(N__69264),
            .I(\c0.n33463 ));
    InMux I__14369 (
            .O(N__69261),
            .I(N__69258));
    LocalMux I__14368 (
            .O(N__69258),
            .I(N__69255));
    Span4Mux_h I__14367 (
            .O(N__69255),
            .I(N__69252));
    Odrv4 I__14366 (
            .O(N__69252),
            .I(\c0.n35250 ));
    InMux I__14365 (
            .O(N__69249),
            .I(N__69245));
    CascadeMux I__14364 (
            .O(N__69248),
            .I(N__69241));
    LocalMux I__14363 (
            .O(N__69245),
            .I(N__69238));
    InMux I__14362 (
            .O(N__69244),
            .I(N__69235));
    InMux I__14361 (
            .O(N__69241),
            .I(N__69232));
    Span4Mux_h I__14360 (
            .O(N__69238),
            .I(N__69229));
    LocalMux I__14359 (
            .O(N__69235),
            .I(N__69226));
    LocalMux I__14358 (
            .O(N__69232),
            .I(N__69221));
    Span4Mux_v I__14357 (
            .O(N__69229),
            .I(N__69221));
    Span4Mux_v I__14356 (
            .O(N__69226),
            .I(N__69218));
    Odrv4 I__14355 (
            .O(N__69221),
            .I(\c0.data_in_frame_26_0 ));
    Odrv4 I__14354 (
            .O(N__69218),
            .I(\c0.data_in_frame_26_0 ));
    InMux I__14353 (
            .O(N__69213),
            .I(N__69209));
    InMux I__14352 (
            .O(N__69212),
            .I(N__69206));
    LocalMux I__14351 (
            .O(N__69209),
            .I(N__69203));
    LocalMux I__14350 (
            .O(N__69206),
            .I(N__69200));
    Odrv12 I__14349 (
            .O(N__69203),
            .I(\c0.n33846 ));
    Odrv4 I__14348 (
            .O(N__69200),
            .I(\c0.n33846 ));
    InMux I__14347 (
            .O(N__69195),
            .I(N__69192));
    LocalMux I__14346 (
            .O(N__69192),
            .I(N__69189));
    Odrv4 I__14345 (
            .O(N__69189),
            .I(\c0.n33490 ));
    InMux I__14344 (
            .O(N__69186),
            .I(N__69183));
    LocalMux I__14343 (
            .O(N__69183),
            .I(\c0.n33816 ));
    CascadeMux I__14342 (
            .O(N__69180),
            .I(N__69176));
    CascadeMux I__14341 (
            .O(N__69179),
            .I(N__69173));
    InMux I__14340 (
            .O(N__69176),
            .I(N__69170));
    InMux I__14339 (
            .O(N__69173),
            .I(N__69167));
    LocalMux I__14338 (
            .O(N__69170),
            .I(\c0.data_in_frame_28_7 ));
    LocalMux I__14337 (
            .O(N__69167),
            .I(\c0.data_in_frame_28_7 ));
    InMux I__14336 (
            .O(N__69162),
            .I(N__69159));
    LocalMux I__14335 (
            .O(N__69159),
            .I(N__69155));
    InMux I__14334 (
            .O(N__69158),
            .I(N__69152));
    Odrv4 I__14333 (
            .O(N__69155),
            .I(\c0.n33976 ));
    LocalMux I__14332 (
            .O(N__69152),
            .I(\c0.n33976 ));
    CascadeMux I__14331 (
            .O(N__69147),
            .I(\c0.n16_adj_4750_cascade_ ));
    InMux I__14330 (
            .O(N__69144),
            .I(N__69141));
    LocalMux I__14329 (
            .O(N__69141),
            .I(\c0.n18_adj_4752 ));
    InMux I__14328 (
            .O(N__69138),
            .I(N__69135));
    LocalMux I__14327 (
            .O(N__69135),
            .I(N__69131));
    InMux I__14326 (
            .O(N__69134),
            .I(N__69126));
    Span4Mux_h I__14325 (
            .O(N__69131),
            .I(N__69123));
    InMux I__14324 (
            .O(N__69130),
            .I(N__69118));
    InMux I__14323 (
            .O(N__69129),
            .I(N__69118));
    LocalMux I__14322 (
            .O(N__69126),
            .I(\c0.data_in_frame_27_4 ));
    Odrv4 I__14321 (
            .O(N__69123),
            .I(\c0.data_in_frame_27_4 ));
    LocalMux I__14320 (
            .O(N__69118),
            .I(\c0.data_in_frame_27_4 ));
    InMux I__14319 (
            .O(N__69111),
            .I(N__69106));
    InMux I__14318 (
            .O(N__69110),
            .I(N__69101));
    InMux I__14317 (
            .O(N__69109),
            .I(N__69101));
    LocalMux I__14316 (
            .O(N__69106),
            .I(\c0.data_in_frame_27_0 ));
    LocalMux I__14315 (
            .O(N__69101),
            .I(\c0.data_in_frame_27_0 ));
    CascadeMux I__14314 (
            .O(N__69096),
            .I(N__69092));
    InMux I__14313 (
            .O(N__69095),
            .I(N__69087));
    InMux I__14312 (
            .O(N__69092),
            .I(N__69087));
    LocalMux I__14311 (
            .O(N__69087),
            .I(\c0.data_in_frame_26_6 ));
    InMux I__14310 (
            .O(N__69084),
            .I(N__69080));
    InMux I__14309 (
            .O(N__69083),
            .I(N__69076));
    LocalMux I__14308 (
            .O(N__69080),
            .I(N__69072));
    InMux I__14307 (
            .O(N__69079),
            .I(N__69069));
    LocalMux I__14306 (
            .O(N__69076),
            .I(N__69066));
    InMux I__14305 (
            .O(N__69075),
            .I(N__69063));
    Span4Mux_v I__14304 (
            .O(N__69072),
            .I(N__69058));
    LocalMux I__14303 (
            .O(N__69069),
            .I(N__69058));
    Span4Mux_h I__14302 (
            .O(N__69066),
            .I(N__69055));
    LocalMux I__14301 (
            .O(N__69063),
            .I(N__69050));
    Span4Mux_h I__14300 (
            .O(N__69058),
            .I(N__69050));
    Odrv4 I__14299 (
            .O(N__69055),
            .I(\c0.n33374 ));
    Odrv4 I__14298 (
            .O(N__69050),
            .I(\c0.n33374 ));
    InMux I__14297 (
            .O(N__69045),
            .I(N__69041));
    InMux I__14296 (
            .O(N__69044),
            .I(N__69038));
    LocalMux I__14295 (
            .O(N__69041),
            .I(N__69035));
    LocalMux I__14294 (
            .O(N__69038),
            .I(N__69029));
    Span4Mux_h I__14293 (
            .O(N__69035),
            .I(N__69029));
    InMux I__14292 (
            .O(N__69034),
            .I(N__69026));
    Odrv4 I__14291 (
            .O(N__69029),
            .I(\c0.data_in_frame_26_4 ));
    LocalMux I__14290 (
            .O(N__69026),
            .I(\c0.data_in_frame_26_4 ));
    CascadeMux I__14289 (
            .O(N__69021),
            .I(N__69018));
    InMux I__14288 (
            .O(N__69018),
            .I(N__69014));
    InMux I__14287 (
            .O(N__69017),
            .I(N__69009));
    LocalMux I__14286 (
            .O(N__69014),
            .I(N__69006));
    InMux I__14285 (
            .O(N__69013),
            .I(N__69001));
    InMux I__14284 (
            .O(N__69012),
            .I(N__69001));
    LocalMux I__14283 (
            .O(N__69009),
            .I(N__68998));
    Odrv12 I__14282 (
            .O(N__69006),
            .I(\c0.data_in_frame_22_2 ));
    LocalMux I__14281 (
            .O(N__69001),
            .I(\c0.data_in_frame_22_2 ));
    Odrv4 I__14280 (
            .O(N__68998),
            .I(\c0.data_in_frame_22_2 ));
    InMux I__14279 (
            .O(N__68991),
            .I(N__68988));
    LocalMux I__14278 (
            .O(N__68988),
            .I(N__68985));
    Span4Mux_h I__14277 (
            .O(N__68985),
            .I(N__68981));
    InMux I__14276 (
            .O(N__68984),
            .I(N__68978));
    Odrv4 I__14275 (
            .O(N__68981),
            .I(\c0.n33849 ));
    LocalMux I__14274 (
            .O(N__68978),
            .I(\c0.n33849 ));
    InMux I__14273 (
            .O(N__68973),
            .I(N__68969));
    InMux I__14272 (
            .O(N__68972),
            .I(N__68966));
    LocalMux I__14271 (
            .O(N__68969),
            .I(N__68963));
    LocalMux I__14270 (
            .O(N__68966),
            .I(N__68960));
    Odrv12 I__14269 (
            .O(N__68963),
            .I(\c0.n18193 ));
    Odrv4 I__14268 (
            .O(N__68960),
            .I(\c0.n18193 ));
    InMux I__14267 (
            .O(N__68955),
            .I(N__68948));
    InMux I__14266 (
            .O(N__68954),
            .I(N__68948));
    InMux I__14265 (
            .O(N__68953),
            .I(N__68945));
    LocalMux I__14264 (
            .O(N__68948),
            .I(\c0.n33775 ));
    LocalMux I__14263 (
            .O(N__68945),
            .I(\c0.n33775 ));
    CascadeMux I__14262 (
            .O(N__68940),
            .I(N__68936));
    CascadeMux I__14261 (
            .O(N__68939),
            .I(N__68933));
    InMux I__14260 (
            .O(N__68936),
            .I(N__68930));
    InMux I__14259 (
            .O(N__68933),
            .I(N__68927));
    LocalMux I__14258 (
            .O(N__68930),
            .I(N__68924));
    LocalMux I__14257 (
            .O(N__68927),
            .I(N__68921));
    Span4Mux_h I__14256 (
            .O(N__68924),
            .I(N__68918));
    Odrv12 I__14255 (
            .O(N__68921),
            .I(\c0.n33350 ));
    Odrv4 I__14254 (
            .O(N__68918),
            .I(\c0.n33350 ));
    InMux I__14253 (
            .O(N__68913),
            .I(N__68905));
    InMux I__14252 (
            .O(N__68912),
            .I(N__68905));
    InMux I__14251 (
            .O(N__68911),
            .I(N__68902));
    InMux I__14250 (
            .O(N__68910),
            .I(N__68899));
    LocalMux I__14249 (
            .O(N__68905),
            .I(N__68896));
    LocalMux I__14248 (
            .O(N__68902),
            .I(N__68892));
    LocalMux I__14247 (
            .O(N__68899),
            .I(N__68887));
    Span4Mux_h I__14246 (
            .O(N__68896),
            .I(N__68887));
    InMux I__14245 (
            .O(N__68895),
            .I(N__68884));
    Span4Mux_h I__14244 (
            .O(N__68892),
            .I(N__68881));
    Span4Mux_h I__14243 (
            .O(N__68887),
            .I(N__68878));
    LocalMux I__14242 (
            .O(N__68884),
            .I(\c0.n32339 ));
    Odrv4 I__14241 (
            .O(N__68881),
            .I(\c0.n32339 ));
    Odrv4 I__14240 (
            .O(N__68878),
            .I(\c0.n32339 ));
    InMux I__14239 (
            .O(N__68871),
            .I(N__68868));
    LocalMux I__14238 (
            .O(N__68868),
            .I(N__68865));
    Span4Mux_h I__14237 (
            .O(N__68865),
            .I(N__68862));
    Span4Mux_h I__14236 (
            .O(N__68862),
            .I(N__68859));
    Odrv4 I__14235 (
            .O(N__68859),
            .I(\c0.n8_adj_4540 ));
    InMux I__14234 (
            .O(N__68856),
            .I(N__68853));
    LocalMux I__14233 (
            .O(N__68853),
            .I(N__68850));
    Odrv4 I__14232 (
            .O(N__68850),
            .I(\c0.n18596 ));
    InMux I__14231 (
            .O(N__68847),
            .I(N__68844));
    LocalMux I__14230 (
            .O(N__68844),
            .I(N__68841));
    Odrv4 I__14229 (
            .O(N__68841),
            .I(\c0.n16120 ));
    InMux I__14228 (
            .O(N__68838),
            .I(N__68835));
    LocalMux I__14227 (
            .O(N__68835),
            .I(N__68832));
    Span4Mux_h I__14226 (
            .O(N__68832),
            .I(N__68829));
    Odrv4 I__14225 (
            .O(N__68829),
            .I(\c0.n6_adj_4756 ));
    CascadeMux I__14224 (
            .O(N__68826),
            .I(N__68822));
    InMux I__14223 (
            .O(N__68825),
            .I(N__68818));
    InMux I__14222 (
            .O(N__68822),
            .I(N__68813));
    InMux I__14221 (
            .O(N__68821),
            .I(N__68813));
    LocalMux I__14220 (
            .O(N__68818),
            .I(N__68808));
    LocalMux I__14219 (
            .O(N__68813),
            .I(N__68808));
    Span4Mux_h I__14218 (
            .O(N__68808),
            .I(N__68804));
    InMux I__14217 (
            .O(N__68807),
            .I(N__68801));
    Span4Mux_h I__14216 (
            .O(N__68804),
            .I(N__68798));
    LocalMux I__14215 (
            .O(N__68801),
            .I(\c0.data_in_frame_27_2 ));
    Odrv4 I__14214 (
            .O(N__68798),
            .I(\c0.data_in_frame_27_2 ));
    InMux I__14213 (
            .O(N__68793),
            .I(N__68790));
    LocalMux I__14212 (
            .O(N__68790),
            .I(N__68786));
    InMux I__14211 (
            .O(N__68789),
            .I(N__68782));
    Span4Mux_v I__14210 (
            .O(N__68786),
            .I(N__68779));
    InMux I__14209 (
            .O(N__68785),
            .I(N__68776));
    LocalMux I__14208 (
            .O(N__68782),
            .I(N__68773));
    Odrv4 I__14207 (
            .O(N__68779),
            .I(\c0.n18568 ));
    LocalMux I__14206 (
            .O(N__68776),
            .I(\c0.n18568 ));
    Odrv12 I__14205 (
            .O(N__68773),
            .I(\c0.n18568 ));
    InMux I__14204 (
            .O(N__68766),
            .I(N__68763));
    LocalMux I__14203 (
            .O(N__68763),
            .I(N__68760));
    Span4Mux_v I__14202 (
            .O(N__68760),
            .I(N__68757));
    Span4Mux_h I__14201 (
            .O(N__68757),
            .I(N__68754));
    Odrv4 I__14200 (
            .O(N__68754),
            .I(\c0.n35416 ));
    InMux I__14199 (
            .O(N__68751),
            .I(N__68748));
    LocalMux I__14198 (
            .O(N__68748),
            .I(N__68745));
    Odrv4 I__14197 (
            .O(N__68745),
            .I(n2315));
    InMux I__14196 (
            .O(N__68742),
            .I(N__68739));
    LocalMux I__14195 (
            .O(N__68739),
            .I(N__68735));
    CascadeMux I__14194 (
            .O(N__68738),
            .I(N__68732));
    Span4Mux_h I__14193 (
            .O(N__68735),
            .I(N__68728));
    InMux I__14192 (
            .O(N__68732),
            .I(N__68723));
    InMux I__14191 (
            .O(N__68731),
            .I(N__68723));
    Odrv4 I__14190 (
            .O(N__68728),
            .I(\c0.data_in_frame_27_7 ));
    LocalMux I__14189 (
            .O(N__68723),
            .I(\c0.data_in_frame_27_7 ));
    CascadeMux I__14188 (
            .O(N__68718),
            .I(N__68715));
    InMux I__14187 (
            .O(N__68715),
            .I(N__68711));
    CascadeMux I__14186 (
            .O(N__68714),
            .I(N__68707));
    LocalMux I__14185 (
            .O(N__68711),
            .I(N__68703));
    InMux I__14184 (
            .O(N__68710),
            .I(N__68700));
    InMux I__14183 (
            .O(N__68707),
            .I(N__68695));
    InMux I__14182 (
            .O(N__68706),
            .I(N__68695));
    Odrv4 I__14181 (
            .O(N__68703),
            .I(\c0.data_in_frame_25_4 ));
    LocalMux I__14180 (
            .O(N__68700),
            .I(\c0.data_in_frame_25_4 ));
    LocalMux I__14179 (
            .O(N__68695),
            .I(\c0.data_in_frame_25_4 ));
    InMux I__14178 (
            .O(N__68688),
            .I(N__68684));
    InMux I__14177 (
            .O(N__68687),
            .I(N__68681));
    LocalMux I__14176 (
            .O(N__68684),
            .I(N__68678));
    LocalMux I__14175 (
            .O(N__68681),
            .I(N__68675));
    Span4Mux_h I__14174 (
            .O(N__68678),
            .I(N__68672));
    Odrv4 I__14173 (
            .O(N__68675),
            .I(\c0.n33594 ));
    Odrv4 I__14172 (
            .O(N__68672),
            .I(\c0.n33594 ));
    InMux I__14171 (
            .O(N__68667),
            .I(N__68664));
    LocalMux I__14170 (
            .O(N__68664),
            .I(N__68659));
    InMux I__14169 (
            .O(N__68663),
            .I(N__68656));
    InMux I__14168 (
            .O(N__68662),
            .I(N__68652));
    Span4Mux_v I__14167 (
            .O(N__68659),
            .I(N__68647));
    LocalMux I__14166 (
            .O(N__68656),
            .I(N__68647));
    InMux I__14165 (
            .O(N__68655),
            .I(N__68644));
    LocalMux I__14164 (
            .O(N__68652),
            .I(N__68641));
    Span4Mux_v I__14163 (
            .O(N__68647),
            .I(N__68638));
    LocalMux I__14162 (
            .O(N__68644),
            .I(\c0.data_in_frame_24_4 ));
    Odrv12 I__14161 (
            .O(N__68641),
            .I(\c0.data_in_frame_24_4 ));
    Odrv4 I__14160 (
            .O(N__68638),
            .I(\c0.data_in_frame_24_4 ));
    InMux I__14159 (
            .O(N__68631),
            .I(N__68625));
    InMux I__14158 (
            .O(N__68630),
            .I(N__68625));
    LocalMux I__14157 (
            .O(N__68625),
            .I(\c0.n34009 ));
    CascadeMux I__14156 (
            .O(N__68622),
            .I(\c0.n34009_cascade_ ));
    InMux I__14155 (
            .O(N__68619),
            .I(N__68615));
    InMux I__14154 (
            .O(N__68618),
            .I(N__68612));
    LocalMux I__14153 (
            .O(N__68615),
            .I(N__68609));
    LocalMux I__14152 (
            .O(N__68612),
            .I(\c0.n31355 ));
    Odrv12 I__14151 (
            .O(N__68609),
            .I(\c0.n31355 ));
    CascadeMux I__14150 (
            .O(N__68604),
            .I(N__68601));
    InMux I__14149 (
            .O(N__68601),
            .I(N__68595));
    InMux I__14148 (
            .O(N__68600),
            .I(N__68595));
    LocalMux I__14147 (
            .O(N__68595),
            .I(N__68591));
    InMux I__14146 (
            .O(N__68594),
            .I(N__68585));
    Span4Mux_h I__14145 (
            .O(N__68591),
            .I(N__68582));
    InMux I__14144 (
            .O(N__68590),
            .I(N__68575));
    InMux I__14143 (
            .O(N__68589),
            .I(N__68575));
    InMux I__14142 (
            .O(N__68588),
            .I(N__68572));
    LocalMux I__14141 (
            .O(N__68585),
            .I(N__68567));
    Span4Mux_h I__14140 (
            .O(N__68582),
            .I(N__68567));
    InMux I__14139 (
            .O(N__68581),
            .I(N__68564));
    InMux I__14138 (
            .O(N__68580),
            .I(N__68560));
    LocalMux I__14137 (
            .O(N__68575),
            .I(N__68557));
    LocalMux I__14136 (
            .O(N__68572),
            .I(N__68554));
    Span4Mux_v I__14135 (
            .O(N__68567),
            .I(N__68551));
    LocalMux I__14134 (
            .O(N__68564),
            .I(N__68548));
    InMux I__14133 (
            .O(N__68563),
            .I(N__68545));
    LocalMux I__14132 (
            .O(N__68560),
            .I(N__68540));
    Span4Mux_v I__14131 (
            .O(N__68557),
            .I(N__68540));
    Span4Mux_h I__14130 (
            .O(N__68554),
            .I(N__68535));
    Span4Mux_h I__14129 (
            .O(N__68551),
            .I(N__68535));
    Span4Mux_h I__14128 (
            .O(N__68548),
            .I(N__68532));
    LocalMux I__14127 (
            .O(N__68545),
            .I(\c0.n12_adj_4526 ));
    Odrv4 I__14126 (
            .O(N__68540),
            .I(\c0.n12_adj_4526 ));
    Odrv4 I__14125 (
            .O(N__68535),
            .I(\c0.n12_adj_4526 ));
    Odrv4 I__14124 (
            .O(N__68532),
            .I(\c0.n12_adj_4526 ));
    InMux I__14123 (
            .O(N__68523),
            .I(N__68520));
    LocalMux I__14122 (
            .O(N__68520),
            .I(N__68516));
    CascadeMux I__14121 (
            .O(N__68519),
            .I(N__68511));
    Span4Mux_h I__14120 (
            .O(N__68516),
            .I(N__68508));
    InMux I__14119 (
            .O(N__68515),
            .I(N__68505));
    InMux I__14118 (
            .O(N__68514),
            .I(N__68502));
    InMux I__14117 (
            .O(N__68511),
            .I(N__68499));
    Span4Mux_h I__14116 (
            .O(N__68508),
            .I(N__68496));
    LocalMux I__14115 (
            .O(N__68505),
            .I(N__68491));
    LocalMux I__14114 (
            .O(N__68502),
            .I(N__68491));
    LocalMux I__14113 (
            .O(N__68499),
            .I(\c0.data_in_frame_13_4 ));
    Odrv4 I__14112 (
            .O(N__68496),
            .I(\c0.data_in_frame_13_4 ));
    Odrv12 I__14111 (
            .O(N__68491),
            .I(\c0.data_in_frame_13_4 ));
    InMux I__14110 (
            .O(N__68484),
            .I(N__68481));
    LocalMux I__14109 (
            .O(N__68481),
            .I(N__68478));
    Odrv4 I__14108 (
            .O(N__68478),
            .I(n2330));
    CascadeMux I__14107 (
            .O(N__68475),
            .I(N__68470));
    InMux I__14106 (
            .O(N__68474),
            .I(N__68467));
    InMux I__14105 (
            .O(N__68473),
            .I(N__68464));
    InMux I__14104 (
            .O(N__68470),
            .I(N__68461));
    LocalMux I__14103 (
            .O(N__68467),
            .I(N__68458));
    LocalMux I__14102 (
            .O(N__68464),
            .I(N__68455));
    LocalMux I__14101 (
            .O(N__68461),
            .I(N__68448));
    Span4Mux_h I__14100 (
            .O(N__68458),
            .I(N__68448));
    Span4Mux_v I__14099 (
            .O(N__68455),
            .I(N__68448));
    Odrv4 I__14098 (
            .O(N__68448),
            .I(\c0.data_in_frame_24_2 ));
    InMux I__14097 (
            .O(N__68445),
            .I(N__68442));
    LocalMux I__14096 (
            .O(N__68442),
            .I(N__68439));
    Span4Mux_h I__14095 (
            .O(N__68439),
            .I(N__68436));
    Odrv4 I__14094 (
            .O(N__68436),
            .I(n2335));
    InMux I__14093 (
            .O(N__68433),
            .I(N__68430));
    LocalMux I__14092 (
            .O(N__68430),
            .I(N__68427));
    Span4Mux_h I__14091 (
            .O(N__68427),
            .I(N__68424));
    Odrv4 I__14090 (
            .O(N__68424),
            .I(n2337));
    InMux I__14089 (
            .O(N__68421),
            .I(N__68415));
    InMux I__14088 (
            .O(N__68420),
            .I(N__68415));
    LocalMux I__14087 (
            .O(N__68415),
            .I(data_out_frame_8_4));
    InMux I__14086 (
            .O(N__68412),
            .I(N__68409));
    LocalMux I__14085 (
            .O(N__68409),
            .I(N__68406));
    Span4Mux_h I__14084 (
            .O(N__68406),
            .I(N__68403));
    Odrv4 I__14083 (
            .O(N__68403),
            .I(\c0.n35812 ));
    InMux I__14082 (
            .O(N__68400),
            .I(N__68396));
    InMux I__14081 (
            .O(N__68399),
            .I(N__68393));
    LocalMux I__14080 (
            .O(N__68396),
            .I(data_out_frame_9_4));
    LocalMux I__14079 (
            .O(N__68393),
            .I(data_out_frame_9_4));
    InMux I__14078 (
            .O(N__68388),
            .I(N__68384));
    InMux I__14077 (
            .O(N__68387),
            .I(N__68381));
    LocalMux I__14076 (
            .O(N__68384),
            .I(data_out_frame_6_4));
    LocalMux I__14075 (
            .O(N__68381),
            .I(data_out_frame_6_4));
    InMux I__14074 (
            .O(N__68376),
            .I(N__68373));
    LocalMux I__14073 (
            .O(N__68373),
            .I(N__68370));
    Odrv4 I__14072 (
            .O(N__68370),
            .I(n2344));
    InMux I__14071 (
            .O(N__68367),
            .I(N__68363));
    InMux I__14070 (
            .O(N__68366),
            .I(N__68360));
    LocalMux I__14069 (
            .O(N__68363),
            .I(data_out_frame_13_4));
    LocalMux I__14068 (
            .O(N__68360),
            .I(data_out_frame_13_4));
    InMux I__14067 (
            .O(N__68355),
            .I(N__68352));
    LocalMux I__14066 (
            .O(N__68352),
            .I(N__68349));
    Span4Mux_v I__14065 (
            .O(N__68349),
            .I(N__68346));
    Odrv4 I__14064 (
            .O(N__68346),
            .I(n2327));
    InMux I__14063 (
            .O(N__68343),
            .I(N__68340));
    LocalMux I__14062 (
            .O(N__68340),
            .I(N__68337));
    Span12Mux_h I__14061 (
            .O(N__68337),
            .I(N__68334));
    Odrv12 I__14060 (
            .O(N__68334),
            .I(n2314));
    InMux I__14059 (
            .O(N__68331),
            .I(N__68328));
    LocalMux I__14058 (
            .O(N__68328),
            .I(N__68325));
    Odrv4 I__14057 (
            .O(N__68325),
            .I(n2338));
    InMux I__14056 (
            .O(N__68322),
            .I(N__68319));
    LocalMux I__14055 (
            .O(N__68319),
            .I(N__68316));
    Span4Mux_h I__14054 (
            .O(N__68316),
            .I(N__68313));
    Span4Mux_v I__14053 (
            .O(N__68313),
            .I(N__68310));
    Odrv4 I__14052 (
            .O(N__68310),
            .I(\c0.n35140 ));
    InMux I__14051 (
            .O(N__68307),
            .I(N__68298));
    InMux I__14050 (
            .O(N__68306),
            .I(N__68298));
    InMux I__14049 (
            .O(N__68305),
            .I(N__68293));
    InMux I__14048 (
            .O(N__68304),
            .I(N__68290));
    InMux I__14047 (
            .O(N__68303),
            .I(N__68287));
    LocalMux I__14046 (
            .O(N__68298),
            .I(N__68284));
    InMux I__14045 (
            .O(N__68297),
            .I(N__68281));
    CascadeMux I__14044 (
            .O(N__68296),
            .I(N__68278));
    LocalMux I__14043 (
            .O(N__68293),
            .I(N__68273));
    LocalMux I__14042 (
            .O(N__68290),
            .I(N__68273));
    LocalMux I__14041 (
            .O(N__68287),
            .I(N__68269));
    Span4Mux_h I__14040 (
            .O(N__68284),
            .I(N__68266));
    LocalMux I__14039 (
            .O(N__68281),
            .I(N__68262));
    InMux I__14038 (
            .O(N__68278),
            .I(N__68259));
    Span4Mux_v I__14037 (
            .O(N__68273),
            .I(N__68256));
    InMux I__14036 (
            .O(N__68272),
            .I(N__68253));
    Span4Mux_v I__14035 (
            .O(N__68269),
            .I(N__68248));
    Span4Mux_h I__14034 (
            .O(N__68266),
            .I(N__68248));
    InMux I__14033 (
            .O(N__68265),
            .I(N__68245));
    Span12Mux_v I__14032 (
            .O(N__68262),
            .I(N__68242));
    LocalMux I__14031 (
            .O(N__68259),
            .I(N__68235));
    Span4Mux_h I__14030 (
            .O(N__68256),
            .I(N__68235));
    LocalMux I__14029 (
            .O(N__68253),
            .I(N__68235));
    Span4Mux_v I__14028 (
            .O(N__68248),
            .I(N__68232));
    LocalMux I__14027 (
            .O(N__68245),
            .I(N__68227));
    Span12Mux_h I__14026 (
            .O(N__68242),
            .I(N__68227));
    Span4Mux_v I__14025 (
            .O(N__68235),
            .I(N__68224));
    Odrv4 I__14024 (
            .O(N__68232),
            .I(\c0.n12_adj_4536 ));
    Odrv12 I__14023 (
            .O(N__68227),
            .I(\c0.n12_adj_4536 ));
    Odrv4 I__14022 (
            .O(N__68224),
            .I(\c0.n12_adj_4536 ));
    InMux I__14021 (
            .O(N__68217),
            .I(N__68214));
    LocalMux I__14020 (
            .O(N__68214),
            .I(N__68210));
    CascadeMux I__14019 (
            .O(N__68213),
            .I(N__68207));
    Span4Mux_h I__14018 (
            .O(N__68210),
            .I(N__68204));
    InMux I__14017 (
            .O(N__68207),
            .I(N__68201));
    Span4Mux_h I__14016 (
            .O(N__68204),
            .I(N__68198));
    LocalMux I__14015 (
            .O(N__68201),
            .I(\c0.data_in_frame_5_4 ));
    Odrv4 I__14014 (
            .O(N__68198),
            .I(\c0.data_in_frame_5_4 ));
    InMux I__14013 (
            .O(N__68193),
            .I(N__68190));
    LocalMux I__14012 (
            .O(N__68190),
            .I(N__68187));
    Odrv12 I__14011 (
            .O(N__68187),
            .I(n2332));
    CascadeMux I__14010 (
            .O(N__68184),
            .I(N__68180));
    CascadeMux I__14009 (
            .O(N__68183),
            .I(N__68177));
    InMux I__14008 (
            .O(N__68180),
            .I(N__68174));
    InMux I__14007 (
            .O(N__68177),
            .I(N__68171));
    LocalMux I__14006 (
            .O(N__68174),
            .I(N__68165));
    LocalMux I__14005 (
            .O(N__68171),
            .I(N__68162));
    InMux I__14004 (
            .O(N__68170),
            .I(N__68159));
    InMux I__14003 (
            .O(N__68169),
            .I(N__68156));
    InMux I__14002 (
            .O(N__68168),
            .I(N__68153));
    Span4Mux_h I__14001 (
            .O(N__68165),
            .I(N__68150));
    Sp12to4 I__14000 (
            .O(N__68162),
            .I(N__68145));
    LocalMux I__13999 (
            .O(N__68159),
            .I(N__68145));
    LocalMux I__13998 (
            .O(N__68156),
            .I(N__68142));
    LocalMux I__13997 (
            .O(N__68153),
            .I(encoder1_position_15));
    Odrv4 I__13996 (
            .O(N__68150),
            .I(encoder1_position_15));
    Odrv12 I__13995 (
            .O(N__68145),
            .I(encoder1_position_15));
    Odrv4 I__13994 (
            .O(N__68142),
            .I(encoder1_position_15));
    InMux I__13993 (
            .O(N__68133),
            .I(N__68130));
    LocalMux I__13992 (
            .O(N__68130),
            .I(\c0.n11_adj_4576 ));
    InMux I__13991 (
            .O(N__68127),
            .I(N__68121));
    InMux I__13990 (
            .O(N__68126),
            .I(N__68121));
    LocalMux I__13989 (
            .O(N__68121),
            .I(data_out_frame_12_4));
    InMux I__13988 (
            .O(N__68118),
            .I(N__68115));
    LocalMux I__13987 (
            .O(N__68115),
            .I(N__68112));
    Span4Mux_h I__13986 (
            .O(N__68112),
            .I(N__68108));
    InMux I__13985 (
            .O(N__68111),
            .I(N__68105));
    Span4Mux_v I__13984 (
            .O(N__68108),
            .I(N__68102));
    LocalMux I__13983 (
            .O(N__68105),
            .I(data_out_frame_5_3));
    Odrv4 I__13982 (
            .O(N__68102),
            .I(data_out_frame_5_3));
    InMux I__13981 (
            .O(N__68097),
            .I(N__68094));
    LocalMux I__13980 (
            .O(N__68094),
            .I(N__68089));
    InMux I__13979 (
            .O(N__68093),
            .I(N__68086));
    InMux I__13978 (
            .O(N__68092),
            .I(N__68083));
    Span4Mux_h I__13977 (
            .O(N__68089),
            .I(N__68080));
    LocalMux I__13976 (
            .O(N__68086),
            .I(N__68074));
    LocalMux I__13975 (
            .O(N__68083),
            .I(N__68074));
    Span4Mux_h I__13974 (
            .O(N__68080),
            .I(N__68069));
    InMux I__13973 (
            .O(N__68079),
            .I(N__68066));
    Span4Mux_h I__13972 (
            .O(N__68074),
            .I(N__68063));
    InMux I__13971 (
            .O(N__68073),
            .I(N__68058));
    InMux I__13970 (
            .O(N__68072),
            .I(N__68058));
    Odrv4 I__13969 (
            .O(N__68069),
            .I(data_in_frame_1_1));
    LocalMux I__13968 (
            .O(N__68066),
            .I(data_in_frame_1_1));
    Odrv4 I__13967 (
            .O(N__68063),
            .I(data_in_frame_1_1));
    LocalMux I__13966 (
            .O(N__68058),
            .I(data_in_frame_1_1));
    InMux I__13965 (
            .O(N__68049),
            .I(N__68045));
    InMux I__13964 (
            .O(N__68048),
            .I(N__68042));
    LocalMux I__13963 (
            .O(N__68045),
            .I(data_out_frame_5_4));
    LocalMux I__13962 (
            .O(N__68042),
            .I(data_out_frame_5_4));
    CascadeMux I__13961 (
            .O(N__68037),
            .I(N__68034));
    InMux I__13960 (
            .O(N__68034),
            .I(N__68031));
    LocalMux I__13959 (
            .O(N__68031),
            .I(N__68025));
    InMux I__13958 (
            .O(N__68030),
            .I(N__68022));
    InMux I__13957 (
            .O(N__68029),
            .I(N__68019));
    InMux I__13956 (
            .O(N__68028),
            .I(N__68015));
    Span4Mux_v I__13955 (
            .O(N__68025),
            .I(N__68010));
    LocalMux I__13954 (
            .O(N__68022),
            .I(N__68010));
    LocalMux I__13953 (
            .O(N__68019),
            .I(N__68007));
    InMux I__13952 (
            .O(N__68018),
            .I(N__68004));
    LocalMux I__13951 (
            .O(N__68015),
            .I(encoder1_position_24));
    Odrv4 I__13950 (
            .O(N__68010),
            .I(encoder1_position_24));
    Odrv4 I__13949 (
            .O(N__68007),
            .I(encoder1_position_24));
    LocalMux I__13948 (
            .O(N__68004),
            .I(encoder1_position_24));
    InMux I__13947 (
            .O(N__67995),
            .I(N__67991));
    InMux I__13946 (
            .O(N__67994),
            .I(N__67988));
    LocalMux I__13945 (
            .O(N__67991),
            .I(N__67985));
    LocalMux I__13944 (
            .O(N__67988),
            .I(data_out_frame_12_5));
    Odrv12 I__13943 (
            .O(N__67985),
            .I(data_out_frame_12_5));
    InMux I__13942 (
            .O(N__67980),
            .I(N__67977));
    LocalMux I__13941 (
            .O(N__67977),
            .I(N__67974));
    Odrv12 I__13940 (
            .O(N__67974),
            .I(\c0.n11_adj_4621 ));
    InMux I__13939 (
            .O(N__67971),
            .I(N__67965));
    InMux I__13938 (
            .O(N__67970),
            .I(N__67965));
    LocalMux I__13937 (
            .O(N__67965),
            .I(data_out_frame_13_5));
    InMux I__13936 (
            .O(N__67962),
            .I(N__67959));
    LocalMux I__13935 (
            .O(N__67959),
            .I(n2250));
    InMux I__13934 (
            .O(N__67956),
            .I(N__67953));
    LocalMux I__13933 (
            .O(N__67953),
            .I(\c0.n43_adj_4569 ));
    InMux I__13932 (
            .O(N__67950),
            .I(N__67947));
    LocalMux I__13931 (
            .O(N__67947),
            .I(n2254));
    InMux I__13930 (
            .O(N__67944),
            .I(N__67941));
    LocalMux I__13929 (
            .O(N__67941),
            .I(N__67933));
    InMux I__13928 (
            .O(N__67940),
            .I(N__67930));
    InMux I__13927 (
            .O(N__67939),
            .I(N__67925));
    InMux I__13926 (
            .O(N__67938),
            .I(N__67925));
    InMux I__13925 (
            .O(N__67937),
            .I(N__67922));
    CascadeMux I__13924 (
            .O(N__67936),
            .I(N__67919));
    Span4Mux_v I__13923 (
            .O(N__67933),
            .I(N__67914));
    LocalMux I__13922 (
            .O(N__67930),
            .I(N__67914));
    LocalMux I__13921 (
            .O(N__67925),
            .I(N__67909));
    LocalMux I__13920 (
            .O(N__67922),
            .I(N__67909));
    InMux I__13919 (
            .O(N__67919),
            .I(N__67906));
    Span4Mux_v I__13918 (
            .O(N__67914),
            .I(N__67903));
    Span12Mux_v I__13917 (
            .O(N__67909),
            .I(N__67900));
    LocalMux I__13916 (
            .O(N__67906),
            .I(\c0.data_in_frame_21_5 ));
    Odrv4 I__13915 (
            .O(N__67903),
            .I(\c0.data_in_frame_21_5 ));
    Odrv12 I__13914 (
            .O(N__67900),
            .I(\c0.data_in_frame_21_5 ));
    InMux I__13913 (
            .O(N__67893),
            .I(N__67890));
    LocalMux I__13912 (
            .O(N__67890),
            .I(N__67886));
    InMux I__13911 (
            .O(N__67889),
            .I(N__67883));
    Span4Mux_h I__13910 (
            .O(N__67886),
            .I(N__67880));
    LocalMux I__13909 (
            .O(N__67883),
            .I(\c0.data_in_frame_5_1 ));
    Odrv4 I__13908 (
            .O(N__67880),
            .I(\c0.data_in_frame_5_1 ));
    CascadeMux I__13907 (
            .O(N__67875),
            .I(N__67872));
    InMux I__13906 (
            .O(N__67872),
            .I(N__67867));
    CascadeMux I__13905 (
            .O(N__67871),
            .I(N__67863));
    CascadeMux I__13904 (
            .O(N__67870),
            .I(N__67860));
    LocalMux I__13903 (
            .O(N__67867),
            .I(N__67857));
    InMux I__13902 (
            .O(N__67866),
            .I(N__67852));
    InMux I__13901 (
            .O(N__67863),
            .I(N__67852));
    InMux I__13900 (
            .O(N__67860),
            .I(N__67849));
    Span4Mux_v I__13899 (
            .O(N__67857),
            .I(N__67846));
    LocalMux I__13898 (
            .O(N__67852),
            .I(encoder1_position_23));
    LocalMux I__13897 (
            .O(N__67849),
            .I(encoder1_position_23));
    Odrv4 I__13896 (
            .O(N__67846),
            .I(encoder1_position_23));
    CascadeMux I__13895 (
            .O(N__67839),
            .I(N__67835));
    InMux I__13894 (
            .O(N__67838),
            .I(N__67830));
    InMux I__13893 (
            .O(N__67835),
            .I(N__67830));
    LocalMux I__13892 (
            .O(N__67830),
            .I(N__67827));
    Odrv4 I__13891 (
            .O(N__67827),
            .I(\c0.n33400 ));
    InMux I__13890 (
            .O(N__67824),
            .I(N__67821));
    LocalMux I__13889 (
            .O(N__67821),
            .I(N__67818));
    Odrv4 I__13888 (
            .O(N__67818),
            .I(n2261));
    CascadeMux I__13887 (
            .O(N__67815),
            .I(N__67811));
    InMux I__13886 (
            .O(N__67814),
            .I(N__67808));
    InMux I__13885 (
            .O(N__67811),
            .I(N__67805));
    LocalMux I__13884 (
            .O(N__67808),
            .I(N__67802));
    LocalMux I__13883 (
            .O(N__67805),
            .I(N__67799));
    Span4Mux_h I__13882 (
            .O(N__67802),
            .I(N__67793));
    Span4Mux_h I__13881 (
            .O(N__67799),
            .I(N__67793));
    CascadeMux I__13880 (
            .O(N__67798),
            .I(N__67790));
    Span4Mux_v I__13879 (
            .O(N__67793),
            .I(N__67785));
    InMux I__13878 (
            .O(N__67790),
            .I(N__67782));
    InMux I__13877 (
            .O(N__67789),
            .I(N__67777));
    InMux I__13876 (
            .O(N__67788),
            .I(N__67777));
    Odrv4 I__13875 (
            .O(N__67785),
            .I(encoder1_position_25));
    LocalMux I__13874 (
            .O(N__67782),
            .I(encoder1_position_25));
    LocalMux I__13873 (
            .O(N__67777),
            .I(encoder1_position_25));
    CascadeMux I__13872 (
            .O(N__67770),
            .I(\c0.n18357_cascade_ ));
    CascadeMux I__13871 (
            .O(N__67767),
            .I(N__67764));
    InMux I__13870 (
            .O(N__67764),
            .I(N__67760));
    InMux I__13869 (
            .O(N__67763),
            .I(N__67757));
    LocalMux I__13868 (
            .O(N__67760),
            .I(N__67754));
    LocalMux I__13867 (
            .O(N__67757),
            .I(data_out_frame_10_7));
    Odrv4 I__13866 (
            .O(N__67754),
            .I(data_out_frame_10_7));
    InMux I__13865 (
            .O(N__67749),
            .I(N__67746));
    LocalMux I__13864 (
            .O(N__67746),
            .I(n2263));
    InMux I__13863 (
            .O(N__67743),
            .I(N__67740));
    LocalMux I__13862 (
            .O(N__67740),
            .I(n2265));
    InMux I__13861 (
            .O(N__67737),
            .I(N__67734));
    LocalMux I__13860 (
            .O(N__67734),
            .I(n2258));
    CascadeMux I__13859 (
            .O(N__67731),
            .I(\c0.n18689_cascade_ ));
    CascadeMux I__13858 (
            .O(N__67728),
            .I(\c0.n38_adj_4568_cascade_ ));
    CascadeMux I__13857 (
            .O(N__67725),
            .I(\c0.n36179_cascade_ ));
    InMux I__13856 (
            .O(N__67722),
            .I(N__67719));
    LocalMux I__13855 (
            .O(N__67719),
            .I(N__67716));
    Span4Mux_v I__13854 (
            .O(N__67716),
            .I(N__67712));
    InMux I__13853 (
            .O(N__67715),
            .I(N__67709));
    Span4Mux_h I__13852 (
            .O(N__67712),
            .I(N__67706));
    LocalMux I__13851 (
            .O(N__67709),
            .I(data_out_frame_9_5));
    Odrv4 I__13850 (
            .O(N__67706),
            .I(data_out_frame_9_5));
    CascadeMux I__13849 (
            .O(N__67701),
            .I(\c0.n36182_cascade_ ));
    CascadeMux I__13848 (
            .O(N__67698),
            .I(n36098_cascade_));
    InMux I__13847 (
            .O(N__67695),
            .I(N__67692));
    LocalMux I__13846 (
            .O(N__67692),
            .I(n2270));
    InMux I__13845 (
            .O(N__67689),
            .I(N__67686));
    LocalMux I__13844 (
            .O(N__67686),
            .I(n2268));
    InMux I__13843 (
            .O(N__67683),
            .I(N__67680));
    LocalMux I__13842 (
            .O(N__67680),
            .I(n2266));
    CascadeMux I__13841 (
            .O(N__67677),
            .I(N__67674));
    InMux I__13840 (
            .O(N__67674),
            .I(N__67670));
    InMux I__13839 (
            .O(N__67673),
            .I(N__67667));
    LocalMux I__13838 (
            .O(N__67670),
            .I(data_out_frame_8_5));
    LocalMux I__13837 (
            .O(N__67667),
            .I(data_out_frame_8_5));
    InMux I__13836 (
            .O(N__67662),
            .I(N__67659));
    LocalMux I__13835 (
            .O(N__67659),
            .I(N__67656));
    Odrv12 I__13834 (
            .O(N__67656),
            .I(\quad_counter1.n28_adj_4488 ));
    CascadeMux I__13833 (
            .O(N__67653),
            .I(N__67639));
    CascadeMux I__13832 (
            .O(N__67652),
            .I(N__67636));
    CascadeMux I__13831 (
            .O(N__67651),
            .I(N__67630));
    CascadeMux I__13830 (
            .O(N__67650),
            .I(N__67627));
    CascadeMux I__13829 (
            .O(N__67649),
            .I(N__67624));
    CascadeMux I__13828 (
            .O(N__67648),
            .I(N__67621));
    CascadeMux I__13827 (
            .O(N__67647),
            .I(N__67618));
    CascadeMux I__13826 (
            .O(N__67646),
            .I(N__67615));
    CascadeMux I__13825 (
            .O(N__67645),
            .I(N__67612));
    CascadeMux I__13824 (
            .O(N__67644),
            .I(N__67609));
    CascadeMux I__13823 (
            .O(N__67643),
            .I(N__67606));
    CascadeMux I__13822 (
            .O(N__67642),
            .I(N__67603));
    InMux I__13821 (
            .O(N__67639),
            .I(N__67598));
    InMux I__13820 (
            .O(N__67636),
            .I(N__67598));
    CascadeMux I__13819 (
            .O(N__67635),
            .I(N__67595));
    CascadeMux I__13818 (
            .O(N__67634),
            .I(N__67592));
    CascadeMux I__13817 (
            .O(N__67633),
            .I(N__67589));
    InMux I__13816 (
            .O(N__67630),
            .I(N__67583));
    InMux I__13815 (
            .O(N__67627),
            .I(N__67583));
    InMux I__13814 (
            .O(N__67624),
            .I(N__67574));
    InMux I__13813 (
            .O(N__67621),
            .I(N__67574));
    InMux I__13812 (
            .O(N__67618),
            .I(N__67574));
    InMux I__13811 (
            .O(N__67615),
            .I(N__67574));
    InMux I__13810 (
            .O(N__67612),
            .I(N__67565));
    InMux I__13809 (
            .O(N__67609),
            .I(N__67565));
    InMux I__13808 (
            .O(N__67606),
            .I(N__67565));
    InMux I__13807 (
            .O(N__67603),
            .I(N__67565));
    LocalMux I__13806 (
            .O(N__67598),
            .I(N__67562));
    InMux I__13805 (
            .O(N__67595),
            .I(N__67553));
    InMux I__13804 (
            .O(N__67592),
            .I(N__67553));
    InMux I__13803 (
            .O(N__67589),
            .I(N__67553));
    InMux I__13802 (
            .O(N__67588),
            .I(N__67553));
    LocalMux I__13801 (
            .O(N__67583),
            .I(\quad_counter1.n3233 ));
    LocalMux I__13800 (
            .O(N__67574),
            .I(\quad_counter1.n3233 ));
    LocalMux I__13799 (
            .O(N__67565),
            .I(\quad_counter1.n3233 ));
    Odrv4 I__13798 (
            .O(N__67562),
            .I(\quad_counter1.n3233 ));
    LocalMux I__13797 (
            .O(N__67553),
            .I(\quad_counter1.n3233 ));
    InMux I__13796 (
            .O(N__67542),
            .I(N__67539));
    LocalMux I__13795 (
            .O(N__67539),
            .I(n2278));
    InMux I__13794 (
            .O(N__67536),
            .I(N__67532));
    InMux I__13793 (
            .O(N__67535),
            .I(N__67529));
    LocalMux I__13792 (
            .O(N__67532),
            .I(data_out_frame_12_3));
    LocalMux I__13791 (
            .O(N__67529),
            .I(data_out_frame_12_3));
    InMux I__13790 (
            .O(N__67524),
            .I(N__67521));
    LocalMux I__13789 (
            .O(N__67521),
            .I(N__67518));
    Span4Mux_v I__13788 (
            .O(N__67518),
            .I(N__67515));
    Span4Mux_h I__13787 (
            .O(N__67515),
            .I(N__67512));
    Odrv4 I__13786 (
            .O(N__67512),
            .I(\c0.n11_adj_4517 ));
    InMux I__13785 (
            .O(N__67509),
            .I(N__67506));
    LocalMux I__13784 (
            .O(N__67506),
            .I(N__67503));
    Odrv4 I__13783 (
            .O(N__67503),
            .I(n2264));
    InMux I__13782 (
            .O(N__67500),
            .I(N__67497));
    LocalMux I__13781 (
            .O(N__67497),
            .I(n2276));
    InMux I__13780 (
            .O(N__67494),
            .I(N__67491));
    LocalMux I__13779 (
            .O(N__67491),
            .I(N__67488));
    Span4Mux_v I__13778 (
            .O(N__67488),
            .I(N__67485));
    Span4Mux_h I__13777 (
            .O(N__67485),
            .I(N__67482));
    Odrv4 I__13776 (
            .O(N__67482),
            .I(\c0.n11_adj_4507 ));
    InMux I__13775 (
            .O(N__67479),
            .I(N__67473));
    InMux I__13774 (
            .O(N__67478),
            .I(N__67473));
    LocalMux I__13773 (
            .O(N__67473),
            .I(data_out_frame_12_1));
    InMux I__13772 (
            .O(N__67470),
            .I(N__67467));
    LocalMux I__13771 (
            .O(N__67467),
            .I(N__67464));
    Sp12to4 I__13770 (
            .O(N__67464),
            .I(N__67460));
    InMux I__13769 (
            .O(N__67463),
            .I(N__67457));
    Span12Mux_h I__13768 (
            .O(N__67460),
            .I(N__67454));
    LocalMux I__13767 (
            .O(N__67457),
            .I(data_out_frame_11_5));
    Odrv12 I__13766 (
            .O(N__67454),
            .I(data_out_frame_11_5));
    InMux I__13765 (
            .O(N__67449),
            .I(\quad_counter1.n30647 ));
    InMux I__13764 (
            .O(N__67446),
            .I(\quad_counter1.n30648 ));
    InMux I__13763 (
            .O(N__67443),
            .I(bfn_19_13_0_));
    InMux I__13762 (
            .O(N__67440),
            .I(\quad_counter1.n30650 ));
    InMux I__13761 (
            .O(N__67437),
            .I(\quad_counter1.n30651 ));
    InMux I__13760 (
            .O(N__67434),
            .I(\quad_counter1.n30652 ));
    InMux I__13759 (
            .O(N__67431),
            .I(\quad_counter1.n30653 ));
    CascadeMux I__13758 (
            .O(N__67428),
            .I(N__67420));
    CascadeMux I__13757 (
            .O(N__67427),
            .I(N__67417));
    CascadeMux I__13756 (
            .O(N__67426),
            .I(N__67414));
    CascadeMux I__13755 (
            .O(N__67425),
            .I(N__67411));
    CascadeMux I__13754 (
            .O(N__67424),
            .I(N__67408));
    CascadeMux I__13753 (
            .O(N__67423),
            .I(N__67405));
    InMux I__13752 (
            .O(N__67420),
            .I(N__67400));
    InMux I__13751 (
            .O(N__67417),
            .I(N__67400));
    InMux I__13750 (
            .O(N__67414),
            .I(N__67391));
    InMux I__13749 (
            .O(N__67411),
            .I(N__67391));
    InMux I__13748 (
            .O(N__67408),
            .I(N__67391));
    InMux I__13747 (
            .O(N__67405),
            .I(N__67391));
    LocalMux I__13746 (
            .O(N__67400),
            .I(N__67386));
    LocalMux I__13745 (
            .O(N__67391),
            .I(N__67386));
    Odrv4 I__13744 (
            .O(N__67386),
            .I(\quad_counter1.n36148 ));
    InMux I__13743 (
            .O(N__67383),
            .I(N__67380));
    LocalMux I__13742 (
            .O(N__67380),
            .I(N__67377));
    Odrv12 I__13741 (
            .O(N__67377),
            .I(\quad_counter1.n24_adj_4487 ));
    CascadeMux I__13740 (
            .O(N__67374),
            .I(N__67371));
    InMux I__13739 (
            .O(N__67371),
            .I(N__67368));
    LocalMux I__13738 (
            .O(N__67368),
            .I(N__67365));
    Odrv12 I__13737 (
            .O(N__67365),
            .I(\quad_counter1.n16_adj_4486 ));
    InMux I__13736 (
            .O(N__67362),
            .I(\quad_counter1.n30637 ));
    InMux I__13735 (
            .O(N__67359),
            .I(\quad_counter1.n30638 ));
    InMux I__13734 (
            .O(N__67356),
            .I(\quad_counter1.n30639 ));
    InMux I__13733 (
            .O(N__67353),
            .I(\quad_counter1.n30640 ));
    InMux I__13732 (
            .O(N__67350),
            .I(bfn_19_12_0_));
    InMux I__13731 (
            .O(N__67347),
            .I(\quad_counter1.n30642 ));
    InMux I__13730 (
            .O(N__67344),
            .I(\quad_counter1.n30643 ));
    InMux I__13729 (
            .O(N__67341),
            .I(\quad_counter1.n30644 ));
    InMux I__13728 (
            .O(N__67338),
            .I(\quad_counter1.n30645 ));
    InMux I__13727 (
            .O(N__67335),
            .I(\quad_counter1.n30646 ));
    InMux I__13726 (
            .O(N__67332),
            .I(N__67329));
    LocalMux I__13725 (
            .O(N__67329),
            .I(\quad_counter1.n19_adj_4485 ));
    CascadeMux I__13724 (
            .O(N__67326),
            .I(\quad_counter1.n26_adj_4484_cascade_ ));
    InMux I__13723 (
            .O(N__67323),
            .I(bfn_19_11_0_));
    InMux I__13722 (
            .O(N__67320),
            .I(\quad_counter1.n30634 ));
    InMux I__13721 (
            .O(N__67317),
            .I(\quad_counter1.n30635 ));
    InMux I__13720 (
            .O(N__67314),
            .I(\quad_counter1.n30636 ));
    InMux I__13719 (
            .O(N__67311),
            .I(N__67306));
    InMux I__13718 (
            .O(N__67310),
            .I(N__67303));
    CascadeMux I__13717 (
            .O(N__67309),
            .I(N__67300));
    LocalMux I__13716 (
            .O(N__67306),
            .I(N__67295));
    LocalMux I__13715 (
            .O(N__67303),
            .I(N__67295));
    InMux I__13714 (
            .O(N__67300),
            .I(N__67292));
    Odrv4 I__13713 (
            .O(N__67295),
            .I(\quad_counter1.n3006 ));
    LocalMux I__13712 (
            .O(N__67292),
            .I(\quad_counter1.n3006 ));
    InMux I__13711 (
            .O(N__67287),
            .I(\quad_counter1.n30610 ));
    InMux I__13710 (
            .O(N__67284),
            .I(N__67279));
    InMux I__13709 (
            .O(N__67283),
            .I(N__67276));
    CascadeMux I__13708 (
            .O(N__67282),
            .I(N__67273));
    LocalMux I__13707 (
            .O(N__67279),
            .I(N__67268));
    LocalMux I__13706 (
            .O(N__67276),
            .I(N__67268));
    InMux I__13705 (
            .O(N__67273),
            .I(N__67265));
    Odrv4 I__13704 (
            .O(N__67268),
            .I(\quad_counter1.n3005 ));
    LocalMux I__13703 (
            .O(N__67265),
            .I(\quad_counter1.n3005 ));
    InMux I__13702 (
            .O(N__67260),
            .I(\quad_counter1.n30611 ));
    InMux I__13701 (
            .O(N__67257),
            .I(N__67253));
    InMux I__13700 (
            .O(N__67256),
            .I(N__67250));
    LocalMux I__13699 (
            .O(N__67253),
            .I(N__67245));
    LocalMux I__13698 (
            .O(N__67250),
            .I(N__67245));
    Span4Mux_h I__13697 (
            .O(N__67245),
            .I(N__67241));
    InMux I__13696 (
            .O(N__67244),
            .I(N__67238));
    Odrv4 I__13695 (
            .O(N__67241),
            .I(\quad_counter1.n3004 ));
    LocalMux I__13694 (
            .O(N__67238),
            .I(\quad_counter1.n3004 ));
    InMux I__13693 (
            .O(N__67233),
            .I(bfn_19_7_0_));
    InMux I__13692 (
            .O(N__67230),
            .I(N__67226));
    InMux I__13691 (
            .O(N__67229),
            .I(N__67223));
    LocalMux I__13690 (
            .O(N__67226),
            .I(N__67217));
    LocalMux I__13689 (
            .O(N__67223),
            .I(N__67217));
    InMux I__13688 (
            .O(N__67222),
            .I(N__67214));
    Odrv4 I__13687 (
            .O(N__67217),
            .I(\quad_counter1.n3003 ));
    LocalMux I__13686 (
            .O(N__67214),
            .I(\quad_counter1.n3003 ));
    InMux I__13685 (
            .O(N__67209),
            .I(\quad_counter1.n30613 ));
    InMux I__13684 (
            .O(N__67206),
            .I(N__67202));
    InMux I__13683 (
            .O(N__67205),
            .I(N__67199));
    LocalMux I__13682 (
            .O(N__67202),
            .I(N__67196));
    LocalMux I__13681 (
            .O(N__67199),
            .I(N__67192));
    Span4Mux_h I__13680 (
            .O(N__67196),
            .I(N__67189));
    InMux I__13679 (
            .O(N__67195),
            .I(N__67186));
    Odrv4 I__13678 (
            .O(N__67192),
            .I(\quad_counter1.n3002 ));
    Odrv4 I__13677 (
            .O(N__67189),
            .I(\quad_counter1.n3002 ));
    LocalMux I__13676 (
            .O(N__67186),
            .I(\quad_counter1.n3002 ));
    CascadeMux I__13675 (
            .O(N__67179),
            .I(N__67164));
    CascadeMux I__13674 (
            .O(N__67178),
            .I(N__67161));
    CascadeMux I__13673 (
            .O(N__67177),
            .I(N__67158));
    CascadeMux I__13672 (
            .O(N__67176),
            .I(N__67155));
    CascadeMux I__13671 (
            .O(N__67175),
            .I(N__67152));
    CascadeMux I__13670 (
            .O(N__67174),
            .I(N__67149));
    CascadeMux I__13669 (
            .O(N__67173),
            .I(N__67146));
    CascadeMux I__13668 (
            .O(N__67172),
            .I(N__67143));
    CascadeMux I__13667 (
            .O(N__67171),
            .I(N__67140));
    CascadeMux I__13666 (
            .O(N__67170),
            .I(N__67137));
    CascadeMux I__13665 (
            .O(N__67169),
            .I(N__67134));
    CascadeMux I__13664 (
            .O(N__67168),
            .I(N__67131));
    CascadeMux I__13663 (
            .O(N__67167),
            .I(N__67128));
    InMux I__13662 (
            .O(N__67164),
            .I(N__67123));
    InMux I__13661 (
            .O(N__67161),
            .I(N__67123));
    InMux I__13660 (
            .O(N__67158),
            .I(N__67120));
    InMux I__13659 (
            .O(N__67155),
            .I(N__67115));
    InMux I__13658 (
            .O(N__67152),
            .I(N__67115));
    InMux I__13657 (
            .O(N__67149),
            .I(N__67106));
    InMux I__13656 (
            .O(N__67146),
            .I(N__67106));
    InMux I__13655 (
            .O(N__67143),
            .I(N__67106));
    InMux I__13654 (
            .O(N__67140),
            .I(N__67106));
    InMux I__13653 (
            .O(N__67137),
            .I(N__67097));
    InMux I__13652 (
            .O(N__67134),
            .I(N__67097));
    InMux I__13651 (
            .O(N__67131),
            .I(N__67097));
    InMux I__13650 (
            .O(N__67128),
            .I(N__67097));
    LocalMux I__13649 (
            .O(N__67123),
            .I(N__67094));
    LocalMux I__13648 (
            .O(N__67120),
            .I(\quad_counter1.n3035 ));
    LocalMux I__13647 (
            .O(N__67115),
            .I(\quad_counter1.n3035 ));
    LocalMux I__13646 (
            .O(N__67106),
            .I(\quad_counter1.n3035 ));
    LocalMux I__13645 (
            .O(N__67097),
            .I(\quad_counter1.n3035 ));
    Odrv4 I__13644 (
            .O(N__67094),
            .I(\quad_counter1.n3035 ));
    InMux I__13643 (
            .O(N__67083),
            .I(\quad_counter1.n30614 ));
    CascadeMux I__13642 (
            .O(N__67080),
            .I(\quad_counter1.n18_adj_4479_cascade_ ));
    InMux I__13641 (
            .O(N__67077),
            .I(N__67074));
    LocalMux I__13640 (
            .O(N__67074),
            .I(\quad_counter1.n24_adj_4480 ));
    InMux I__13639 (
            .O(N__67071),
            .I(N__67067));
    InMux I__13638 (
            .O(N__67070),
            .I(N__67064));
    LocalMux I__13637 (
            .O(N__67067),
            .I(N__67058));
    LocalMux I__13636 (
            .O(N__67064),
            .I(N__67058));
    InMux I__13635 (
            .O(N__67063),
            .I(N__67055));
    Odrv4 I__13634 (
            .O(N__67058),
            .I(\quad_counter1.n3014 ));
    LocalMux I__13633 (
            .O(N__67055),
            .I(\quad_counter1.n3014 ));
    CascadeMux I__13632 (
            .O(N__67050),
            .I(N__67042));
    CascadeMux I__13631 (
            .O(N__67049),
            .I(N__67039));
    CascadeMux I__13630 (
            .O(N__67048),
            .I(N__67036));
    CascadeMux I__13629 (
            .O(N__67047),
            .I(N__67033));
    CascadeMux I__13628 (
            .O(N__67046),
            .I(N__67030));
    CascadeMux I__13627 (
            .O(N__67045),
            .I(N__67027));
    InMux I__13626 (
            .O(N__67042),
            .I(N__67022));
    InMux I__13625 (
            .O(N__67039),
            .I(N__67022));
    InMux I__13624 (
            .O(N__67036),
            .I(N__67013));
    InMux I__13623 (
            .O(N__67033),
            .I(N__67013));
    InMux I__13622 (
            .O(N__67030),
            .I(N__67013));
    InMux I__13621 (
            .O(N__67027),
            .I(N__67013));
    LocalMux I__13620 (
            .O(N__67022),
            .I(\quad_counter1.n36156 ));
    LocalMux I__13619 (
            .O(N__67013),
            .I(\quad_counter1.n36156 ));
    InMux I__13618 (
            .O(N__67008),
            .I(\quad_counter1.n30602 ));
    InMux I__13617 (
            .O(N__67005),
            .I(N__67001));
    InMux I__13616 (
            .O(N__67004),
            .I(N__66998));
    LocalMux I__13615 (
            .O(N__67001),
            .I(N__66992));
    LocalMux I__13614 (
            .O(N__66998),
            .I(N__66992));
    InMux I__13613 (
            .O(N__66997),
            .I(N__66989));
    Span4Mux_v I__13612 (
            .O(N__66992),
            .I(N__66986));
    LocalMux I__13611 (
            .O(N__66989),
            .I(N__66983));
    Odrv4 I__13610 (
            .O(N__66986),
            .I(\quad_counter1.n3013 ));
    Odrv4 I__13609 (
            .O(N__66983),
            .I(\quad_counter1.n3013 ));
    InMux I__13608 (
            .O(N__66978),
            .I(\quad_counter1.n30603 ));
    InMux I__13607 (
            .O(N__66975),
            .I(N__66971));
    InMux I__13606 (
            .O(N__66974),
            .I(N__66968));
    LocalMux I__13605 (
            .O(N__66971),
            .I(N__66962));
    LocalMux I__13604 (
            .O(N__66968),
            .I(N__66962));
    InMux I__13603 (
            .O(N__66967),
            .I(N__66959));
    Odrv4 I__13602 (
            .O(N__66962),
            .I(\quad_counter1.n3012 ));
    LocalMux I__13601 (
            .O(N__66959),
            .I(\quad_counter1.n3012 ));
    InMux I__13600 (
            .O(N__66954),
            .I(bfn_19_6_0_));
    InMux I__13599 (
            .O(N__66951),
            .I(N__66947));
    InMux I__13598 (
            .O(N__66950),
            .I(N__66944));
    LocalMux I__13597 (
            .O(N__66947),
            .I(N__66938));
    LocalMux I__13596 (
            .O(N__66944),
            .I(N__66938));
    InMux I__13595 (
            .O(N__66943),
            .I(N__66935));
    Span4Mux_h I__13594 (
            .O(N__66938),
            .I(N__66930));
    LocalMux I__13593 (
            .O(N__66935),
            .I(N__66930));
    Odrv4 I__13592 (
            .O(N__66930),
            .I(\quad_counter1.n3011 ));
    InMux I__13591 (
            .O(N__66927),
            .I(\quad_counter1.n30605 ));
    InMux I__13590 (
            .O(N__66924),
            .I(N__66920));
    InMux I__13589 (
            .O(N__66923),
            .I(N__66917));
    LocalMux I__13588 (
            .O(N__66920),
            .I(N__66911));
    LocalMux I__13587 (
            .O(N__66917),
            .I(N__66911));
    InMux I__13586 (
            .O(N__66916),
            .I(N__66908));
    Span4Mux_v I__13585 (
            .O(N__66911),
            .I(N__66905));
    LocalMux I__13584 (
            .O(N__66908),
            .I(N__66902));
    Odrv4 I__13583 (
            .O(N__66905),
            .I(\quad_counter1.n3010 ));
    Odrv4 I__13582 (
            .O(N__66902),
            .I(\quad_counter1.n3010 ));
    InMux I__13581 (
            .O(N__66897),
            .I(\quad_counter1.n30606 ));
    InMux I__13580 (
            .O(N__66894),
            .I(N__66889));
    InMux I__13579 (
            .O(N__66893),
            .I(N__66886));
    CascadeMux I__13578 (
            .O(N__66892),
            .I(N__66883));
    LocalMux I__13577 (
            .O(N__66889),
            .I(N__66878));
    LocalMux I__13576 (
            .O(N__66886),
            .I(N__66878));
    InMux I__13575 (
            .O(N__66883),
            .I(N__66875));
    Span4Mux_v I__13574 (
            .O(N__66878),
            .I(N__66872));
    LocalMux I__13573 (
            .O(N__66875),
            .I(N__66869));
    Odrv4 I__13572 (
            .O(N__66872),
            .I(\quad_counter1.n3009 ));
    Odrv4 I__13571 (
            .O(N__66869),
            .I(\quad_counter1.n3009 ));
    InMux I__13570 (
            .O(N__66864),
            .I(\quad_counter1.n30607 ));
    InMux I__13569 (
            .O(N__66861),
            .I(N__66857));
    InMux I__13568 (
            .O(N__66860),
            .I(N__66854));
    LocalMux I__13567 (
            .O(N__66857),
            .I(N__66849));
    LocalMux I__13566 (
            .O(N__66854),
            .I(N__66849));
    Span4Mux_v I__13565 (
            .O(N__66849),
            .I(N__66845));
    InMux I__13564 (
            .O(N__66848),
            .I(N__66842));
    Odrv4 I__13563 (
            .O(N__66845),
            .I(\quad_counter1.n3008 ));
    LocalMux I__13562 (
            .O(N__66842),
            .I(\quad_counter1.n3008 ));
    InMux I__13561 (
            .O(N__66837),
            .I(\quad_counter1.n30608 ));
    InMux I__13560 (
            .O(N__66834),
            .I(N__66830));
    InMux I__13559 (
            .O(N__66833),
            .I(N__66827));
    LocalMux I__13558 (
            .O(N__66830),
            .I(N__66822));
    LocalMux I__13557 (
            .O(N__66827),
            .I(N__66822));
    Span4Mux_v I__13556 (
            .O(N__66822),
            .I(N__66818));
    InMux I__13555 (
            .O(N__66821),
            .I(N__66815));
    Odrv4 I__13554 (
            .O(N__66818),
            .I(\quad_counter1.n3007 ));
    LocalMux I__13553 (
            .O(N__66815),
            .I(\quad_counter1.n3007 ));
    InMux I__13552 (
            .O(N__66810),
            .I(\quad_counter1.n30609 ));
    InMux I__13551 (
            .O(N__66807),
            .I(\quad_counter1.n30577 ));
    InMux I__13550 (
            .O(N__66804),
            .I(N__66801));
    LocalMux I__13549 (
            .O(N__66801),
            .I(N__66796));
    InMux I__13548 (
            .O(N__66800),
            .I(N__66791));
    InMux I__13547 (
            .O(N__66799),
            .I(N__66791));
    Span4Mux_h I__13546 (
            .O(N__66796),
            .I(N__66788));
    LocalMux I__13545 (
            .O(N__66791),
            .I(N__66785));
    Odrv4 I__13544 (
            .O(N__66788),
            .I(\quad_counter1.n2904 ));
    Odrv4 I__13543 (
            .O(N__66785),
            .I(\quad_counter1.n2904 ));
    InMux I__13542 (
            .O(N__66780),
            .I(\quad_counter1.n30578 ));
    InMux I__13541 (
            .O(N__66777),
            .I(bfn_19_4_0_));
    InMux I__13540 (
            .O(N__66774),
            .I(N__66769));
    InMux I__13539 (
            .O(N__66773),
            .I(N__66766));
    InMux I__13538 (
            .O(N__66772),
            .I(N__66763));
    LocalMux I__13537 (
            .O(N__66769),
            .I(N__66760));
    LocalMux I__13536 (
            .O(N__66766),
            .I(\quad_counter1.n2903 ));
    LocalMux I__13535 (
            .O(N__66763),
            .I(\quad_counter1.n2903 ));
    Odrv4 I__13534 (
            .O(N__66760),
            .I(\quad_counter1.n2903 ));
    InMux I__13533 (
            .O(N__66753),
            .I(bfn_19_5_0_));
    InMux I__13532 (
            .O(N__66750),
            .I(N__66746));
    InMux I__13531 (
            .O(N__66749),
            .I(N__66743));
    LocalMux I__13530 (
            .O(N__66746),
            .I(N__66738));
    LocalMux I__13529 (
            .O(N__66743),
            .I(N__66738));
    Span4Mux_v I__13528 (
            .O(N__66738),
            .I(N__66734));
    InMux I__13527 (
            .O(N__66737),
            .I(N__66731));
    Odrv4 I__13526 (
            .O(N__66734),
            .I(\quad_counter1.n3019 ));
    LocalMux I__13525 (
            .O(N__66731),
            .I(\quad_counter1.n3019 ));
    InMux I__13524 (
            .O(N__66726),
            .I(\quad_counter1.n30597 ));
    InMux I__13523 (
            .O(N__66723),
            .I(N__66719));
    InMux I__13522 (
            .O(N__66722),
            .I(N__66716));
    LocalMux I__13521 (
            .O(N__66719),
            .I(N__66711));
    LocalMux I__13520 (
            .O(N__66716),
            .I(N__66711));
    Span4Mux_v I__13519 (
            .O(N__66711),
            .I(N__66707));
    InMux I__13518 (
            .O(N__66710),
            .I(N__66704));
    Odrv4 I__13517 (
            .O(N__66707),
            .I(\quad_counter1.n3018 ));
    LocalMux I__13516 (
            .O(N__66704),
            .I(\quad_counter1.n3018 ));
    InMux I__13515 (
            .O(N__66699),
            .I(\quad_counter1.n30598 ));
    InMux I__13514 (
            .O(N__66696),
            .I(N__66692));
    InMux I__13513 (
            .O(N__66695),
            .I(N__66689));
    LocalMux I__13512 (
            .O(N__66692),
            .I(N__66683));
    LocalMux I__13511 (
            .O(N__66689),
            .I(N__66683));
    InMux I__13510 (
            .O(N__66688),
            .I(N__66680));
    Odrv4 I__13509 (
            .O(N__66683),
            .I(\quad_counter1.n3017 ));
    LocalMux I__13508 (
            .O(N__66680),
            .I(\quad_counter1.n3017 ));
    InMux I__13507 (
            .O(N__66675),
            .I(\quad_counter1.n30599 ));
    InMux I__13506 (
            .O(N__66672),
            .I(N__66668));
    InMux I__13505 (
            .O(N__66671),
            .I(N__66665));
    LocalMux I__13504 (
            .O(N__66668),
            .I(N__66659));
    LocalMux I__13503 (
            .O(N__66665),
            .I(N__66659));
    InMux I__13502 (
            .O(N__66664),
            .I(N__66656));
    Odrv4 I__13501 (
            .O(N__66659),
            .I(\quad_counter1.n3016 ));
    LocalMux I__13500 (
            .O(N__66656),
            .I(\quad_counter1.n3016 ));
    InMux I__13499 (
            .O(N__66651),
            .I(\quad_counter1.n30600 ));
    InMux I__13498 (
            .O(N__66648),
            .I(N__66644));
    InMux I__13497 (
            .O(N__66647),
            .I(N__66641));
    LocalMux I__13496 (
            .O(N__66644),
            .I(N__66635));
    LocalMux I__13495 (
            .O(N__66641),
            .I(N__66635));
    InMux I__13494 (
            .O(N__66640),
            .I(N__66632));
    Odrv4 I__13493 (
            .O(N__66635),
            .I(\quad_counter1.n3015 ));
    LocalMux I__13492 (
            .O(N__66632),
            .I(\quad_counter1.n3015 ));
    InMux I__13491 (
            .O(N__66627),
            .I(\quad_counter1.n30601 ));
    CascadeMux I__13490 (
            .O(N__66624),
            .I(N__66619));
    InMux I__13489 (
            .O(N__66623),
            .I(N__66616));
    InMux I__13488 (
            .O(N__66622),
            .I(N__66613));
    InMux I__13487 (
            .O(N__66619),
            .I(N__66610));
    LocalMux I__13486 (
            .O(N__66616),
            .I(\quad_counter1.n2913 ));
    LocalMux I__13485 (
            .O(N__66613),
            .I(\quad_counter1.n2913 ));
    LocalMux I__13484 (
            .O(N__66610),
            .I(\quad_counter1.n2913 ));
    InMux I__13483 (
            .O(N__66603),
            .I(\quad_counter1.n30569 ));
    InMux I__13482 (
            .O(N__66600),
            .I(N__66597));
    LocalMux I__13481 (
            .O(N__66597),
            .I(N__66594));
    Span4Mux_v I__13480 (
            .O(N__66594),
            .I(N__66590));
    InMux I__13479 (
            .O(N__66593),
            .I(N__66587));
    Span4Mux_s0_v I__13478 (
            .O(N__66590),
            .I(N__66581));
    LocalMux I__13477 (
            .O(N__66587),
            .I(N__66581));
    InMux I__13476 (
            .O(N__66586),
            .I(N__66578));
    Odrv4 I__13475 (
            .O(N__66581),
            .I(\quad_counter1.n2912 ));
    LocalMux I__13474 (
            .O(N__66578),
            .I(\quad_counter1.n2912 ));
    InMux I__13473 (
            .O(N__66573),
            .I(\quad_counter1.n30570 ));
    InMux I__13472 (
            .O(N__66570),
            .I(N__66565));
    InMux I__13471 (
            .O(N__66569),
            .I(N__66562));
    InMux I__13470 (
            .O(N__66568),
            .I(N__66559));
    LocalMux I__13469 (
            .O(N__66565),
            .I(\quad_counter1.n2911 ));
    LocalMux I__13468 (
            .O(N__66562),
            .I(\quad_counter1.n2911 ));
    LocalMux I__13467 (
            .O(N__66559),
            .I(\quad_counter1.n2911 ));
    InMux I__13466 (
            .O(N__66552),
            .I(bfn_19_3_0_));
    InMux I__13465 (
            .O(N__66549),
            .I(N__66544));
    InMux I__13464 (
            .O(N__66548),
            .I(N__66541));
    InMux I__13463 (
            .O(N__66547),
            .I(N__66538));
    LocalMux I__13462 (
            .O(N__66544),
            .I(N__66535));
    LocalMux I__13461 (
            .O(N__66541),
            .I(\quad_counter1.n2910 ));
    LocalMux I__13460 (
            .O(N__66538),
            .I(\quad_counter1.n2910 ));
    Odrv4 I__13459 (
            .O(N__66535),
            .I(\quad_counter1.n2910 ));
    InMux I__13458 (
            .O(N__66528),
            .I(\quad_counter1.n30572 ));
    InMux I__13457 (
            .O(N__66525),
            .I(N__66521));
    InMux I__13456 (
            .O(N__66524),
            .I(N__66517));
    LocalMux I__13455 (
            .O(N__66521),
            .I(N__66514));
    CascadeMux I__13454 (
            .O(N__66520),
            .I(N__66511));
    LocalMux I__13453 (
            .O(N__66517),
            .I(N__66506));
    Span4Mux_h I__13452 (
            .O(N__66514),
            .I(N__66506));
    InMux I__13451 (
            .O(N__66511),
            .I(N__66503));
    Odrv4 I__13450 (
            .O(N__66506),
            .I(\quad_counter1.n2909 ));
    LocalMux I__13449 (
            .O(N__66503),
            .I(\quad_counter1.n2909 ));
    InMux I__13448 (
            .O(N__66498),
            .I(\quad_counter1.n30573 ));
    CascadeMux I__13447 (
            .O(N__66495),
            .I(N__66492));
    InMux I__13446 (
            .O(N__66492),
            .I(N__66487));
    InMux I__13445 (
            .O(N__66491),
            .I(N__66484));
    InMux I__13444 (
            .O(N__66490),
            .I(N__66481));
    LocalMux I__13443 (
            .O(N__66487),
            .I(N__66478));
    LocalMux I__13442 (
            .O(N__66484),
            .I(\quad_counter1.n2908 ));
    LocalMux I__13441 (
            .O(N__66481),
            .I(\quad_counter1.n2908 ));
    Odrv4 I__13440 (
            .O(N__66478),
            .I(\quad_counter1.n2908 ));
    InMux I__13439 (
            .O(N__66471),
            .I(\quad_counter1.n30574 ));
    InMux I__13438 (
            .O(N__66468),
            .I(N__66463));
    InMux I__13437 (
            .O(N__66467),
            .I(N__66460));
    InMux I__13436 (
            .O(N__66466),
            .I(N__66457));
    LocalMux I__13435 (
            .O(N__66463),
            .I(\quad_counter1.n2907 ));
    LocalMux I__13434 (
            .O(N__66460),
            .I(\quad_counter1.n2907 ));
    LocalMux I__13433 (
            .O(N__66457),
            .I(\quad_counter1.n2907 ));
    InMux I__13432 (
            .O(N__66450),
            .I(\quad_counter1.n30575 ));
    InMux I__13431 (
            .O(N__66447),
            .I(N__66442));
    InMux I__13430 (
            .O(N__66446),
            .I(N__66439));
    InMux I__13429 (
            .O(N__66445),
            .I(N__66436));
    LocalMux I__13428 (
            .O(N__66442),
            .I(\quad_counter1.n2906 ));
    LocalMux I__13427 (
            .O(N__66439),
            .I(\quad_counter1.n2906 ));
    LocalMux I__13426 (
            .O(N__66436),
            .I(\quad_counter1.n2906 ));
    InMux I__13425 (
            .O(N__66429),
            .I(\quad_counter1.n30576 ));
    InMux I__13424 (
            .O(N__66426),
            .I(N__66421));
    InMux I__13423 (
            .O(N__66425),
            .I(N__66418));
    InMux I__13422 (
            .O(N__66424),
            .I(N__66415));
    LocalMux I__13421 (
            .O(N__66421),
            .I(\quad_counter1.n2905 ));
    LocalMux I__13420 (
            .O(N__66418),
            .I(\quad_counter1.n2905 ));
    LocalMux I__13419 (
            .O(N__66415),
            .I(\quad_counter1.n2905 ));
    InMux I__13418 (
            .O(N__66408),
            .I(N__66405));
    LocalMux I__13417 (
            .O(N__66405),
            .I(N__66402));
    Span4Mux_h I__13416 (
            .O(N__66402),
            .I(N__66398));
    InMux I__13415 (
            .O(N__66401),
            .I(N__66395));
    Odrv4 I__13414 (
            .O(N__66398),
            .I(\c0.n33991 ));
    LocalMux I__13413 (
            .O(N__66395),
            .I(\c0.n33991 ));
    InMux I__13412 (
            .O(N__66390),
            .I(N__66387));
    LocalMux I__13411 (
            .O(N__66387),
            .I(N__66383));
    InMux I__13410 (
            .O(N__66386),
            .I(N__66380));
    Odrv12 I__13409 (
            .O(N__66383),
            .I(\c0.n33858 ));
    LocalMux I__13408 (
            .O(N__66380),
            .I(\c0.n33858 ));
    CascadeMux I__13407 (
            .O(N__66375),
            .I(\c0.n10_adj_4673_cascade_ ));
    InMux I__13406 (
            .O(N__66372),
            .I(N__66368));
    InMux I__13405 (
            .O(N__66371),
            .I(N__66364));
    LocalMux I__13404 (
            .O(N__66368),
            .I(N__66361));
    InMux I__13403 (
            .O(N__66367),
            .I(N__66358));
    LocalMux I__13402 (
            .O(N__66364),
            .I(N__66355));
    Span4Mux_v I__13401 (
            .O(N__66361),
            .I(N__66350));
    LocalMux I__13400 (
            .O(N__66358),
            .I(N__66350));
    Odrv4 I__13399 (
            .O(N__66355),
            .I(\c0.n32310 ));
    Odrv4 I__13398 (
            .O(N__66350),
            .I(\c0.n32310 ));
    InMux I__13397 (
            .O(N__66345),
            .I(N__66342));
    LocalMux I__13396 (
            .O(N__66342),
            .I(N__66337));
    InMux I__13395 (
            .O(N__66341),
            .I(N__66334));
    InMux I__13394 (
            .O(N__66340),
            .I(N__66331));
    Span4Mux_h I__13393 (
            .O(N__66337),
            .I(N__66328));
    LocalMux I__13392 (
            .O(N__66334),
            .I(\quad_counter1.n2919 ));
    LocalMux I__13391 (
            .O(N__66331),
            .I(\quad_counter1.n2919 ));
    Odrv4 I__13390 (
            .O(N__66328),
            .I(\quad_counter1.n2919 ));
    InMux I__13389 (
            .O(N__66321),
            .I(bfn_19_2_0_));
    InMux I__13388 (
            .O(N__66318),
            .I(N__66314));
    InMux I__13387 (
            .O(N__66317),
            .I(N__66310));
    LocalMux I__13386 (
            .O(N__66314),
            .I(N__66307));
    CascadeMux I__13385 (
            .O(N__66313),
            .I(N__66304));
    LocalMux I__13384 (
            .O(N__66310),
            .I(N__66299));
    Span4Mux_h I__13383 (
            .O(N__66307),
            .I(N__66299));
    InMux I__13382 (
            .O(N__66304),
            .I(N__66296));
    Odrv4 I__13381 (
            .O(N__66299),
            .I(\quad_counter1.n2918 ));
    LocalMux I__13380 (
            .O(N__66296),
            .I(\quad_counter1.n2918 ));
    InMux I__13379 (
            .O(N__66291),
            .I(\quad_counter1.n30564 ));
    InMux I__13378 (
            .O(N__66288),
            .I(N__66284));
    InMux I__13377 (
            .O(N__66287),
            .I(N__66280));
    LocalMux I__13376 (
            .O(N__66284),
            .I(N__66277));
    InMux I__13375 (
            .O(N__66283),
            .I(N__66274));
    LocalMux I__13374 (
            .O(N__66280),
            .I(\quad_counter1.n2917 ));
    Odrv4 I__13373 (
            .O(N__66277),
            .I(\quad_counter1.n2917 ));
    LocalMux I__13372 (
            .O(N__66274),
            .I(\quad_counter1.n2917 ));
    InMux I__13371 (
            .O(N__66267),
            .I(\quad_counter1.n30565 ));
    InMux I__13370 (
            .O(N__66264),
            .I(N__66259));
    InMux I__13369 (
            .O(N__66263),
            .I(N__66256));
    InMux I__13368 (
            .O(N__66262),
            .I(N__66253));
    LocalMux I__13367 (
            .O(N__66259),
            .I(\quad_counter1.n2916 ));
    LocalMux I__13366 (
            .O(N__66256),
            .I(\quad_counter1.n2916 ));
    LocalMux I__13365 (
            .O(N__66253),
            .I(\quad_counter1.n2916 ));
    InMux I__13364 (
            .O(N__66246),
            .I(\quad_counter1.n30566 ));
    InMux I__13363 (
            .O(N__66243),
            .I(N__66238));
    InMux I__13362 (
            .O(N__66242),
            .I(N__66235));
    InMux I__13361 (
            .O(N__66241),
            .I(N__66232));
    LocalMux I__13360 (
            .O(N__66238),
            .I(\quad_counter1.n2915 ));
    LocalMux I__13359 (
            .O(N__66235),
            .I(\quad_counter1.n2915 ));
    LocalMux I__13358 (
            .O(N__66232),
            .I(\quad_counter1.n2915 ));
    InMux I__13357 (
            .O(N__66225),
            .I(\quad_counter1.n30567 ));
    InMux I__13356 (
            .O(N__66222),
            .I(N__66217));
    InMux I__13355 (
            .O(N__66221),
            .I(N__66214));
    InMux I__13354 (
            .O(N__66220),
            .I(N__66211));
    LocalMux I__13353 (
            .O(N__66217),
            .I(\quad_counter1.n2914 ));
    LocalMux I__13352 (
            .O(N__66214),
            .I(\quad_counter1.n2914 ));
    LocalMux I__13351 (
            .O(N__66211),
            .I(\quad_counter1.n2914 ));
    InMux I__13350 (
            .O(N__66204),
            .I(\quad_counter1.n30568 ));
    InMux I__13349 (
            .O(N__66201),
            .I(N__66198));
    LocalMux I__13348 (
            .O(N__66198),
            .I(\c0.n8_adj_4622 ));
    InMux I__13347 (
            .O(N__66195),
            .I(N__66192));
    LocalMux I__13346 (
            .O(N__66192),
            .I(N__66189));
    Span4Mux_h I__13345 (
            .O(N__66189),
            .I(N__66186));
    Odrv4 I__13344 (
            .O(N__66186),
            .I(\c0.n7_adj_4662 ));
    InMux I__13343 (
            .O(N__66183),
            .I(N__66180));
    LocalMux I__13342 (
            .O(N__66180),
            .I(\c0.n32316 ));
    CascadeMux I__13341 (
            .O(N__66177),
            .I(\c0.n32316_cascade_ ));
    InMux I__13340 (
            .O(N__66174),
            .I(N__66170));
    InMux I__13339 (
            .O(N__66173),
            .I(N__66167));
    LocalMux I__13338 (
            .O(N__66170),
            .I(\c0.n31451 ));
    LocalMux I__13337 (
            .O(N__66167),
            .I(\c0.n31451 ));
    InMux I__13336 (
            .O(N__66162),
            .I(N__66159));
    LocalMux I__13335 (
            .O(N__66159),
            .I(\c0.n21_adj_4659 ));
    CascadeMux I__13334 (
            .O(N__66156),
            .I(\c0.n19_adj_4658_cascade_ ));
    InMux I__13333 (
            .O(N__66153),
            .I(N__66150));
    LocalMux I__13332 (
            .O(N__66150),
            .I(N__66147));
    Span4Mux_v I__13331 (
            .O(N__66147),
            .I(N__66144));
    Odrv4 I__13330 (
            .O(N__66144),
            .I(\c0.n20_adj_4656 ));
    CascadeMux I__13329 (
            .O(N__66141),
            .I(\c0.n5_adj_4660_cascade_ ));
    CascadeMux I__13328 (
            .O(N__66138),
            .I(N__66135));
    InMux I__13327 (
            .O(N__66135),
            .I(N__66130));
    InMux I__13326 (
            .O(N__66134),
            .I(N__66127));
    InMux I__13325 (
            .O(N__66133),
            .I(N__66124));
    LocalMux I__13324 (
            .O(N__66130),
            .I(N__66121));
    LocalMux I__13323 (
            .O(N__66127),
            .I(N__66116));
    LocalMux I__13322 (
            .O(N__66124),
            .I(N__66116));
    Span4Mux_h I__13321 (
            .O(N__66121),
            .I(N__66113));
    Span4Mux_v I__13320 (
            .O(N__66116),
            .I(N__66110));
    Odrv4 I__13319 (
            .O(N__66113),
            .I(\c0.n16118 ));
    Odrv4 I__13318 (
            .O(N__66110),
            .I(\c0.n16118 ));
    InMux I__13317 (
            .O(N__66105),
            .I(N__66101));
    InMux I__13316 (
            .O(N__66104),
            .I(N__66098));
    LocalMux I__13315 (
            .O(N__66101),
            .I(N__66095));
    LocalMux I__13314 (
            .O(N__66098),
            .I(N__66092));
    Span4Mux_h I__13313 (
            .O(N__66095),
            .I(N__66089));
    Odrv4 I__13312 (
            .O(N__66092),
            .I(\c0.n33792 ));
    Odrv4 I__13311 (
            .O(N__66089),
            .I(\c0.n33792 ));
    CascadeMux I__13310 (
            .O(N__66084),
            .I(N__66080));
    InMux I__13309 (
            .O(N__66083),
            .I(N__66076));
    InMux I__13308 (
            .O(N__66080),
            .I(N__66070));
    InMux I__13307 (
            .O(N__66079),
            .I(N__66070));
    LocalMux I__13306 (
            .O(N__66076),
            .I(N__66067));
    InMux I__13305 (
            .O(N__66075),
            .I(N__66064));
    LocalMux I__13304 (
            .O(N__66070),
            .I(\c0.data_in_frame_24_3 ));
    Odrv4 I__13303 (
            .O(N__66067),
            .I(\c0.data_in_frame_24_3 ));
    LocalMux I__13302 (
            .O(N__66064),
            .I(\c0.data_in_frame_24_3 ));
    InMux I__13301 (
            .O(N__66057),
            .I(N__66053));
    InMux I__13300 (
            .O(N__66056),
            .I(N__66050));
    LocalMux I__13299 (
            .O(N__66053),
            .I(N__66047));
    LocalMux I__13298 (
            .O(N__66050),
            .I(\c0.n34006 ));
    Odrv4 I__13297 (
            .O(N__66047),
            .I(\c0.n34006 ));
    InMux I__13296 (
            .O(N__66042),
            .I(N__66036));
    InMux I__13295 (
            .O(N__66041),
            .I(N__66036));
    LocalMux I__13294 (
            .O(N__66036),
            .I(\c0.data_in_frame_28_5 ));
    InMux I__13293 (
            .O(N__66033),
            .I(N__66030));
    LocalMux I__13292 (
            .O(N__66030),
            .I(\c0.n10_adj_4755 ));
    CascadeMux I__13291 (
            .O(N__66027),
            .I(N__66022));
    CascadeMux I__13290 (
            .O(N__66026),
            .I(N__66019));
    CascadeMux I__13289 (
            .O(N__66025),
            .I(N__66014));
    InMux I__13288 (
            .O(N__66022),
            .I(N__66011));
    InMux I__13287 (
            .O(N__66019),
            .I(N__66008));
    InMux I__13286 (
            .O(N__66018),
            .I(N__66005));
    InMux I__13285 (
            .O(N__66017),
            .I(N__66002));
    InMux I__13284 (
            .O(N__66014),
            .I(N__65999));
    LocalMux I__13283 (
            .O(N__66011),
            .I(N__65996));
    LocalMux I__13282 (
            .O(N__66008),
            .I(N__65991));
    LocalMux I__13281 (
            .O(N__66005),
            .I(N__65991));
    LocalMux I__13280 (
            .O(N__66002),
            .I(N__65988));
    LocalMux I__13279 (
            .O(N__65999),
            .I(\c0.data_in_frame_22_0 ));
    Odrv12 I__13278 (
            .O(N__65996),
            .I(\c0.data_in_frame_22_0 ));
    Odrv12 I__13277 (
            .O(N__65991),
            .I(\c0.data_in_frame_22_0 ));
    Odrv4 I__13276 (
            .O(N__65988),
            .I(\c0.data_in_frame_22_0 ));
    InMux I__13275 (
            .O(N__65979),
            .I(N__65976));
    LocalMux I__13274 (
            .O(N__65976),
            .I(\c0.n35142 ));
    InMux I__13273 (
            .O(N__65973),
            .I(N__65970));
    LocalMux I__13272 (
            .O(N__65970),
            .I(N__65967));
    Odrv12 I__13271 (
            .O(N__65967),
            .I(\c0.n35787 ));
    CascadeMux I__13270 (
            .O(N__65964),
            .I(N__65961));
    InMux I__13269 (
            .O(N__65961),
            .I(N__65957));
    InMux I__13268 (
            .O(N__65960),
            .I(N__65954));
    LocalMux I__13267 (
            .O(N__65957),
            .I(N__65949));
    LocalMux I__13266 (
            .O(N__65954),
            .I(N__65949));
    Odrv12 I__13265 (
            .O(N__65949),
            .I(\c0.data_in_frame_26_1 ));
    InMux I__13264 (
            .O(N__65946),
            .I(N__65943));
    LocalMux I__13263 (
            .O(N__65943),
            .I(N__65939));
    InMux I__13262 (
            .O(N__65942),
            .I(N__65934));
    Span4Mux_h I__13261 (
            .O(N__65939),
            .I(N__65931));
    CascadeMux I__13260 (
            .O(N__65938),
            .I(N__65928));
    InMux I__13259 (
            .O(N__65937),
            .I(N__65925));
    LocalMux I__13258 (
            .O(N__65934),
            .I(N__65920));
    Span4Mux_h I__13257 (
            .O(N__65931),
            .I(N__65920));
    InMux I__13256 (
            .O(N__65928),
            .I(N__65917));
    LocalMux I__13255 (
            .O(N__65925),
            .I(\c0.data_in_frame_25_5 ));
    Odrv4 I__13254 (
            .O(N__65920),
            .I(\c0.data_in_frame_25_5 ));
    LocalMux I__13253 (
            .O(N__65917),
            .I(\c0.data_in_frame_25_5 ));
    InMux I__13252 (
            .O(N__65910),
            .I(N__65907));
    LocalMux I__13251 (
            .O(N__65907),
            .I(N__65904));
    Span4Mux_h I__13250 (
            .O(N__65904),
            .I(N__65901));
    Odrv4 I__13249 (
            .O(N__65901),
            .I(\c0.n30_adj_4706 ));
    InMux I__13248 (
            .O(N__65898),
            .I(N__65895));
    LocalMux I__13247 (
            .O(N__65895),
            .I(N__65892));
    Span4Mux_h I__13246 (
            .O(N__65892),
            .I(N__65888));
    InMux I__13245 (
            .O(N__65891),
            .I(N__65885));
    Odrv4 I__13244 (
            .O(N__65888),
            .I(\c0.n33632 ));
    LocalMux I__13243 (
            .O(N__65885),
            .I(\c0.n33632 ));
    InMux I__13242 (
            .O(N__65880),
            .I(N__65876));
    InMux I__13241 (
            .O(N__65879),
            .I(N__65872));
    LocalMux I__13240 (
            .O(N__65876),
            .I(N__65869));
    InMux I__13239 (
            .O(N__65875),
            .I(N__65866));
    LocalMux I__13238 (
            .O(N__65872),
            .I(N__65863));
    Span4Mux_v I__13237 (
            .O(N__65869),
            .I(N__65860));
    LocalMux I__13236 (
            .O(N__65866),
            .I(N__65857));
    Span4Mux_h I__13235 (
            .O(N__65863),
            .I(N__65852));
    Span4Mux_h I__13234 (
            .O(N__65860),
            .I(N__65852));
    Odrv4 I__13233 (
            .O(N__65857),
            .I(\c0.n18405 ));
    Odrv4 I__13232 (
            .O(N__65852),
            .I(\c0.n18405 ));
    CascadeMux I__13231 (
            .O(N__65847),
            .I(N__65843));
    CascadeMux I__13230 (
            .O(N__65846),
            .I(N__65840));
    InMux I__13229 (
            .O(N__65843),
            .I(N__65837));
    InMux I__13228 (
            .O(N__65840),
            .I(N__65833));
    LocalMux I__13227 (
            .O(N__65837),
            .I(N__65830));
    InMux I__13226 (
            .O(N__65836),
            .I(N__65827));
    LocalMux I__13225 (
            .O(N__65833),
            .I(\c0.data_in_frame_25_6 ));
    Odrv12 I__13224 (
            .O(N__65830),
            .I(\c0.data_in_frame_25_6 ));
    LocalMux I__13223 (
            .O(N__65827),
            .I(\c0.data_in_frame_25_6 ));
    CascadeMux I__13222 (
            .O(N__65820),
            .I(N__65817));
    InMux I__13221 (
            .O(N__65817),
            .I(N__65814));
    LocalMux I__13220 (
            .O(N__65814),
            .I(N__65811));
    Odrv4 I__13219 (
            .O(N__65811),
            .I(\c0.n13 ));
    InMux I__13218 (
            .O(N__65808),
            .I(N__65805));
    LocalMux I__13217 (
            .O(N__65805),
            .I(N__65802));
    Span12Mux_h I__13216 (
            .O(N__65802),
            .I(N__65799));
    Odrv12 I__13215 (
            .O(N__65799),
            .I(\c0.n33994 ));
    CascadeMux I__13214 (
            .O(N__65796),
            .I(\c0.n32294_cascade_ ));
    InMux I__13213 (
            .O(N__65793),
            .I(N__65790));
    LocalMux I__13212 (
            .O(N__65790),
            .I(N__65787));
    Span4Mux_v I__13211 (
            .O(N__65787),
            .I(N__65784));
    Odrv4 I__13210 (
            .O(N__65784),
            .I(\c0.n37 ));
    InMux I__13209 (
            .O(N__65781),
            .I(N__65778));
    LocalMux I__13208 (
            .O(N__65778),
            .I(\c0.n18961 ));
    CascadeMux I__13207 (
            .O(N__65775),
            .I(N__65772));
    InMux I__13206 (
            .O(N__65772),
            .I(N__65768));
    CascadeMux I__13205 (
            .O(N__65771),
            .I(N__65765));
    LocalMux I__13204 (
            .O(N__65768),
            .I(N__65762));
    InMux I__13203 (
            .O(N__65765),
            .I(N__65758));
    Span4Mux_h I__13202 (
            .O(N__65762),
            .I(N__65755));
    InMux I__13201 (
            .O(N__65761),
            .I(N__65752));
    LocalMux I__13200 (
            .O(N__65758),
            .I(\c0.data_in_frame_23_1 ));
    Odrv4 I__13199 (
            .O(N__65755),
            .I(\c0.data_in_frame_23_1 ));
    LocalMux I__13198 (
            .O(N__65752),
            .I(\c0.data_in_frame_23_1 ));
    InMux I__13197 (
            .O(N__65745),
            .I(N__65739));
    InMux I__13196 (
            .O(N__65744),
            .I(N__65739));
    LocalMux I__13195 (
            .O(N__65739),
            .I(\c0.n33577 ));
    CascadeMux I__13194 (
            .O(N__65736),
            .I(N__65732));
    InMux I__13193 (
            .O(N__65735),
            .I(N__65728));
    InMux I__13192 (
            .O(N__65732),
            .I(N__65723));
    InMux I__13191 (
            .O(N__65731),
            .I(N__65723));
    LocalMux I__13190 (
            .O(N__65728),
            .I(N__65719));
    LocalMux I__13189 (
            .O(N__65723),
            .I(N__65716));
    InMux I__13188 (
            .O(N__65722),
            .I(N__65713));
    Odrv4 I__13187 (
            .O(N__65719),
            .I(\c0.data_in_frame_23_5 ));
    Odrv4 I__13186 (
            .O(N__65716),
            .I(\c0.data_in_frame_23_5 ));
    LocalMux I__13185 (
            .O(N__65713),
            .I(\c0.data_in_frame_23_5 ));
    InMux I__13184 (
            .O(N__65706),
            .I(N__65703));
    LocalMux I__13183 (
            .O(N__65703),
            .I(N__65700));
    Odrv4 I__13182 (
            .O(N__65700),
            .I(\c0.n35314 ));
    InMux I__13181 (
            .O(N__65697),
            .I(N__65694));
    LocalMux I__13180 (
            .O(N__65694),
            .I(N__65691));
    Span4Mux_h I__13179 (
            .O(N__65691),
            .I(N__65688));
    Odrv4 I__13178 (
            .O(N__65688),
            .I(\c0.n25_adj_4758 ));
    InMux I__13177 (
            .O(N__65685),
            .I(N__65682));
    LocalMux I__13176 (
            .O(N__65682),
            .I(\c0.n31_adj_4763 ));
    InMux I__13175 (
            .O(N__65679),
            .I(N__65674));
    InMux I__13174 (
            .O(N__65678),
            .I(N__65668));
    InMux I__13173 (
            .O(N__65677),
            .I(N__65668));
    LocalMux I__13172 (
            .O(N__65674),
            .I(N__65665));
    CascadeMux I__13171 (
            .O(N__65673),
            .I(N__65662));
    LocalMux I__13170 (
            .O(N__65668),
            .I(N__65659));
    Span4Mux_v I__13169 (
            .O(N__65665),
            .I(N__65656));
    InMux I__13168 (
            .O(N__65662),
            .I(N__65653));
    Span4Mux_h I__13167 (
            .O(N__65659),
            .I(N__65650));
    Span4Mux_h I__13166 (
            .O(N__65656),
            .I(N__65647));
    LocalMux I__13165 (
            .O(N__65653),
            .I(\c0.data_in_frame_22_7 ));
    Odrv4 I__13164 (
            .O(N__65650),
            .I(\c0.data_in_frame_22_7 ));
    Odrv4 I__13163 (
            .O(N__65647),
            .I(\c0.data_in_frame_22_7 ));
    InMux I__13162 (
            .O(N__65640),
            .I(N__65636));
    InMux I__13161 (
            .O(N__65639),
            .I(N__65633));
    LocalMux I__13160 (
            .O(N__65636),
            .I(N__65630));
    LocalMux I__13159 (
            .O(N__65633),
            .I(N__65627));
    Span12Mux_v I__13158 (
            .O(N__65630),
            .I(N__65624));
    Span4Mux_v I__13157 (
            .O(N__65627),
            .I(N__65621));
    Odrv12 I__13156 (
            .O(N__65624),
            .I(\c0.n31374 ));
    Odrv4 I__13155 (
            .O(N__65621),
            .I(\c0.n31374 ));
    InMux I__13154 (
            .O(N__65616),
            .I(N__65613));
    LocalMux I__13153 (
            .O(N__65613),
            .I(N__65610));
    Span4Mux_v I__13152 (
            .O(N__65610),
            .I(N__65607));
    Odrv4 I__13151 (
            .O(N__65607),
            .I(\c0.n33864 ));
    CascadeMux I__13150 (
            .O(N__65604),
            .I(\c0.n18961_cascade_ ));
    InMux I__13149 (
            .O(N__65601),
            .I(N__65598));
    LocalMux I__13148 (
            .O(N__65598),
            .I(N__65595));
    Span4Mux_v I__13147 (
            .O(N__65595),
            .I(N__65592));
    Odrv4 I__13146 (
            .O(N__65592),
            .I(\c0.n14_adj_4668 ));
    InMux I__13145 (
            .O(N__65589),
            .I(N__65585));
    InMux I__13144 (
            .O(N__65588),
            .I(N__65581));
    LocalMux I__13143 (
            .O(N__65585),
            .I(N__65578));
    InMux I__13142 (
            .O(N__65584),
            .I(N__65575));
    LocalMux I__13141 (
            .O(N__65581),
            .I(N__65572));
    Span4Mux_h I__13140 (
            .O(N__65578),
            .I(N__65569));
    LocalMux I__13139 (
            .O(N__65575),
            .I(N__65564));
    Span12Mux_v I__13138 (
            .O(N__65572),
            .I(N__65564));
    Odrv4 I__13137 (
            .O(N__65569),
            .I(\c0.n33665 ));
    Odrv12 I__13136 (
            .O(N__65564),
            .I(\c0.n33665 ));
    CascadeMux I__13135 (
            .O(N__65559),
            .I(N__65556));
    InMux I__13134 (
            .O(N__65556),
            .I(N__65553));
    LocalMux I__13133 (
            .O(N__65553),
            .I(N__65550));
    Span4Mux_h I__13132 (
            .O(N__65550),
            .I(N__65546));
    InMux I__13131 (
            .O(N__65549),
            .I(N__65543));
    Span4Mux_h I__13130 (
            .O(N__65546),
            .I(N__65540));
    LocalMux I__13129 (
            .O(N__65543),
            .I(\c0.n32263 ));
    Odrv4 I__13128 (
            .O(N__65540),
            .I(\c0.n32263 ));
    CascadeMux I__13127 (
            .O(N__65535),
            .I(\c0.n32263_cascade_ ));
    InMux I__13126 (
            .O(N__65532),
            .I(N__65529));
    LocalMux I__13125 (
            .O(N__65529),
            .I(\c0.n33576 ));
    CascadeMux I__13124 (
            .O(N__65526),
            .I(N__65518));
    InMux I__13123 (
            .O(N__65525),
            .I(N__65511));
    InMux I__13122 (
            .O(N__65524),
            .I(N__65511));
    InMux I__13121 (
            .O(N__65523),
            .I(N__65511));
    InMux I__13120 (
            .O(N__65522),
            .I(N__65508));
    CascadeMux I__13119 (
            .O(N__65521),
            .I(N__65505));
    InMux I__13118 (
            .O(N__65518),
            .I(N__65502));
    LocalMux I__13117 (
            .O(N__65511),
            .I(N__65499));
    LocalMux I__13116 (
            .O(N__65508),
            .I(N__65496));
    InMux I__13115 (
            .O(N__65505),
            .I(N__65493));
    LocalMux I__13114 (
            .O(N__65502),
            .I(N__65488));
    Sp12to4 I__13113 (
            .O(N__65499),
            .I(N__65488));
    Span4Mux_h I__13112 (
            .O(N__65496),
            .I(N__65485));
    LocalMux I__13111 (
            .O(N__65493),
            .I(\c0.data_in_frame_19_2 ));
    Odrv12 I__13110 (
            .O(N__65488),
            .I(\c0.data_in_frame_19_2 ));
    Odrv4 I__13109 (
            .O(N__65485),
            .I(\c0.data_in_frame_19_2 ));
    InMux I__13108 (
            .O(N__65478),
            .I(N__65475));
    LocalMux I__13107 (
            .O(N__65475),
            .I(N__65468));
    InMux I__13106 (
            .O(N__65474),
            .I(N__65465));
    InMux I__13105 (
            .O(N__65473),
            .I(N__65458));
    InMux I__13104 (
            .O(N__65472),
            .I(N__65458));
    InMux I__13103 (
            .O(N__65471),
            .I(N__65458));
    Span4Mux_h I__13102 (
            .O(N__65468),
            .I(N__65455));
    LocalMux I__13101 (
            .O(N__65465),
            .I(N__65450));
    LocalMux I__13100 (
            .O(N__65458),
            .I(N__65450));
    Odrv4 I__13099 (
            .O(N__65455),
            .I(\c0.n6215 ));
    Odrv12 I__13098 (
            .O(N__65450),
            .I(\c0.n6215 ));
    CascadeMux I__13097 (
            .O(N__65445),
            .I(\c0.n33576_cascade_ ));
    CascadeMux I__13096 (
            .O(N__65442),
            .I(\c0.n33577_cascade_ ));
    InMux I__13095 (
            .O(N__65439),
            .I(N__65436));
    LocalMux I__13094 (
            .O(N__65436),
            .I(N__65432));
    InMux I__13093 (
            .O(N__65435),
            .I(N__65429));
    Span4Mux_h I__13092 (
            .O(N__65432),
            .I(N__65424));
    LocalMux I__13091 (
            .O(N__65429),
            .I(N__65424));
    Span4Mux_h I__13090 (
            .O(N__65424),
            .I(N__65421));
    Odrv4 I__13089 (
            .O(N__65421),
            .I(\c0.n33638 ));
    InMux I__13088 (
            .O(N__65418),
            .I(N__65415));
    LocalMux I__13087 (
            .O(N__65415),
            .I(\c0.n14_adj_4757 ));
    CascadeMux I__13086 (
            .O(N__65412),
            .I(N__65408));
    InMux I__13085 (
            .O(N__65411),
            .I(N__65405));
    InMux I__13084 (
            .O(N__65408),
            .I(N__65402));
    LocalMux I__13083 (
            .O(N__65405),
            .I(N__65399));
    LocalMux I__13082 (
            .O(N__65402),
            .I(N__65396));
    Span4Mux_h I__13081 (
            .O(N__65399),
            .I(N__65393));
    Span4Mux_v I__13080 (
            .O(N__65396),
            .I(N__65390));
    Span4Mux_v I__13079 (
            .O(N__65393),
            .I(N__65387));
    Span4Mux_v I__13078 (
            .O(N__65390),
            .I(N__65384));
    Odrv4 I__13077 (
            .O(N__65387),
            .I(\c0.n33407 ));
    Odrv4 I__13076 (
            .O(N__65384),
            .I(\c0.n33407 ));
    InMux I__13075 (
            .O(N__65379),
            .I(N__65376));
    LocalMux I__13074 (
            .O(N__65376),
            .I(n2331));
    InMux I__13073 (
            .O(N__65373),
            .I(N__65370));
    LocalMux I__13072 (
            .O(N__65370),
            .I(N__65367));
    Odrv12 I__13071 (
            .O(N__65367),
            .I(\c0.n27862 ));
    InMux I__13070 (
            .O(N__65364),
            .I(N__65360));
    InMux I__13069 (
            .O(N__65363),
            .I(N__65357));
    LocalMux I__13068 (
            .O(N__65360),
            .I(N__65351));
    LocalMux I__13067 (
            .O(N__65357),
            .I(N__65351));
    InMux I__13066 (
            .O(N__65356),
            .I(N__65348));
    Span4Mux_v I__13065 (
            .O(N__65351),
            .I(N__65345));
    LocalMux I__13064 (
            .O(N__65348),
            .I(N__65342));
    Span4Mux_v I__13063 (
            .O(N__65345),
            .I(N__65339));
    Span4Mux_h I__13062 (
            .O(N__65342),
            .I(N__65336));
    Span4Mux_h I__13061 (
            .O(N__65339),
            .I(N__65331));
    Span4Mux_v I__13060 (
            .O(N__65336),
            .I(N__65331));
    Odrv4 I__13059 (
            .O(N__65331),
            .I(\c0.n18084 ));
    InMux I__13058 (
            .O(N__65328),
            .I(N__65325));
    LocalMux I__13057 (
            .O(N__65325),
            .I(N__65321));
    CascadeMux I__13056 (
            .O(N__65324),
            .I(N__65318));
    Span4Mux_h I__13055 (
            .O(N__65321),
            .I(N__65314));
    InMux I__13054 (
            .O(N__65318),
            .I(N__65309));
    InMux I__13053 (
            .O(N__65317),
            .I(N__65309));
    Odrv4 I__13052 (
            .O(N__65314),
            .I(\c0.data_in_frame_25_7 ));
    LocalMux I__13051 (
            .O(N__65309),
            .I(\c0.data_in_frame_25_7 ));
    InMux I__13050 (
            .O(N__65304),
            .I(N__65301));
    LocalMux I__13049 (
            .O(N__65301),
            .I(N__65298));
    Odrv12 I__13048 (
            .O(N__65298),
            .I(\c0.n33_adj_4764 ));
    CascadeMux I__13047 (
            .O(N__65295),
            .I(\c0.n28_adj_4762_cascade_ ));
    InMux I__13046 (
            .O(N__65292),
            .I(N__65289));
    LocalMux I__13045 (
            .O(N__65289),
            .I(N__65286));
    Odrv12 I__13044 (
            .O(N__65286),
            .I(n2249));
    InMux I__13043 (
            .O(N__65283),
            .I(N__65280));
    LocalMux I__13042 (
            .O(N__65280),
            .I(n2339));
    InMux I__13041 (
            .O(N__65277),
            .I(N__65274));
    LocalMux I__13040 (
            .O(N__65274),
            .I(N__65269));
    InMux I__13039 (
            .O(N__65273),
            .I(N__65266));
    InMux I__13038 (
            .O(N__65272),
            .I(N__65263));
    Span4Mux_v I__13037 (
            .O(N__65269),
            .I(N__65259));
    LocalMux I__13036 (
            .O(N__65266),
            .I(N__65254));
    LocalMux I__13035 (
            .O(N__65263),
            .I(N__65254));
    CascadeMux I__13034 (
            .O(N__65262),
            .I(N__65251));
    Span4Mux_h I__13033 (
            .O(N__65259),
            .I(N__65246));
    Span4Mux_v I__13032 (
            .O(N__65254),
            .I(N__65246));
    InMux I__13031 (
            .O(N__65251),
            .I(N__65243));
    Span4Mux_h I__13030 (
            .O(N__65246),
            .I(N__65240));
    LocalMux I__13029 (
            .O(N__65243),
            .I(\c0.data_in_frame_5_3 ));
    Odrv4 I__13028 (
            .O(N__65240),
            .I(\c0.data_in_frame_5_3 ));
    InMux I__13027 (
            .O(N__65235),
            .I(N__65232));
    LocalMux I__13026 (
            .O(N__65232),
            .I(N__65229));
    Odrv12 I__13025 (
            .O(N__65229),
            .I(n2262));
    InMux I__13024 (
            .O(N__65226),
            .I(N__65223));
    LocalMux I__13023 (
            .O(N__65223),
            .I(N__65220));
    Odrv12 I__13022 (
            .O(N__65220),
            .I(n2255));
    InMux I__13021 (
            .O(N__65217),
            .I(N__65213));
    InMux I__13020 (
            .O(N__65216),
            .I(N__65210));
    LocalMux I__13019 (
            .O(N__65213),
            .I(data_out_frame_11_4));
    LocalMux I__13018 (
            .O(N__65210),
            .I(data_out_frame_11_4));
    InMux I__13017 (
            .O(N__65205),
            .I(N__65201));
    InMux I__13016 (
            .O(N__65204),
            .I(N__65198));
    LocalMux I__13015 (
            .O(N__65201),
            .I(data_out_frame_10_4));
    LocalMux I__13014 (
            .O(N__65198),
            .I(data_out_frame_10_4));
    InMux I__13013 (
            .O(N__65193),
            .I(N__65190));
    LocalMux I__13012 (
            .O(N__65190),
            .I(\c0.n35813 ));
    InMux I__13011 (
            .O(N__65187),
            .I(N__65184));
    LocalMux I__13010 (
            .O(N__65184),
            .I(\c0.n35964 ));
    InMux I__13009 (
            .O(N__65181),
            .I(N__65178));
    LocalMux I__13008 (
            .O(N__65178),
            .I(n2325));
    InMux I__13007 (
            .O(N__65175),
            .I(N__65172));
    LocalMux I__13006 (
            .O(N__65172),
            .I(N__65169));
    Span4Mux_h I__13005 (
            .O(N__65169),
            .I(N__65165));
    InMux I__13004 (
            .O(N__65168),
            .I(N__65162));
    Span4Mux_v I__13003 (
            .O(N__65165),
            .I(N__65159));
    LocalMux I__13002 (
            .O(N__65162),
            .I(\c0.data_out_frame_0_4 ));
    Odrv4 I__13001 (
            .O(N__65159),
            .I(\c0.data_out_frame_0_4 ));
    CascadeMux I__13000 (
            .O(N__65154),
            .I(\c0.n36173_cascade_ ));
    CascadeMux I__12999 (
            .O(N__65151),
            .I(\c0.n35814_cascade_ ));
    InMux I__12998 (
            .O(N__65148),
            .I(N__65142));
    InMux I__12997 (
            .O(N__65147),
            .I(N__65139));
    InMux I__12996 (
            .O(N__65146),
            .I(N__65130));
    InMux I__12995 (
            .O(N__65145),
            .I(N__65130));
    LocalMux I__12994 (
            .O(N__65142),
            .I(N__65127));
    LocalMux I__12993 (
            .O(N__65139),
            .I(N__65124));
    InMux I__12992 (
            .O(N__65138),
            .I(N__65116));
    InMux I__12991 (
            .O(N__65137),
            .I(N__65116));
    InMux I__12990 (
            .O(N__65136),
            .I(N__65111));
    InMux I__12989 (
            .O(N__65135),
            .I(N__65111));
    LocalMux I__12988 (
            .O(N__65130),
            .I(N__65104));
    Span4Mux_v I__12987 (
            .O(N__65127),
            .I(N__65104));
    Span4Mux_v I__12986 (
            .O(N__65124),
            .I(N__65104));
    InMux I__12985 (
            .O(N__65123),
            .I(N__65097));
    InMux I__12984 (
            .O(N__65122),
            .I(N__65097));
    InMux I__12983 (
            .O(N__65121),
            .I(N__65097));
    LocalMux I__12982 (
            .O(N__65116),
            .I(r_SM_Main_1));
    LocalMux I__12981 (
            .O(N__65111),
            .I(r_SM_Main_1));
    Odrv4 I__12980 (
            .O(N__65104),
            .I(r_SM_Main_1));
    LocalMux I__12979 (
            .O(N__65097),
            .I(r_SM_Main_1));
    InMux I__12978 (
            .O(N__65088),
            .I(N__65085));
    LocalMux I__12977 (
            .O(N__65085),
            .I(N__65082));
    Span4Mux_h I__12976 (
            .O(N__65082),
            .I(N__65070));
    InMux I__12975 (
            .O(N__65081),
            .I(N__65063));
    InMux I__12974 (
            .O(N__65080),
            .I(N__65063));
    InMux I__12973 (
            .O(N__65079),
            .I(N__65063));
    InMux I__12972 (
            .O(N__65078),
            .I(N__65058));
    InMux I__12971 (
            .O(N__65077),
            .I(N__65058));
    InMux I__12970 (
            .O(N__65076),
            .I(N__65053));
    InMux I__12969 (
            .O(N__65075),
            .I(N__65053));
    InMux I__12968 (
            .O(N__65074),
            .I(N__65048));
    InMux I__12967 (
            .O(N__65073),
            .I(N__65048));
    Odrv4 I__12966 (
            .O(N__65070),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__12965 (
            .O(N__65063),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__12964 (
            .O(N__65058),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__12963 (
            .O(N__65053),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__12962 (
            .O(N__65048),
            .I(\c0.rx.r_SM_Main_0 ));
    InMux I__12961 (
            .O(N__65037),
            .I(N__65033));
    InMux I__12960 (
            .O(N__65036),
            .I(N__65030));
    LocalMux I__12959 (
            .O(N__65033),
            .I(data_out_frame_7_4));
    LocalMux I__12958 (
            .O(N__65030),
            .I(data_out_frame_7_4));
    InMux I__12957 (
            .O(N__65025),
            .I(N__65022));
    LocalMux I__12956 (
            .O(N__65022),
            .I(\c0.n5_adj_4707 ));
    InMux I__12955 (
            .O(N__65019),
            .I(N__65016));
    LocalMux I__12954 (
            .O(N__65016),
            .I(n2345));
    InMux I__12953 (
            .O(N__65013),
            .I(N__65010));
    LocalMux I__12952 (
            .O(N__65010),
            .I(n2342));
    InMux I__12951 (
            .O(N__65007),
            .I(\quad_counter1.n30105 ));
    InMux I__12950 (
            .O(N__65004),
            .I(\quad_counter1.n30106 ));
    CascadeMux I__12949 (
            .O(N__65001),
            .I(N__64990));
    CascadeMux I__12948 (
            .O(N__65000),
            .I(N__64986));
    CascadeMux I__12947 (
            .O(N__64999),
            .I(N__64982));
    CascadeMux I__12946 (
            .O(N__64998),
            .I(N__64978));
    CascadeMux I__12945 (
            .O(N__64997),
            .I(N__64974));
    CascadeMux I__12944 (
            .O(N__64996),
            .I(N__64970));
    CascadeMux I__12943 (
            .O(N__64995),
            .I(N__64966));
    CascadeMux I__12942 (
            .O(N__64994),
            .I(N__64962));
    InMux I__12941 (
            .O(N__64993),
            .I(N__64954));
    InMux I__12940 (
            .O(N__64990),
            .I(N__64937));
    InMux I__12939 (
            .O(N__64989),
            .I(N__64937));
    InMux I__12938 (
            .O(N__64986),
            .I(N__64937));
    InMux I__12937 (
            .O(N__64985),
            .I(N__64937));
    InMux I__12936 (
            .O(N__64982),
            .I(N__64937));
    InMux I__12935 (
            .O(N__64981),
            .I(N__64937));
    InMux I__12934 (
            .O(N__64978),
            .I(N__64937));
    InMux I__12933 (
            .O(N__64977),
            .I(N__64937));
    InMux I__12932 (
            .O(N__64974),
            .I(N__64920));
    InMux I__12931 (
            .O(N__64973),
            .I(N__64920));
    InMux I__12930 (
            .O(N__64970),
            .I(N__64920));
    InMux I__12929 (
            .O(N__64969),
            .I(N__64920));
    InMux I__12928 (
            .O(N__64966),
            .I(N__64920));
    InMux I__12927 (
            .O(N__64965),
            .I(N__64920));
    InMux I__12926 (
            .O(N__64962),
            .I(N__64920));
    InMux I__12925 (
            .O(N__64961),
            .I(N__64920));
    CascadeMux I__12924 (
            .O(N__64960),
            .I(N__64917));
    CascadeMux I__12923 (
            .O(N__64959),
            .I(N__64913));
    CascadeMux I__12922 (
            .O(N__64958),
            .I(N__64909));
    CascadeMux I__12921 (
            .O(N__64957),
            .I(N__64905));
    LocalMux I__12920 (
            .O(N__64954),
            .I(N__64896));
    LocalMux I__12919 (
            .O(N__64937),
            .I(N__64896));
    LocalMux I__12918 (
            .O(N__64920),
            .I(N__64896));
    InMux I__12917 (
            .O(N__64917),
            .I(N__64879));
    InMux I__12916 (
            .O(N__64916),
            .I(N__64879));
    InMux I__12915 (
            .O(N__64913),
            .I(N__64879));
    InMux I__12914 (
            .O(N__64912),
            .I(N__64879));
    InMux I__12913 (
            .O(N__64909),
            .I(N__64879));
    InMux I__12912 (
            .O(N__64908),
            .I(N__64879));
    InMux I__12911 (
            .O(N__64905),
            .I(N__64879));
    InMux I__12910 (
            .O(N__64904),
            .I(N__64879));
    CascadeMux I__12909 (
            .O(N__64903),
            .I(N__64873));
    Span4Mux_v I__12908 (
            .O(N__64896),
            .I(N__64864));
    LocalMux I__12907 (
            .O(N__64879),
            .I(N__64864));
    InMux I__12906 (
            .O(N__64878),
            .I(N__64855));
    InMux I__12905 (
            .O(N__64877),
            .I(N__64855));
    InMux I__12904 (
            .O(N__64876),
            .I(N__64855));
    InMux I__12903 (
            .O(N__64873),
            .I(N__64855));
    InMux I__12902 (
            .O(N__64872),
            .I(N__64846));
    InMux I__12901 (
            .O(N__64871),
            .I(N__64846));
    InMux I__12900 (
            .O(N__64870),
            .I(N__64846));
    InMux I__12899 (
            .O(N__64869),
            .I(N__64846));
    Sp12to4 I__12898 (
            .O(N__64864),
            .I(N__64839));
    LocalMux I__12897 (
            .O(N__64855),
            .I(N__64839));
    LocalMux I__12896 (
            .O(N__64846),
            .I(N__64839));
    Span12Mux_v I__12895 (
            .O(N__64839),
            .I(N__64836));
    Odrv12 I__12894 (
            .O(N__64836),
            .I(\quad_counter1.n2230 ));
    InMux I__12893 (
            .O(N__64833),
            .I(bfn_18_20_0_));
    InMux I__12892 (
            .O(N__64830),
            .I(N__64822));
    InMux I__12891 (
            .O(N__64829),
            .I(N__64819));
    InMux I__12890 (
            .O(N__64828),
            .I(N__64816));
    InMux I__12889 (
            .O(N__64827),
            .I(N__64813));
    InMux I__12888 (
            .O(N__64826),
            .I(N__64810));
    CascadeMux I__12887 (
            .O(N__64825),
            .I(N__64807));
    LocalMux I__12886 (
            .O(N__64822),
            .I(N__64804));
    LocalMux I__12885 (
            .O(N__64819),
            .I(N__64801));
    LocalMux I__12884 (
            .O(N__64816),
            .I(N__64794));
    LocalMux I__12883 (
            .O(N__64813),
            .I(N__64794));
    LocalMux I__12882 (
            .O(N__64810),
            .I(N__64794));
    InMux I__12881 (
            .O(N__64807),
            .I(N__64791));
    Span4Mux_h I__12880 (
            .O(N__64804),
            .I(N__64788));
    Span4Mux_h I__12879 (
            .O(N__64801),
            .I(N__64783));
    Span4Mux_h I__12878 (
            .O(N__64794),
            .I(N__64783));
    LocalMux I__12877 (
            .O(N__64791),
            .I(data_in_frame_1_6));
    Odrv4 I__12876 (
            .O(N__64788),
            .I(data_in_frame_1_6));
    Odrv4 I__12875 (
            .O(N__64783),
            .I(data_in_frame_1_6));
    InMux I__12874 (
            .O(N__64776),
            .I(N__64773));
    LocalMux I__12873 (
            .O(N__64773),
            .I(n2252));
    InMux I__12872 (
            .O(N__64770),
            .I(N__64767));
    LocalMux I__12871 (
            .O(N__64767),
            .I(N__64764));
    Odrv4 I__12870 (
            .O(N__64764),
            .I(n2257));
    InMux I__12869 (
            .O(N__64761),
            .I(N__64758));
    LocalMux I__12868 (
            .O(N__64758),
            .I(N__64755));
    Sp12to4 I__12867 (
            .O(N__64755),
            .I(N__64751));
    InMux I__12866 (
            .O(N__64754),
            .I(N__64748));
    Span12Mux_v I__12865 (
            .O(N__64751),
            .I(N__64745));
    LocalMux I__12864 (
            .O(N__64748),
            .I(data_out_frame_8_7));
    Odrv12 I__12863 (
            .O(N__64745),
            .I(data_out_frame_8_7));
    CascadeMux I__12862 (
            .O(N__64740),
            .I(N__64735));
    CascadeMux I__12861 (
            .O(N__64739),
            .I(N__64732));
    CascadeMux I__12860 (
            .O(N__64738),
            .I(N__64728));
    InMux I__12859 (
            .O(N__64735),
            .I(N__64725));
    InMux I__12858 (
            .O(N__64732),
            .I(N__64722));
    InMux I__12857 (
            .O(N__64731),
            .I(N__64719));
    InMux I__12856 (
            .O(N__64728),
            .I(N__64716));
    LocalMux I__12855 (
            .O(N__64725),
            .I(N__64713));
    LocalMux I__12854 (
            .O(N__64722),
            .I(N__64706));
    LocalMux I__12853 (
            .O(N__64719),
            .I(N__64706));
    LocalMux I__12852 (
            .O(N__64716),
            .I(N__64701));
    Sp12to4 I__12851 (
            .O(N__64713),
            .I(N__64701));
    InMux I__12850 (
            .O(N__64712),
            .I(N__64698));
    InMux I__12849 (
            .O(N__64711),
            .I(N__64695));
    Span4Mux_h I__12848 (
            .O(N__64706),
            .I(N__64692));
    Odrv12 I__12847 (
            .O(N__64701),
            .I(data_in_frame_1_3));
    LocalMux I__12846 (
            .O(N__64698),
            .I(data_in_frame_1_3));
    LocalMux I__12845 (
            .O(N__64695),
            .I(data_in_frame_1_3));
    Odrv4 I__12844 (
            .O(N__64692),
            .I(data_in_frame_1_3));
    InMux I__12843 (
            .O(N__64683),
            .I(N__64680));
    LocalMux I__12842 (
            .O(N__64680),
            .I(n2251));
    InMux I__12841 (
            .O(N__64677),
            .I(\quad_counter1.n30097 ));
    InMux I__12840 (
            .O(N__64674),
            .I(\quad_counter1.n30098 ));
    InMux I__12839 (
            .O(N__64671),
            .I(N__64668));
    LocalMux I__12838 (
            .O(N__64668),
            .I(n2256));
    InMux I__12837 (
            .O(N__64665),
            .I(bfn_18_19_0_));
    InMux I__12836 (
            .O(N__64662),
            .I(\quad_counter1.n30100 ));
    InMux I__12835 (
            .O(N__64659),
            .I(\quad_counter1.n30101 ));
    InMux I__12834 (
            .O(N__64656),
            .I(N__64653));
    LocalMux I__12833 (
            .O(N__64653),
            .I(N__64650));
    Span4Mux_h I__12832 (
            .O(N__64650),
            .I(N__64647));
    Odrv4 I__12831 (
            .O(N__64647),
            .I(n2253));
    InMux I__12830 (
            .O(N__64644),
            .I(\quad_counter1.n30102 ));
    InMux I__12829 (
            .O(N__64641),
            .I(\quad_counter1.n30103 ));
    InMux I__12828 (
            .O(N__64638),
            .I(\quad_counter1.n30104 ));
    InMux I__12827 (
            .O(N__64635),
            .I(\quad_counter1.n30088 ));
    InMux I__12826 (
            .O(N__64632),
            .I(\quad_counter1.n30089 ));
    InMux I__12825 (
            .O(N__64629),
            .I(\quad_counter1.n30090 ));
    InMux I__12824 (
            .O(N__64626),
            .I(bfn_18_18_0_));
    InMux I__12823 (
            .O(N__64623),
            .I(\quad_counter1.n30092 ));
    InMux I__12822 (
            .O(N__64620),
            .I(\quad_counter1.n30093 ));
    InMux I__12821 (
            .O(N__64617),
            .I(\quad_counter1.n30094 ));
    InMux I__12820 (
            .O(N__64614),
            .I(N__64611));
    LocalMux I__12819 (
            .O(N__64611),
            .I(n2260));
    InMux I__12818 (
            .O(N__64608),
            .I(\quad_counter1.n30095 ));
    InMux I__12817 (
            .O(N__64605),
            .I(\quad_counter1.n30096 ));
    InMux I__12816 (
            .O(N__64602),
            .I(\quad_counter1.n30079 ));
    InMux I__12815 (
            .O(N__64599),
            .I(\quad_counter1.n30080 ));
    InMux I__12814 (
            .O(N__64596),
            .I(\quad_counter1.n30081 ));
    InMux I__12813 (
            .O(N__64593),
            .I(\quad_counter1.n30082 ));
    InMux I__12812 (
            .O(N__64590),
            .I(N__64587));
    LocalMux I__12811 (
            .O(N__64587),
            .I(n2272));
    InMux I__12810 (
            .O(N__64584),
            .I(bfn_18_17_0_));
    InMux I__12809 (
            .O(N__64581),
            .I(\quad_counter1.n30084 ));
    InMux I__12808 (
            .O(N__64578),
            .I(\quad_counter1.n30085 ));
    InMux I__12807 (
            .O(N__64575),
            .I(N__64572));
    LocalMux I__12806 (
            .O(N__64572),
            .I(N__64569));
    Odrv4 I__12805 (
            .O(N__64569),
            .I(n2269));
    InMux I__12804 (
            .O(N__64566),
            .I(\quad_counter1.n30086 ));
    InMux I__12803 (
            .O(N__64563),
            .I(\quad_counter1.n30087 ));
    InMux I__12802 (
            .O(N__64560),
            .I(N__64555));
    InMux I__12801 (
            .O(N__64559),
            .I(N__64552));
    InMux I__12800 (
            .O(N__64558),
            .I(N__64549));
    LocalMux I__12799 (
            .O(N__64555),
            .I(\quad_counter0.n2508 ));
    LocalMux I__12798 (
            .O(N__64552),
            .I(\quad_counter0.n2508 ));
    LocalMux I__12797 (
            .O(N__64549),
            .I(\quad_counter0.n2508 ));
    InMux I__12796 (
            .O(N__64542),
            .I(N__64538));
    InMux I__12795 (
            .O(N__64541),
            .I(N__64534));
    LocalMux I__12794 (
            .O(N__64538),
            .I(N__64531));
    InMux I__12793 (
            .O(N__64537),
            .I(N__64528));
    LocalMux I__12792 (
            .O(N__64534),
            .I(\quad_counter0.n2507 ));
    Odrv4 I__12791 (
            .O(N__64531),
            .I(\quad_counter0.n2507 ));
    LocalMux I__12790 (
            .O(N__64528),
            .I(\quad_counter0.n2507 ));
    InMux I__12789 (
            .O(N__64521),
            .I(N__64518));
    LocalMux I__12788 (
            .O(N__64518),
            .I(\quad_counter0.n14 ));
    CascadeMux I__12787 (
            .O(N__64515),
            .I(N__64505));
    CascadeMux I__12786 (
            .O(N__64514),
            .I(N__64502));
    CascadeMux I__12785 (
            .O(N__64513),
            .I(N__64499));
    CascadeMux I__12784 (
            .O(N__64512),
            .I(N__64496));
    CascadeMux I__12783 (
            .O(N__64511),
            .I(N__64493));
    CascadeMux I__12782 (
            .O(N__64510),
            .I(N__64490));
    CascadeMux I__12781 (
            .O(N__64509),
            .I(N__64487));
    CascadeMux I__12780 (
            .O(N__64508),
            .I(N__64484));
    InMux I__12779 (
            .O(N__64505),
            .I(N__64477));
    InMux I__12778 (
            .O(N__64502),
            .I(N__64477));
    InMux I__12777 (
            .O(N__64499),
            .I(N__64477));
    InMux I__12776 (
            .O(N__64496),
            .I(N__64472));
    InMux I__12775 (
            .O(N__64493),
            .I(N__64472));
    InMux I__12774 (
            .O(N__64490),
            .I(N__64465));
    InMux I__12773 (
            .O(N__64487),
            .I(N__64465));
    InMux I__12772 (
            .O(N__64484),
            .I(N__64465));
    LocalMux I__12771 (
            .O(N__64477),
            .I(N__64460));
    LocalMux I__12770 (
            .O(N__64472),
            .I(N__64460));
    LocalMux I__12769 (
            .O(N__64465),
            .I(\quad_counter0.n2540 ));
    Odrv4 I__12768 (
            .O(N__64460),
            .I(\quad_counter0.n2540 ));
    CascadeMux I__12767 (
            .O(N__64455),
            .I(\quad_counter0.n2540_cascade_ ));
    CascadeMux I__12766 (
            .O(N__64452),
            .I(N__64444));
    CascadeMux I__12765 (
            .O(N__64451),
            .I(N__64441));
    CascadeMux I__12764 (
            .O(N__64450),
            .I(N__64438));
    CascadeMux I__12763 (
            .O(N__64449),
            .I(N__64435));
    CascadeMux I__12762 (
            .O(N__64448),
            .I(N__64432));
    CascadeMux I__12761 (
            .O(N__64447),
            .I(N__64429));
    InMux I__12760 (
            .O(N__64444),
            .I(N__64424));
    InMux I__12759 (
            .O(N__64441),
            .I(N__64424));
    InMux I__12758 (
            .O(N__64438),
            .I(N__64415));
    InMux I__12757 (
            .O(N__64435),
            .I(N__64415));
    InMux I__12756 (
            .O(N__64432),
            .I(N__64415));
    InMux I__12755 (
            .O(N__64429),
            .I(N__64415));
    LocalMux I__12754 (
            .O(N__64424),
            .I(N__64410));
    LocalMux I__12753 (
            .O(N__64415),
            .I(N__64410));
    Odrv4 I__12752 (
            .O(N__64410),
            .I(\quad_counter0.n36151 ));
    InMux I__12751 (
            .O(N__64407),
            .I(N__64402));
    InMux I__12750 (
            .O(N__64406),
            .I(N__64399));
    InMux I__12749 (
            .O(N__64405),
            .I(N__64396));
    LocalMux I__12748 (
            .O(N__64402),
            .I(N__64393));
    LocalMux I__12747 (
            .O(N__64399),
            .I(N__64390));
    LocalMux I__12746 (
            .O(N__64396),
            .I(\quad_counter0.n2517 ));
    Odrv4 I__12745 (
            .O(N__64393),
            .I(\quad_counter0.n2517 ));
    Odrv4 I__12744 (
            .O(N__64390),
            .I(\quad_counter0.n2517 ));
    InMux I__12743 (
            .O(N__64383),
            .I(N__64378));
    InMux I__12742 (
            .O(N__64382),
            .I(N__64375));
    InMux I__12741 (
            .O(N__64381),
            .I(N__64372));
    LocalMux I__12740 (
            .O(N__64378),
            .I(N__64369));
    LocalMux I__12739 (
            .O(N__64375),
            .I(\quad_counter0.n2518 ));
    LocalMux I__12738 (
            .O(N__64372),
            .I(\quad_counter0.n2518 ));
    Odrv4 I__12737 (
            .O(N__64369),
            .I(\quad_counter0.n2518 ));
    CascadeMux I__12736 (
            .O(N__64362),
            .I(N__64359));
    InMux I__12735 (
            .O(N__64359),
            .I(N__64356));
    LocalMux I__12734 (
            .O(N__64356),
            .I(\quad_counter0.n28345 ));
    InMux I__12733 (
            .O(N__64353),
            .I(N__64348));
    InMux I__12732 (
            .O(N__64352),
            .I(N__64345));
    InMux I__12731 (
            .O(N__64351),
            .I(N__64342));
    LocalMux I__12730 (
            .O(N__64348),
            .I(N__64339));
    LocalMux I__12729 (
            .O(N__64345),
            .I(\quad_counter0.n2514 ));
    LocalMux I__12728 (
            .O(N__64342),
            .I(\quad_counter0.n2514 ));
    Odrv4 I__12727 (
            .O(N__64339),
            .I(\quad_counter0.n2514 ));
    InMux I__12726 (
            .O(N__64332),
            .I(N__64327));
    InMux I__12725 (
            .O(N__64331),
            .I(N__64324));
    InMux I__12724 (
            .O(N__64330),
            .I(N__64321));
    LocalMux I__12723 (
            .O(N__64327),
            .I(N__64318));
    LocalMux I__12722 (
            .O(N__64324),
            .I(\quad_counter0.n2516 ));
    LocalMux I__12721 (
            .O(N__64321),
            .I(\quad_counter0.n2516 ));
    Odrv4 I__12720 (
            .O(N__64318),
            .I(\quad_counter0.n2516 ));
    InMux I__12719 (
            .O(N__64311),
            .I(N__64306));
    InMux I__12718 (
            .O(N__64310),
            .I(N__64303));
    InMux I__12717 (
            .O(N__64309),
            .I(N__64300));
    LocalMux I__12716 (
            .O(N__64306),
            .I(N__64297));
    LocalMux I__12715 (
            .O(N__64303),
            .I(\quad_counter0.n2515 ));
    LocalMux I__12714 (
            .O(N__64300),
            .I(\quad_counter0.n2515 ));
    Odrv4 I__12713 (
            .O(N__64297),
            .I(\quad_counter0.n2515 ));
    CascadeMux I__12712 (
            .O(N__64290),
            .I(\quad_counter0.n10_adj_4397_cascade_ ));
    InMux I__12711 (
            .O(N__64287),
            .I(N__64282));
    InMux I__12710 (
            .O(N__64286),
            .I(N__64279));
    InMux I__12709 (
            .O(N__64285),
            .I(N__64276));
    LocalMux I__12708 (
            .O(N__64282),
            .I(\quad_counter0.n2510 ));
    LocalMux I__12707 (
            .O(N__64279),
            .I(\quad_counter0.n2510 ));
    LocalMux I__12706 (
            .O(N__64276),
            .I(\quad_counter0.n2510 ));
    CascadeMux I__12705 (
            .O(N__64269),
            .I(N__64266));
    InMux I__12704 (
            .O(N__64266),
            .I(N__64263));
    LocalMux I__12703 (
            .O(N__64263),
            .I(\quad_counter0.n9_adj_4398 ));
    InMux I__12702 (
            .O(N__64260),
            .I(N__64257));
    LocalMux I__12701 (
            .O(N__64257),
            .I(N__64254));
    Span4Mux_v I__12700 (
            .O(N__64254),
            .I(N__64251));
    Span4Mux_v I__12699 (
            .O(N__64251),
            .I(N__64248));
    Span4Mux_v I__12698 (
            .O(N__64248),
            .I(N__64245));
    Odrv4 I__12697 (
            .O(N__64245),
            .I(\quad_counter1.count_direction ));
    InMux I__12696 (
            .O(N__64242),
            .I(N__64239));
    LocalMux I__12695 (
            .O(N__64239),
            .I(n2279));
    InMux I__12694 (
            .O(N__64236),
            .I(\quad_counter1.n30076 ));
    InMux I__12693 (
            .O(N__64233),
            .I(\quad_counter1.n30077 ));
    InMux I__12692 (
            .O(N__64230),
            .I(\quad_counter1.n30078 ));
    CascadeMux I__12691 (
            .O(N__64227),
            .I(N__64219));
    CascadeMux I__12690 (
            .O(N__64226),
            .I(N__64216));
    CascadeMux I__12689 (
            .O(N__64225),
            .I(N__64213));
    CascadeMux I__12688 (
            .O(N__64224),
            .I(N__64210));
    CascadeMux I__12687 (
            .O(N__64223),
            .I(N__64207));
    CascadeMux I__12686 (
            .O(N__64222),
            .I(N__64204));
    InMux I__12685 (
            .O(N__64219),
            .I(N__64199));
    InMux I__12684 (
            .O(N__64216),
            .I(N__64199));
    InMux I__12683 (
            .O(N__64213),
            .I(N__64190));
    InMux I__12682 (
            .O(N__64210),
            .I(N__64190));
    InMux I__12681 (
            .O(N__64207),
            .I(N__64190));
    InMux I__12680 (
            .O(N__64204),
            .I(N__64190));
    LocalMux I__12679 (
            .O(N__64199),
            .I(N__64185));
    LocalMux I__12678 (
            .O(N__64190),
            .I(N__64185));
    Odrv12 I__12677 (
            .O(N__64185),
            .I(\quad_counter0.n36153 ));
    InMux I__12676 (
            .O(N__64182),
            .I(\quad_counter0.n30265 ));
    InMux I__12675 (
            .O(N__64179),
            .I(N__64176));
    LocalMux I__12674 (
            .O(N__64176),
            .I(N__64171));
    InMux I__12673 (
            .O(N__64175),
            .I(N__64168));
    InMux I__12672 (
            .O(N__64174),
            .I(N__64165));
    Span4Mux_h I__12671 (
            .O(N__64171),
            .I(N__64160));
    LocalMux I__12670 (
            .O(N__64168),
            .I(N__64160));
    LocalMux I__12669 (
            .O(N__64165),
            .I(N__64157));
    Span4Mux_h I__12668 (
            .O(N__64160),
            .I(N__64154));
    Odrv4 I__12667 (
            .O(N__64157),
            .I(\quad_counter0.n2413 ));
    Odrv4 I__12666 (
            .O(N__64154),
            .I(\quad_counter0.n2413 ));
    InMux I__12665 (
            .O(N__64149),
            .I(\quad_counter0.n30266 ));
    CascadeMux I__12664 (
            .O(N__64146),
            .I(N__64141));
    InMux I__12663 (
            .O(N__64145),
            .I(N__64138));
    InMux I__12662 (
            .O(N__64144),
            .I(N__64135));
    InMux I__12661 (
            .O(N__64141),
            .I(N__64132));
    LocalMux I__12660 (
            .O(N__64138),
            .I(N__64127));
    LocalMux I__12659 (
            .O(N__64135),
            .I(N__64127));
    LocalMux I__12658 (
            .O(N__64132),
            .I(N__64124));
    Span4Mux_v I__12657 (
            .O(N__64127),
            .I(N__64119));
    Span4Mux_h I__12656 (
            .O(N__64124),
            .I(N__64119));
    Odrv4 I__12655 (
            .O(N__64119),
            .I(\quad_counter0.n2412 ));
    InMux I__12654 (
            .O(N__64116),
            .I(bfn_18_14_0_));
    CascadeMux I__12653 (
            .O(N__64113),
            .I(N__64110));
    InMux I__12652 (
            .O(N__64110),
            .I(N__64105));
    InMux I__12651 (
            .O(N__64109),
            .I(N__64102));
    InMux I__12650 (
            .O(N__64108),
            .I(N__64099));
    LocalMux I__12649 (
            .O(N__64105),
            .I(N__64096));
    LocalMux I__12648 (
            .O(N__64102),
            .I(N__64093));
    LocalMux I__12647 (
            .O(N__64099),
            .I(N__64088));
    Span4Mux_h I__12646 (
            .O(N__64096),
            .I(N__64088));
    Odrv4 I__12645 (
            .O(N__64093),
            .I(\quad_counter0.n2411 ));
    Odrv4 I__12644 (
            .O(N__64088),
            .I(\quad_counter0.n2411 ));
    InMux I__12643 (
            .O(N__64083),
            .I(\quad_counter0.n30268 ));
    InMux I__12642 (
            .O(N__64080),
            .I(N__64075));
    InMux I__12641 (
            .O(N__64079),
            .I(N__64072));
    InMux I__12640 (
            .O(N__64078),
            .I(N__64069));
    LocalMux I__12639 (
            .O(N__64075),
            .I(N__64066));
    LocalMux I__12638 (
            .O(N__64072),
            .I(N__64061));
    LocalMux I__12637 (
            .O(N__64069),
            .I(N__64061));
    Span4Mux_h I__12636 (
            .O(N__64066),
            .I(N__64058));
    Odrv12 I__12635 (
            .O(N__64061),
            .I(\quad_counter0.n2410 ));
    Odrv4 I__12634 (
            .O(N__64058),
            .I(\quad_counter0.n2410 ));
    InMux I__12633 (
            .O(N__64053),
            .I(\quad_counter0.n30269 ));
    InMux I__12632 (
            .O(N__64050),
            .I(N__64045));
    InMux I__12631 (
            .O(N__64049),
            .I(N__64042));
    InMux I__12630 (
            .O(N__64048),
            .I(N__64039));
    LocalMux I__12629 (
            .O(N__64045),
            .I(N__64036));
    LocalMux I__12628 (
            .O(N__64042),
            .I(N__64031));
    LocalMux I__12627 (
            .O(N__64039),
            .I(N__64031));
    Span4Mux_v I__12626 (
            .O(N__64036),
            .I(N__64028));
    Odrv4 I__12625 (
            .O(N__64031),
            .I(\quad_counter0.n2409 ));
    Odrv4 I__12624 (
            .O(N__64028),
            .I(\quad_counter0.n2409 ));
    InMux I__12623 (
            .O(N__64023),
            .I(\quad_counter0.n30270 ));
    InMux I__12622 (
            .O(N__64020),
            .I(N__64015));
    InMux I__12621 (
            .O(N__64019),
            .I(N__64012));
    InMux I__12620 (
            .O(N__64018),
            .I(N__64009));
    LocalMux I__12619 (
            .O(N__64015),
            .I(N__64006));
    LocalMux I__12618 (
            .O(N__64012),
            .I(N__64003));
    LocalMux I__12617 (
            .O(N__64009),
            .I(N__64000));
    Span4Mux_v I__12616 (
            .O(N__64006),
            .I(N__63997));
    Odrv4 I__12615 (
            .O(N__64003),
            .I(\quad_counter0.n2408 ));
    Odrv4 I__12614 (
            .O(N__64000),
            .I(\quad_counter0.n2408 ));
    Odrv4 I__12613 (
            .O(N__63997),
            .I(\quad_counter0.n2408 ));
    CascadeMux I__12612 (
            .O(N__63990),
            .I(N__63983));
    CascadeMux I__12611 (
            .O(N__63989),
            .I(N__63980));
    CascadeMux I__12610 (
            .O(N__63988),
            .I(N__63977));
    CascadeMux I__12609 (
            .O(N__63987),
            .I(N__63974));
    CascadeMux I__12608 (
            .O(N__63986),
            .I(N__63971));
    InMux I__12607 (
            .O(N__63983),
            .I(N__63964));
    InMux I__12606 (
            .O(N__63980),
            .I(N__63964));
    InMux I__12605 (
            .O(N__63977),
            .I(N__63957));
    InMux I__12604 (
            .O(N__63974),
            .I(N__63957));
    InMux I__12603 (
            .O(N__63971),
            .I(N__63957));
    CascadeMux I__12602 (
            .O(N__63970),
            .I(N__63954));
    CascadeMux I__12601 (
            .O(N__63969),
            .I(N__63951));
    LocalMux I__12600 (
            .O(N__63964),
            .I(N__63946));
    LocalMux I__12599 (
            .O(N__63957),
            .I(N__63946));
    InMux I__12598 (
            .O(N__63954),
            .I(N__63941));
    InMux I__12597 (
            .O(N__63951),
            .I(N__63941));
    Span4Mux_h I__12596 (
            .O(N__63946),
            .I(N__63938));
    LocalMux I__12595 (
            .O(N__63941),
            .I(N__63935));
    Odrv4 I__12594 (
            .O(N__63938),
            .I(\quad_counter0.n2441 ));
    Odrv12 I__12593 (
            .O(N__63935),
            .I(\quad_counter0.n2441 ));
    InMux I__12592 (
            .O(N__63930),
            .I(\quad_counter0.n30271 ));
    InMux I__12591 (
            .O(N__63927),
            .I(N__63922));
    InMux I__12590 (
            .O(N__63926),
            .I(N__63918));
    InMux I__12589 (
            .O(N__63925),
            .I(N__63915));
    LocalMux I__12588 (
            .O(N__63922),
            .I(N__63912));
    InMux I__12587 (
            .O(N__63921),
            .I(N__63909));
    LocalMux I__12586 (
            .O(N__63918),
            .I(N__63904));
    LocalMux I__12585 (
            .O(N__63915),
            .I(N__63904));
    Span4Mux_v I__12584 (
            .O(N__63912),
            .I(N__63901));
    LocalMux I__12583 (
            .O(N__63909),
            .I(\quad_counter0.millisecond_counter_18 ));
    Odrv12 I__12582 (
            .O(N__63904),
            .I(\quad_counter0.millisecond_counter_18 ));
    Odrv4 I__12581 (
            .O(N__63901),
            .I(\quad_counter0.millisecond_counter_18 ));
    InMux I__12580 (
            .O(N__63894),
            .I(N__63889));
    InMux I__12579 (
            .O(N__63893),
            .I(N__63886));
    InMux I__12578 (
            .O(N__63892),
            .I(N__63883));
    LocalMux I__12577 (
            .O(N__63889),
            .I(\quad_counter0.n2519 ));
    LocalMux I__12576 (
            .O(N__63886),
            .I(\quad_counter0.n2519 ));
    LocalMux I__12575 (
            .O(N__63883),
            .I(\quad_counter0.n2519 ));
    InMux I__12574 (
            .O(N__63876),
            .I(N__63871));
    InMux I__12573 (
            .O(N__63875),
            .I(N__63868));
    InMux I__12572 (
            .O(N__63874),
            .I(N__63865));
    LocalMux I__12571 (
            .O(N__63871),
            .I(\quad_counter0.n2513 ));
    LocalMux I__12570 (
            .O(N__63868),
            .I(\quad_counter0.n2513 ));
    LocalMux I__12569 (
            .O(N__63865),
            .I(\quad_counter0.n2513 ));
    InMux I__12568 (
            .O(N__63858),
            .I(N__63853));
    InMux I__12567 (
            .O(N__63857),
            .I(N__63850));
    InMux I__12566 (
            .O(N__63856),
            .I(N__63847));
    LocalMux I__12565 (
            .O(N__63853),
            .I(\quad_counter0.n2512 ));
    LocalMux I__12564 (
            .O(N__63850),
            .I(\quad_counter0.n2512 ));
    LocalMux I__12563 (
            .O(N__63847),
            .I(\quad_counter0.n2512 ));
    CascadeMux I__12562 (
            .O(N__63840),
            .I(N__63835));
    InMux I__12561 (
            .O(N__63839),
            .I(N__63832));
    InMux I__12560 (
            .O(N__63838),
            .I(N__63829));
    InMux I__12559 (
            .O(N__63835),
            .I(N__63826));
    LocalMux I__12558 (
            .O(N__63832),
            .I(\quad_counter0.n2511 ));
    LocalMux I__12557 (
            .O(N__63829),
            .I(\quad_counter0.n2511 ));
    LocalMux I__12556 (
            .O(N__63826),
            .I(\quad_counter0.n2511 ));
    InMux I__12555 (
            .O(N__63819),
            .I(N__63814));
    InMux I__12554 (
            .O(N__63818),
            .I(N__63811));
    InMux I__12553 (
            .O(N__63817),
            .I(N__63808));
    LocalMux I__12552 (
            .O(N__63814),
            .I(\quad_counter0.n2509 ));
    LocalMux I__12551 (
            .O(N__63811),
            .I(\quad_counter0.n2509 ));
    LocalMux I__12550 (
            .O(N__63808),
            .I(\quad_counter0.n2509 ));
    InMux I__12549 (
            .O(N__63801),
            .I(N__63797));
    InMux I__12548 (
            .O(N__63800),
            .I(N__63794));
    LocalMux I__12547 (
            .O(N__63797),
            .I(N__63788));
    LocalMux I__12546 (
            .O(N__63794),
            .I(N__63788));
    InMux I__12545 (
            .O(N__63793),
            .I(N__63785));
    Odrv4 I__12544 (
            .O(N__63788),
            .I(\quad_counter0.n2310 ));
    LocalMux I__12543 (
            .O(N__63785),
            .I(\quad_counter0.n2310 ));
    InMux I__12542 (
            .O(N__63780),
            .I(\quad_counter0.n30258 ));
    InMux I__12541 (
            .O(N__63777),
            .I(N__63773));
    InMux I__12540 (
            .O(N__63776),
            .I(N__63770));
    LocalMux I__12539 (
            .O(N__63773),
            .I(N__63764));
    LocalMux I__12538 (
            .O(N__63770),
            .I(N__63764));
    InMux I__12537 (
            .O(N__63769),
            .I(N__63761));
    Odrv12 I__12536 (
            .O(N__63764),
            .I(\quad_counter0.n2309 ));
    LocalMux I__12535 (
            .O(N__63761),
            .I(\quad_counter0.n2309 ));
    CascadeMux I__12534 (
            .O(N__63756),
            .I(N__63750));
    CascadeMux I__12533 (
            .O(N__63755),
            .I(N__63747));
    CascadeMux I__12532 (
            .O(N__63754),
            .I(N__63744));
    CascadeMux I__12531 (
            .O(N__63753),
            .I(N__63741));
    InMux I__12530 (
            .O(N__63750),
            .I(N__63734));
    InMux I__12529 (
            .O(N__63747),
            .I(N__63734));
    InMux I__12528 (
            .O(N__63744),
            .I(N__63729));
    InMux I__12527 (
            .O(N__63741),
            .I(N__63729));
    CascadeMux I__12526 (
            .O(N__63740),
            .I(N__63726));
    CascadeMux I__12525 (
            .O(N__63739),
            .I(N__63723));
    LocalMux I__12524 (
            .O(N__63734),
            .I(N__63718));
    LocalMux I__12523 (
            .O(N__63729),
            .I(N__63718));
    InMux I__12522 (
            .O(N__63726),
            .I(N__63713));
    InMux I__12521 (
            .O(N__63723),
            .I(N__63713));
    Odrv4 I__12520 (
            .O(N__63718),
            .I(\quad_counter0.n2342_adj_4384 ));
    LocalMux I__12519 (
            .O(N__63713),
            .I(\quad_counter0.n2342_adj_4384 ));
    InMux I__12518 (
            .O(N__63708),
            .I(\quad_counter0.n30259 ));
    InMux I__12517 (
            .O(N__63705),
            .I(N__63701));
    InMux I__12516 (
            .O(N__63704),
            .I(N__63698));
    LocalMux I__12515 (
            .O(N__63701),
            .I(N__63692));
    LocalMux I__12514 (
            .O(N__63698),
            .I(N__63692));
    InMux I__12513 (
            .O(N__63697),
            .I(N__63689));
    Span4Mux_h I__12512 (
            .O(N__63692),
            .I(N__63685));
    LocalMux I__12511 (
            .O(N__63689),
            .I(N__63682));
    InMux I__12510 (
            .O(N__63688),
            .I(N__63679));
    Span4Mux_h I__12509 (
            .O(N__63685),
            .I(N__63676));
    Span4Mux_h I__12508 (
            .O(N__63682),
            .I(N__63673));
    LocalMux I__12507 (
            .O(N__63679),
            .I(\quad_counter0.millisecond_counter_19 ));
    Odrv4 I__12506 (
            .O(N__63676),
            .I(\quad_counter0.millisecond_counter_19 ));
    Odrv4 I__12505 (
            .O(N__63673),
            .I(\quad_counter0.millisecond_counter_19 ));
    InMux I__12504 (
            .O(N__63666),
            .I(bfn_18_13_0_));
    CascadeMux I__12503 (
            .O(N__63663),
            .I(N__63659));
    InMux I__12502 (
            .O(N__63662),
            .I(N__63655));
    InMux I__12501 (
            .O(N__63659),
            .I(N__63652));
    InMux I__12500 (
            .O(N__63658),
            .I(N__63649));
    LocalMux I__12499 (
            .O(N__63655),
            .I(N__63646));
    LocalMux I__12498 (
            .O(N__63652),
            .I(N__63643));
    LocalMux I__12497 (
            .O(N__63649),
            .I(N__63640));
    Span4Mux_h I__12496 (
            .O(N__63646),
            .I(N__63637));
    Span4Mux_h I__12495 (
            .O(N__63643),
            .I(N__63634));
    Odrv4 I__12494 (
            .O(N__63640),
            .I(\quad_counter0.n2419 ));
    Odrv4 I__12493 (
            .O(N__63637),
            .I(\quad_counter0.n2419 ));
    Odrv4 I__12492 (
            .O(N__63634),
            .I(\quad_counter0.n2419 ));
    InMux I__12491 (
            .O(N__63627),
            .I(\quad_counter0.n30260 ));
    InMux I__12490 (
            .O(N__63624),
            .I(N__63619));
    InMux I__12489 (
            .O(N__63623),
            .I(N__63616));
    InMux I__12488 (
            .O(N__63622),
            .I(N__63613));
    LocalMux I__12487 (
            .O(N__63619),
            .I(N__63610));
    LocalMux I__12486 (
            .O(N__63616),
            .I(N__63607));
    LocalMux I__12485 (
            .O(N__63613),
            .I(N__63604));
    Odrv12 I__12484 (
            .O(N__63610),
            .I(\quad_counter0.n2418 ));
    Odrv4 I__12483 (
            .O(N__63607),
            .I(\quad_counter0.n2418 ));
    Odrv12 I__12482 (
            .O(N__63604),
            .I(\quad_counter0.n2418 ));
    InMux I__12481 (
            .O(N__63597),
            .I(\quad_counter0.n30261 ));
    InMux I__12480 (
            .O(N__63594),
            .I(\quad_counter0.n30262 ));
    InMux I__12479 (
            .O(N__63591),
            .I(N__63588));
    LocalMux I__12478 (
            .O(N__63588),
            .I(N__63583));
    InMux I__12477 (
            .O(N__63587),
            .I(N__63580));
    InMux I__12476 (
            .O(N__63586),
            .I(N__63577));
    Span4Mux_v I__12475 (
            .O(N__63583),
            .I(N__63574));
    LocalMux I__12474 (
            .O(N__63580),
            .I(N__63569));
    LocalMux I__12473 (
            .O(N__63577),
            .I(N__63569));
    Span4Mux_h I__12472 (
            .O(N__63574),
            .I(N__63566));
    Odrv4 I__12471 (
            .O(N__63569),
            .I(\quad_counter0.n2416 ));
    Odrv4 I__12470 (
            .O(N__63566),
            .I(\quad_counter0.n2416 ));
    InMux I__12469 (
            .O(N__63561),
            .I(\quad_counter0.n30263 ));
    CascadeMux I__12468 (
            .O(N__63558),
            .I(N__63555));
    InMux I__12467 (
            .O(N__63555),
            .I(N__63552));
    LocalMux I__12466 (
            .O(N__63552),
            .I(N__63547));
    InMux I__12465 (
            .O(N__63551),
            .I(N__63544));
    InMux I__12464 (
            .O(N__63550),
            .I(N__63541));
    Span4Mux_h I__12463 (
            .O(N__63547),
            .I(N__63538));
    LocalMux I__12462 (
            .O(N__63544),
            .I(N__63531));
    LocalMux I__12461 (
            .O(N__63541),
            .I(N__63531));
    Span4Mux_h I__12460 (
            .O(N__63538),
            .I(N__63531));
    Odrv4 I__12459 (
            .O(N__63531),
            .I(\quad_counter0.n2415 ));
    InMux I__12458 (
            .O(N__63528),
            .I(\quad_counter0.n30264 ));
    InMux I__12457 (
            .O(N__63525),
            .I(N__63520));
    InMux I__12456 (
            .O(N__63524),
            .I(N__63517));
    InMux I__12455 (
            .O(N__63523),
            .I(N__63514));
    LocalMux I__12454 (
            .O(N__63520),
            .I(N__63511));
    LocalMux I__12453 (
            .O(N__63517),
            .I(N__63508));
    LocalMux I__12452 (
            .O(N__63514),
            .I(N__63505));
    Span4Mux_h I__12451 (
            .O(N__63511),
            .I(N__63502));
    Odrv12 I__12450 (
            .O(N__63508),
            .I(\quad_counter0.n2318_adj_4386 ));
    Odrv4 I__12449 (
            .O(N__63505),
            .I(\quad_counter0.n2318_adj_4386 ));
    Odrv4 I__12448 (
            .O(N__63502),
            .I(\quad_counter0.n2318_adj_4386 ));
    InMux I__12447 (
            .O(N__63495),
            .I(\quad_counter0.n30250 ));
    CascadeMux I__12446 (
            .O(N__63492),
            .I(N__63489));
    InMux I__12445 (
            .O(N__63489),
            .I(N__63484));
    InMux I__12444 (
            .O(N__63488),
            .I(N__63481));
    InMux I__12443 (
            .O(N__63487),
            .I(N__63478));
    LocalMux I__12442 (
            .O(N__63484),
            .I(N__63475));
    LocalMux I__12441 (
            .O(N__63481),
            .I(N__63472));
    LocalMux I__12440 (
            .O(N__63478),
            .I(N__63469));
    Span4Mux_h I__12439 (
            .O(N__63475),
            .I(N__63466));
    Odrv4 I__12438 (
            .O(N__63472),
            .I(\quad_counter0.n2317_adj_4387 ));
    Odrv4 I__12437 (
            .O(N__63469),
            .I(\quad_counter0.n2317_adj_4387 ));
    Odrv4 I__12436 (
            .O(N__63466),
            .I(\quad_counter0.n2317_adj_4387 ));
    InMux I__12435 (
            .O(N__63459),
            .I(\quad_counter0.n30251 ));
    InMux I__12434 (
            .O(N__63456),
            .I(N__63451));
    InMux I__12433 (
            .O(N__63455),
            .I(N__63448));
    InMux I__12432 (
            .O(N__63454),
            .I(N__63445));
    LocalMux I__12431 (
            .O(N__63451),
            .I(N__63442));
    LocalMux I__12430 (
            .O(N__63448),
            .I(N__63437));
    LocalMux I__12429 (
            .O(N__63445),
            .I(N__63437));
    Span4Mux_h I__12428 (
            .O(N__63442),
            .I(N__63434));
    Odrv4 I__12427 (
            .O(N__63437),
            .I(\quad_counter0.n2316_adj_4391 ));
    Odrv4 I__12426 (
            .O(N__63434),
            .I(\quad_counter0.n2316_adj_4391 ));
    InMux I__12425 (
            .O(N__63429),
            .I(\quad_counter0.n30252 ));
    InMux I__12424 (
            .O(N__63426),
            .I(N__63421));
    InMux I__12423 (
            .O(N__63425),
            .I(N__63418));
    InMux I__12422 (
            .O(N__63424),
            .I(N__63415));
    LocalMux I__12421 (
            .O(N__63421),
            .I(N__63412));
    LocalMux I__12420 (
            .O(N__63418),
            .I(N__63409));
    LocalMux I__12419 (
            .O(N__63415),
            .I(N__63406));
    Span4Mux_v I__12418 (
            .O(N__63412),
            .I(N__63403));
    Odrv4 I__12417 (
            .O(N__63409),
            .I(\quad_counter0.n2315_adj_4392 ));
    Odrv12 I__12416 (
            .O(N__63406),
            .I(\quad_counter0.n2315_adj_4392 ));
    Odrv4 I__12415 (
            .O(N__63403),
            .I(\quad_counter0.n2315_adj_4392 ));
    InMux I__12414 (
            .O(N__63396),
            .I(\quad_counter0.n30253 ));
    InMux I__12413 (
            .O(N__63393),
            .I(N__63388));
    InMux I__12412 (
            .O(N__63392),
            .I(N__63385));
    InMux I__12411 (
            .O(N__63391),
            .I(N__63382));
    LocalMux I__12410 (
            .O(N__63388),
            .I(N__63379));
    LocalMux I__12409 (
            .O(N__63385),
            .I(N__63374));
    LocalMux I__12408 (
            .O(N__63382),
            .I(N__63374));
    Span4Mux_v I__12407 (
            .O(N__63379),
            .I(N__63371));
    Odrv4 I__12406 (
            .O(N__63374),
            .I(\quad_counter0.n2314_adj_4388 ));
    Odrv4 I__12405 (
            .O(N__63371),
            .I(\quad_counter0.n2314_adj_4388 ));
    CascadeMux I__12404 (
            .O(N__63366),
            .I(N__63358));
    CascadeMux I__12403 (
            .O(N__63365),
            .I(N__63355));
    CascadeMux I__12402 (
            .O(N__63364),
            .I(N__63352));
    CascadeMux I__12401 (
            .O(N__63363),
            .I(N__63349));
    CascadeMux I__12400 (
            .O(N__63362),
            .I(N__63346));
    CascadeMux I__12399 (
            .O(N__63361),
            .I(N__63343));
    InMux I__12398 (
            .O(N__63358),
            .I(N__63338));
    InMux I__12397 (
            .O(N__63355),
            .I(N__63338));
    InMux I__12396 (
            .O(N__63352),
            .I(N__63329));
    InMux I__12395 (
            .O(N__63349),
            .I(N__63329));
    InMux I__12394 (
            .O(N__63346),
            .I(N__63329));
    InMux I__12393 (
            .O(N__63343),
            .I(N__63329));
    LocalMux I__12392 (
            .O(N__63338),
            .I(\quad_counter0.n36154 ));
    LocalMux I__12391 (
            .O(N__63329),
            .I(\quad_counter0.n36154 ));
    InMux I__12390 (
            .O(N__63324),
            .I(\quad_counter0.n30254 ));
    InMux I__12389 (
            .O(N__63321),
            .I(N__63316));
    InMux I__12388 (
            .O(N__63320),
            .I(N__63313));
    InMux I__12387 (
            .O(N__63319),
            .I(N__63310));
    LocalMux I__12386 (
            .O(N__63316),
            .I(N__63307));
    LocalMux I__12385 (
            .O(N__63313),
            .I(N__63304));
    LocalMux I__12384 (
            .O(N__63310),
            .I(N__63301));
    Span4Mux_h I__12383 (
            .O(N__63307),
            .I(N__63298));
    Odrv12 I__12382 (
            .O(N__63304),
            .I(\quad_counter0.n2313 ));
    Odrv4 I__12381 (
            .O(N__63301),
            .I(\quad_counter0.n2313 ));
    Odrv4 I__12380 (
            .O(N__63298),
            .I(\quad_counter0.n2313 ));
    InMux I__12379 (
            .O(N__63291),
            .I(\quad_counter0.n30255 ));
    InMux I__12378 (
            .O(N__63288),
            .I(N__63283));
    InMux I__12377 (
            .O(N__63287),
            .I(N__63280));
    CascadeMux I__12376 (
            .O(N__63286),
            .I(N__63277));
    LocalMux I__12375 (
            .O(N__63283),
            .I(N__63272));
    LocalMux I__12374 (
            .O(N__63280),
            .I(N__63272));
    InMux I__12373 (
            .O(N__63277),
            .I(N__63269));
    Odrv4 I__12372 (
            .O(N__63272),
            .I(\quad_counter0.n2312 ));
    LocalMux I__12371 (
            .O(N__63269),
            .I(\quad_counter0.n2312 ));
    InMux I__12370 (
            .O(N__63264),
            .I(bfn_18_12_0_));
    InMux I__12369 (
            .O(N__63261),
            .I(N__63256));
    InMux I__12368 (
            .O(N__63260),
            .I(N__63253));
    CascadeMux I__12367 (
            .O(N__63259),
            .I(N__63250));
    LocalMux I__12366 (
            .O(N__63256),
            .I(N__63245));
    LocalMux I__12365 (
            .O(N__63253),
            .I(N__63245));
    InMux I__12364 (
            .O(N__63250),
            .I(N__63242));
    Odrv12 I__12363 (
            .O(N__63245),
            .I(\quad_counter0.n2311 ));
    LocalMux I__12362 (
            .O(N__63242),
            .I(\quad_counter0.n2311 ));
    InMux I__12361 (
            .O(N__63237),
            .I(\quad_counter0.n30257 ));
    InMux I__12360 (
            .O(N__63234),
            .I(N__63229));
    InMux I__12359 (
            .O(N__63233),
            .I(N__63226));
    InMux I__12358 (
            .O(N__63232),
            .I(N__63223));
    LocalMux I__12357 (
            .O(N__63229),
            .I(N__63218));
    LocalMux I__12356 (
            .O(N__63226),
            .I(N__63218));
    LocalMux I__12355 (
            .O(N__63223),
            .I(N__63215));
    Span4Mux_v I__12354 (
            .O(N__63218),
            .I(N__63212));
    Span4Mux_h I__12353 (
            .O(N__63215),
            .I(N__63209));
    Odrv4 I__12352 (
            .O(N__63212),
            .I(\quad_counter0.n2212 ));
    Odrv4 I__12351 (
            .O(N__63209),
            .I(\quad_counter0.n2212 ));
    InMux I__12350 (
            .O(N__63204),
            .I(bfn_18_10_0_));
    InMux I__12349 (
            .O(N__63201),
            .I(N__63196));
    InMux I__12348 (
            .O(N__63200),
            .I(N__63193));
    InMux I__12347 (
            .O(N__63199),
            .I(N__63190));
    LocalMux I__12346 (
            .O(N__63196),
            .I(N__63187));
    LocalMux I__12345 (
            .O(N__63193),
            .I(N__63184));
    LocalMux I__12344 (
            .O(N__63190),
            .I(N__63181));
    Span4Mux_v I__12343 (
            .O(N__63187),
            .I(N__63176));
    Span4Mux_v I__12342 (
            .O(N__63184),
            .I(N__63176));
    Span4Mux_h I__12341 (
            .O(N__63181),
            .I(N__63173));
    Odrv4 I__12340 (
            .O(N__63176),
            .I(\quad_counter0.n2211 ));
    Odrv4 I__12339 (
            .O(N__63173),
            .I(\quad_counter0.n2211 ));
    InMux I__12338 (
            .O(N__63168),
            .I(\quad_counter0.n30247 ));
    InMux I__12337 (
            .O(N__63165),
            .I(N__63161));
    InMux I__12336 (
            .O(N__63164),
            .I(N__63157));
    LocalMux I__12335 (
            .O(N__63161),
            .I(N__63154));
    InMux I__12334 (
            .O(N__63160),
            .I(N__63151));
    LocalMux I__12333 (
            .O(N__63157),
            .I(N__63148));
    Span4Mux_v I__12332 (
            .O(N__63154),
            .I(N__63145));
    LocalMux I__12331 (
            .O(N__63151),
            .I(N__63142));
    Span4Mux_v I__12330 (
            .O(N__63148),
            .I(N__63137));
    Span4Mux_h I__12329 (
            .O(N__63145),
            .I(N__63137));
    Span4Mux_h I__12328 (
            .O(N__63142),
            .I(N__63134));
    Odrv4 I__12327 (
            .O(N__63137),
            .I(\quad_counter0.n2210 ));
    Odrv4 I__12326 (
            .O(N__63134),
            .I(\quad_counter0.n2210 ));
    CascadeMux I__12325 (
            .O(N__63129),
            .I(N__63124));
    CascadeMux I__12324 (
            .O(N__63128),
            .I(N__63121));
    CascadeMux I__12323 (
            .O(N__63127),
            .I(N__63118));
    InMux I__12322 (
            .O(N__63124),
            .I(N__63113));
    InMux I__12321 (
            .O(N__63121),
            .I(N__63108));
    InMux I__12320 (
            .O(N__63118),
            .I(N__63108));
    CascadeMux I__12319 (
            .O(N__63117),
            .I(N__63105));
    CascadeMux I__12318 (
            .O(N__63116),
            .I(N__63102));
    LocalMux I__12317 (
            .O(N__63113),
            .I(N__63097));
    LocalMux I__12316 (
            .O(N__63108),
            .I(N__63097));
    InMux I__12315 (
            .O(N__63105),
            .I(N__63092));
    InMux I__12314 (
            .O(N__63102),
            .I(N__63092));
    Odrv4 I__12313 (
            .O(N__63097),
            .I(\quad_counter0.n2243 ));
    LocalMux I__12312 (
            .O(N__63092),
            .I(\quad_counter0.n2243 ));
    InMux I__12311 (
            .O(N__63087),
            .I(\quad_counter0.n30248 ));
    InMux I__12310 (
            .O(N__63084),
            .I(N__63081));
    LocalMux I__12309 (
            .O(N__63081),
            .I(N__63078));
    Odrv4 I__12308 (
            .O(N__63078),
            .I(\quad_counter0.n7_adj_4393 ));
    CascadeMux I__12307 (
            .O(N__63075),
            .I(\quad_counter0.n2342_adj_4384_cascade_ ));
    InMux I__12306 (
            .O(N__63072),
            .I(N__63069));
    LocalMux I__12305 (
            .O(N__63069),
            .I(N__63066));
    Odrv4 I__12304 (
            .O(N__63066),
            .I(\quad_counter0.n28361 ));
    InMux I__12303 (
            .O(N__63063),
            .I(N__63060));
    LocalMux I__12302 (
            .O(N__63060),
            .I(\quad_counter0.n8_adj_4390 ));
    InMux I__12301 (
            .O(N__63057),
            .I(N__63054));
    LocalMux I__12300 (
            .O(N__63054),
            .I(N__63049));
    InMux I__12299 (
            .O(N__63053),
            .I(N__63045));
    InMux I__12298 (
            .O(N__63052),
            .I(N__63042));
    Span4Mux_v I__12297 (
            .O(N__63049),
            .I(N__63039));
    InMux I__12296 (
            .O(N__63048),
            .I(N__63036));
    LocalMux I__12295 (
            .O(N__63045),
            .I(\quad_counter0.millisecond_counter_20 ));
    LocalMux I__12294 (
            .O(N__63042),
            .I(\quad_counter0.millisecond_counter_20 ));
    Odrv4 I__12293 (
            .O(N__63039),
            .I(\quad_counter0.millisecond_counter_20 ));
    LocalMux I__12292 (
            .O(N__63036),
            .I(\quad_counter0.millisecond_counter_20 ));
    InMux I__12291 (
            .O(N__63027),
            .I(bfn_18_11_0_));
    InMux I__12290 (
            .O(N__63024),
            .I(N__63020));
    InMux I__12289 (
            .O(N__63023),
            .I(N__63017));
    LocalMux I__12288 (
            .O(N__63020),
            .I(N__63011));
    LocalMux I__12287 (
            .O(N__63017),
            .I(N__63011));
    InMux I__12286 (
            .O(N__63016),
            .I(N__63008));
    Odrv4 I__12285 (
            .O(N__63011),
            .I(\quad_counter0.n2319_adj_4385 ));
    LocalMux I__12284 (
            .O(N__63008),
            .I(\quad_counter0.n2319_adj_4385 ));
    InMux I__12283 (
            .O(N__63003),
            .I(\quad_counter0.n30249 ));
    InMux I__12282 (
            .O(N__63000),
            .I(N__62994));
    InMux I__12281 (
            .O(N__62999),
            .I(N__62991));
    InMux I__12280 (
            .O(N__62998),
            .I(N__62988));
    InMux I__12279 (
            .O(N__62997),
            .I(N__62985));
    LocalMux I__12278 (
            .O(N__62994),
            .I(N__62982));
    LocalMux I__12277 (
            .O(N__62991),
            .I(\quad_counter0.millisecond_counter_21 ));
    LocalMux I__12276 (
            .O(N__62988),
            .I(\quad_counter0.millisecond_counter_21 ));
    LocalMux I__12275 (
            .O(N__62985),
            .I(\quad_counter0.millisecond_counter_21 ));
    Odrv4 I__12274 (
            .O(N__62982),
            .I(\quad_counter0.millisecond_counter_21 ));
    InMux I__12273 (
            .O(N__62973),
            .I(bfn_18_9_0_));
    InMux I__12272 (
            .O(N__62970),
            .I(N__62966));
    InMux I__12271 (
            .O(N__62969),
            .I(N__62963));
    LocalMux I__12270 (
            .O(N__62966),
            .I(N__62958));
    LocalMux I__12269 (
            .O(N__62963),
            .I(N__62958));
    Span4Mux_v I__12268 (
            .O(N__62958),
            .I(N__62954));
    InMux I__12267 (
            .O(N__62957),
            .I(N__62951));
    Odrv4 I__12266 (
            .O(N__62954),
            .I(\quad_counter0.n2219 ));
    LocalMux I__12265 (
            .O(N__62951),
            .I(\quad_counter0.n2219 ));
    InMux I__12264 (
            .O(N__62946),
            .I(\quad_counter0.n30239 ));
    InMux I__12263 (
            .O(N__62943),
            .I(N__62940));
    LocalMux I__12262 (
            .O(N__62940),
            .I(N__62935));
    InMux I__12261 (
            .O(N__62939),
            .I(N__62932));
    InMux I__12260 (
            .O(N__62938),
            .I(N__62929));
    Span4Mux_v I__12259 (
            .O(N__62935),
            .I(N__62926));
    LocalMux I__12258 (
            .O(N__62932),
            .I(N__62923));
    LocalMux I__12257 (
            .O(N__62929),
            .I(N__62920));
    Span4Mux_h I__12256 (
            .O(N__62926),
            .I(N__62915));
    Span4Mux_v I__12255 (
            .O(N__62923),
            .I(N__62915));
    Span4Mux_h I__12254 (
            .O(N__62920),
            .I(N__62912));
    Odrv4 I__12253 (
            .O(N__62915),
            .I(\quad_counter0.n2218 ));
    Odrv4 I__12252 (
            .O(N__62912),
            .I(\quad_counter0.n2218 ));
    InMux I__12251 (
            .O(N__62907),
            .I(\quad_counter0.n30240 ));
    CascadeMux I__12250 (
            .O(N__62904),
            .I(N__62899));
    InMux I__12249 (
            .O(N__62903),
            .I(N__62896));
    InMux I__12248 (
            .O(N__62902),
            .I(N__62893));
    InMux I__12247 (
            .O(N__62899),
            .I(N__62890));
    LocalMux I__12246 (
            .O(N__62896),
            .I(N__62887));
    LocalMux I__12245 (
            .O(N__62893),
            .I(N__62882));
    LocalMux I__12244 (
            .O(N__62890),
            .I(N__62882));
    Span4Mux_h I__12243 (
            .O(N__62887),
            .I(N__62879));
    Span4Mux_v I__12242 (
            .O(N__62882),
            .I(N__62876));
    Odrv4 I__12241 (
            .O(N__62879),
            .I(\quad_counter0.n2217 ));
    Odrv4 I__12240 (
            .O(N__62876),
            .I(\quad_counter0.n2217 ));
    InMux I__12239 (
            .O(N__62871),
            .I(\quad_counter0.n30241 ));
    InMux I__12238 (
            .O(N__62868),
            .I(N__62863));
    InMux I__12237 (
            .O(N__62867),
            .I(N__62860));
    InMux I__12236 (
            .O(N__62866),
            .I(N__62857));
    LocalMux I__12235 (
            .O(N__62863),
            .I(N__62854));
    LocalMux I__12234 (
            .O(N__62860),
            .I(N__62849));
    LocalMux I__12233 (
            .O(N__62857),
            .I(N__62849));
    Span4Mux_v I__12232 (
            .O(N__62854),
            .I(N__62844));
    Span4Mux_v I__12231 (
            .O(N__62849),
            .I(N__62844));
    Odrv4 I__12230 (
            .O(N__62844),
            .I(\quad_counter0.n2216 ));
    InMux I__12229 (
            .O(N__62841),
            .I(\quad_counter0.n30242 ));
    InMux I__12228 (
            .O(N__62838),
            .I(N__62833));
    InMux I__12227 (
            .O(N__62837),
            .I(N__62830));
    InMux I__12226 (
            .O(N__62836),
            .I(N__62827));
    LocalMux I__12225 (
            .O(N__62833),
            .I(N__62822));
    LocalMux I__12224 (
            .O(N__62830),
            .I(N__62822));
    LocalMux I__12223 (
            .O(N__62827),
            .I(N__62819));
    Span4Mux_h I__12222 (
            .O(N__62822),
            .I(N__62816));
    Span4Mux_h I__12221 (
            .O(N__62819),
            .I(N__62813));
    Odrv4 I__12220 (
            .O(N__62816),
            .I(\quad_counter0.n2215 ));
    Odrv4 I__12219 (
            .O(N__62813),
            .I(\quad_counter0.n2215 ));
    InMux I__12218 (
            .O(N__62808),
            .I(\quad_counter0.n30243 ));
    InMux I__12217 (
            .O(N__62805),
            .I(N__62800));
    InMux I__12216 (
            .O(N__62804),
            .I(N__62797));
    InMux I__12215 (
            .O(N__62803),
            .I(N__62794));
    LocalMux I__12214 (
            .O(N__62800),
            .I(N__62791));
    LocalMux I__12213 (
            .O(N__62797),
            .I(N__62788));
    LocalMux I__12212 (
            .O(N__62794),
            .I(N__62785));
    Span4Mux_h I__12211 (
            .O(N__62791),
            .I(N__62780));
    Span4Mux_h I__12210 (
            .O(N__62788),
            .I(N__62780));
    Span4Mux_h I__12209 (
            .O(N__62785),
            .I(N__62777));
    Odrv4 I__12208 (
            .O(N__62780),
            .I(\quad_counter0.n2214 ));
    Odrv4 I__12207 (
            .O(N__62777),
            .I(\quad_counter0.n2214 ));
    CascadeMux I__12206 (
            .O(N__62772),
            .I(N__62764));
    CascadeMux I__12205 (
            .O(N__62771),
            .I(N__62761));
    CascadeMux I__12204 (
            .O(N__62770),
            .I(N__62758));
    CascadeMux I__12203 (
            .O(N__62769),
            .I(N__62755));
    CascadeMux I__12202 (
            .O(N__62768),
            .I(N__62752));
    CascadeMux I__12201 (
            .O(N__62767),
            .I(N__62749));
    InMux I__12200 (
            .O(N__62764),
            .I(N__62744));
    InMux I__12199 (
            .O(N__62761),
            .I(N__62744));
    InMux I__12198 (
            .O(N__62758),
            .I(N__62735));
    InMux I__12197 (
            .O(N__62755),
            .I(N__62735));
    InMux I__12196 (
            .O(N__62752),
            .I(N__62735));
    InMux I__12195 (
            .O(N__62749),
            .I(N__62735));
    LocalMux I__12194 (
            .O(N__62744),
            .I(\quad_counter0.n36155 ));
    LocalMux I__12193 (
            .O(N__62735),
            .I(\quad_counter0.n36155 ));
    InMux I__12192 (
            .O(N__62730),
            .I(\quad_counter0.n30244 ));
    InMux I__12191 (
            .O(N__62727),
            .I(N__62722));
    InMux I__12190 (
            .O(N__62726),
            .I(N__62719));
    InMux I__12189 (
            .O(N__62725),
            .I(N__62716));
    LocalMux I__12188 (
            .O(N__62722),
            .I(N__62711));
    LocalMux I__12187 (
            .O(N__62719),
            .I(N__62711));
    LocalMux I__12186 (
            .O(N__62716),
            .I(N__62708));
    Span4Mux_h I__12185 (
            .O(N__62711),
            .I(N__62705));
    Span4Mux_h I__12184 (
            .O(N__62708),
            .I(N__62702));
    Odrv4 I__12183 (
            .O(N__62705),
            .I(\quad_counter0.n2213 ));
    Odrv4 I__12182 (
            .O(N__62702),
            .I(\quad_counter0.n2213 ));
    InMux I__12181 (
            .O(N__62697),
            .I(\quad_counter0.n30245 ));
    InMux I__12180 (
            .O(N__62694),
            .I(N__62691));
    LocalMux I__12179 (
            .O(N__62691),
            .I(N__62688));
    Odrv4 I__12178 (
            .O(N__62688),
            .I(\quad_counter1.n18_adj_4459 ));
    InMux I__12177 (
            .O(N__62685),
            .I(N__62682));
    LocalMux I__12176 (
            .O(N__62682),
            .I(N__62679));
    Odrv4 I__12175 (
            .O(N__62679),
            .I(\quad_counter1.n16_adj_4473 ));
    InMux I__12174 (
            .O(N__62676),
            .I(N__62673));
    LocalMux I__12173 (
            .O(N__62673),
            .I(\quad_counter1.n22_adj_4474 ));
    CascadeMux I__12172 (
            .O(N__62670),
            .I(\quad_counter1.n24_adj_4476_cascade_ ));
    InMux I__12171 (
            .O(N__62667),
            .I(N__62664));
    LocalMux I__12170 (
            .O(N__62664),
            .I(\quad_counter1.n20_adj_4475 ));
    CascadeMux I__12169 (
            .O(N__62661),
            .I(\quad_counter1.n3035_cascade_ ));
    InMux I__12168 (
            .O(N__62658),
            .I(N__62655));
    LocalMux I__12167 (
            .O(N__62655),
            .I(\quad_counter0.n28365 ));
    CascadeMux I__12166 (
            .O(N__62652),
            .I(\quad_counter0.n10_adj_4382_cascade_ ));
    CascadeMux I__12165 (
            .O(N__62649),
            .I(\quad_counter0.n7_adj_4383_cascade_ ));
    CascadeMux I__12164 (
            .O(N__62646),
            .I(\quad_counter0.n2243_cascade_ ));
    InMux I__12163 (
            .O(N__62643),
            .I(\quad_counter1.n30588 ));
    InMux I__12162 (
            .O(N__62640),
            .I(\quad_counter1.n30589 ));
    InMux I__12161 (
            .O(N__62637),
            .I(\quad_counter1.n30590 ));
    InMux I__12160 (
            .O(N__62634),
            .I(\quad_counter1.n30591 ));
    InMux I__12159 (
            .O(N__62631),
            .I(\quad_counter1.n30592 ));
    InMux I__12158 (
            .O(N__62628),
            .I(\quad_counter1.n30593 ));
    InMux I__12157 (
            .O(N__62625),
            .I(\quad_counter1.n30594 ));
    InMux I__12156 (
            .O(N__62622),
            .I(bfn_18_5_0_));
    CascadeMux I__12155 (
            .O(N__62619),
            .I(N__62615));
    CascadeMux I__12154 (
            .O(N__62618),
            .I(N__62612));
    InMux I__12153 (
            .O(N__62615),
            .I(N__62601));
    InMux I__12152 (
            .O(N__62612),
            .I(N__62598));
    CascadeMux I__12151 (
            .O(N__62611),
            .I(N__62595));
    CascadeMux I__12150 (
            .O(N__62610),
            .I(N__62592));
    CascadeMux I__12149 (
            .O(N__62609),
            .I(N__62589));
    CascadeMux I__12148 (
            .O(N__62608),
            .I(N__62586));
    CascadeMux I__12147 (
            .O(N__62607),
            .I(N__62583));
    CascadeMux I__12146 (
            .O(N__62606),
            .I(N__62580));
    CascadeMux I__12145 (
            .O(N__62605),
            .I(N__62577));
    CascadeMux I__12144 (
            .O(N__62604),
            .I(N__62574));
    LocalMux I__12143 (
            .O(N__62601),
            .I(N__62567));
    LocalMux I__12142 (
            .O(N__62598),
            .I(N__62567));
    InMux I__12141 (
            .O(N__62595),
            .I(N__62558));
    InMux I__12140 (
            .O(N__62592),
            .I(N__62558));
    InMux I__12139 (
            .O(N__62589),
            .I(N__62558));
    InMux I__12138 (
            .O(N__62586),
            .I(N__62558));
    InMux I__12137 (
            .O(N__62583),
            .I(N__62549));
    InMux I__12136 (
            .O(N__62580),
            .I(N__62549));
    InMux I__12135 (
            .O(N__62577),
            .I(N__62549));
    InMux I__12134 (
            .O(N__62574),
            .I(N__62549));
    CascadeMux I__12133 (
            .O(N__62573),
            .I(N__62546));
    CascadeMux I__12132 (
            .O(N__62572),
            .I(N__62543));
    Span4Mux_v I__12131 (
            .O(N__62567),
            .I(N__62536));
    LocalMux I__12130 (
            .O(N__62558),
            .I(N__62536));
    LocalMux I__12129 (
            .O(N__62549),
            .I(N__62536));
    InMux I__12128 (
            .O(N__62546),
            .I(N__62531));
    InMux I__12127 (
            .O(N__62543),
            .I(N__62531));
    Odrv4 I__12126 (
            .O(N__62536),
            .I(\quad_counter1.n2936 ));
    LocalMux I__12125 (
            .O(N__62531),
            .I(\quad_counter1.n2936 ));
    InMux I__12124 (
            .O(N__62526),
            .I(\quad_counter1.n30596 ));
    InMux I__12123 (
            .O(N__62523),
            .I(bfn_18_3_0_));
    InMux I__12122 (
            .O(N__62520),
            .I(\quad_counter1.n30580 ));
    InMux I__12121 (
            .O(N__62517),
            .I(\quad_counter1.n30581 ));
    InMux I__12120 (
            .O(N__62514),
            .I(\quad_counter1.n30582 ));
    InMux I__12119 (
            .O(N__62511),
            .I(\quad_counter1.n30583 ));
    InMux I__12118 (
            .O(N__62508),
            .I(\quad_counter1.n30584 ));
    CascadeMux I__12117 (
            .O(N__62505),
            .I(N__62501));
    CascadeMux I__12116 (
            .O(N__62504),
            .I(N__62498));
    InMux I__12115 (
            .O(N__62501),
            .I(N__62489));
    InMux I__12114 (
            .O(N__62498),
            .I(N__62489));
    CascadeMux I__12113 (
            .O(N__62497),
            .I(N__62486));
    CascadeMux I__12112 (
            .O(N__62496),
            .I(N__62483));
    CascadeMux I__12111 (
            .O(N__62495),
            .I(N__62480));
    CascadeMux I__12110 (
            .O(N__62494),
            .I(N__62477));
    LocalMux I__12109 (
            .O(N__62489),
            .I(N__62474));
    InMux I__12108 (
            .O(N__62486),
            .I(N__62465));
    InMux I__12107 (
            .O(N__62483),
            .I(N__62465));
    InMux I__12106 (
            .O(N__62480),
            .I(N__62465));
    InMux I__12105 (
            .O(N__62477),
            .I(N__62465));
    Odrv12 I__12104 (
            .O(N__62474),
            .I(\quad_counter1.n36159 ));
    LocalMux I__12103 (
            .O(N__62465),
            .I(\quad_counter1.n36159 ));
    InMux I__12102 (
            .O(N__62460),
            .I(\quad_counter1.n30585 ));
    InMux I__12101 (
            .O(N__62457),
            .I(\quad_counter1.n30586 ));
    InMux I__12100 (
            .O(N__62454),
            .I(bfn_18_4_0_));
    CascadeMux I__12099 (
            .O(N__62451),
            .I(N__62448));
    InMux I__12098 (
            .O(N__62448),
            .I(N__62444));
    CascadeMux I__12097 (
            .O(N__62447),
            .I(N__62441));
    LocalMux I__12096 (
            .O(N__62444),
            .I(N__62438));
    InMux I__12095 (
            .O(N__62441),
            .I(N__62435));
    Span4Mux_h I__12094 (
            .O(N__62438),
            .I(N__62432));
    LocalMux I__12093 (
            .O(N__62435),
            .I(N__62426));
    Span4Mux_v I__12092 (
            .O(N__62432),
            .I(N__62426));
    InMux I__12091 (
            .O(N__62431),
            .I(N__62423));
    Span4Mux_h I__12090 (
            .O(N__62426),
            .I(N__62420));
    LocalMux I__12089 (
            .O(N__62423),
            .I(\c0.data_in_frame_18_4 ));
    Odrv4 I__12088 (
            .O(N__62420),
            .I(\c0.data_in_frame_18_4 ));
    InMux I__12087 (
            .O(N__62415),
            .I(N__62412));
    LocalMux I__12086 (
            .O(N__62412),
            .I(N__62408));
    InMux I__12085 (
            .O(N__62411),
            .I(N__62404));
    Span4Mux_v I__12084 (
            .O(N__62408),
            .I(N__62401));
    InMux I__12083 (
            .O(N__62407),
            .I(N__62398));
    LocalMux I__12082 (
            .O(N__62404),
            .I(N__62395));
    Odrv4 I__12081 (
            .O(N__62401),
            .I(\c0.n18415 ));
    LocalMux I__12080 (
            .O(N__62398),
            .I(\c0.n18415 ));
    Odrv4 I__12079 (
            .O(N__62395),
            .I(\c0.n18415 ));
    InMux I__12078 (
            .O(N__62388),
            .I(N__62385));
    LocalMux I__12077 (
            .O(N__62385),
            .I(\c0.n29 ));
    CascadeMux I__12076 (
            .O(N__62382),
            .I(\quad_counter1.n2936_cascade_ ));
    InMux I__12075 (
            .O(N__62379),
            .I(N__62376));
    LocalMux I__12074 (
            .O(N__62376),
            .I(\quad_counter1.n28263 ));
    CascadeMux I__12073 (
            .O(N__62373),
            .I(\quad_counter1.n10_adj_4458_cascade_ ));
    InMux I__12072 (
            .O(N__62370),
            .I(N__62367));
    LocalMux I__12071 (
            .O(N__62367),
            .I(\quad_counter1.n20 ));
    CascadeMux I__12070 (
            .O(N__62364),
            .I(\quad_counter1.n13_cascade_ ));
    InMux I__12069 (
            .O(N__62361),
            .I(N__62358));
    LocalMux I__12068 (
            .O(N__62358),
            .I(\quad_counter1.n22 ));
    CascadeMux I__12067 (
            .O(N__62355),
            .I(\c0.n32431_cascade_ ));
    InMux I__12066 (
            .O(N__62352),
            .I(N__62349));
    LocalMux I__12065 (
            .O(N__62349),
            .I(\c0.n32431 ));
    CascadeMux I__12064 (
            .O(N__62346),
            .I(N__62342));
    CascadeMux I__12063 (
            .O(N__62345),
            .I(N__62339));
    InMux I__12062 (
            .O(N__62342),
            .I(N__62336));
    InMux I__12061 (
            .O(N__62339),
            .I(N__62333));
    LocalMux I__12060 (
            .O(N__62336),
            .I(N__62330));
    LocalMux I__12059 (
            .O(N__62333),
            .I(\c0.data_in_frame_29_4 ));
    Odrv12 I__12058 (
            .O(N__62330),
            .I(\c0.data_in_frame_29_4 ));
    InMux I__12057 (
            .O(N__62325),
            .I(N__62321));
    InMux I__12056 (
            .O(N__62324),
            .I(N__62317));
    LocalMux I__12055 (
            .O(N__62321),
            .I(N__62313));
    InMux I__12054 (
            .O(N__62320),
            .I(N__62310));
    LocalMux I__12053 (
            .O(N__62317),
            .I(N__62306));
    InMux I__12052 (
            .O(N__62316),
            .I(N__62303));
    Span4Mux_v I__12051 (
            .O(N__62313),
            .I(N__62300));
    LocalMux I__12050 (
            .O(N__62310),
            .I(N__62297));
    CascadeMux I__12049 (
            .O(N__62309),
            .I(N__62294));
    Span4Mux_v I__12048 (
            .O(N__62306),
            .I(N__62291));
    LocalMux I__12047 (
            .O(N__62303),
            .I(N__62284));
    Span4Mux_v I__12046 (
            .O(N__62300),
            .I(N__62284));
    Span4Mux_v I__12045 (
            .O(N__62297),
            .I(N__62284));
    InMux I__12044 (
            .O(N__62294),
            .I(N__62281));
    Span4Mux_h I__12043 (
            .O(N__62291),
            .I(N__62278));
    Span4Mux_h I__12042 (
            .O(N__62284),
            .I(N__62275));
    LocalMux I__12041 (
            .O(N__62281),
            .I(\c0.data_in_frame_17_3 ));
    Odrv4 I__12040 (
            .O(N__62278),
            .I(\c0.data_in_frame_17_3 ));
    Odrv4 I__12039 (
            .O(N__62275),
            .I(\c0.data_in_frame_17_3 ));
    CascadeMux I__12038 (
            .O(N__62268),
            .I(N__62262));
    CascadeMux I__12037 (
            .O(N__62267),
            .I(N__62255));
    InMux I__12036 (
            .O(N__62266),
            .I(N__62250));
    CascadeMux I__12035 (
            .O(N__62265),
            .I(N__62247));
    InMux I__12034 (
            .O(N__62262),
            .I(N__62242));
    InMux I__12033 (
            .O(N__62261),
            .I(N__62236));
    InMux I__12032 (
            .O(N__62260),
            .I(N__62233));
    CascadeMux I__12031 (
            .O(N__62259),
            .I(N__62230));
    InMux I__12030 (
            .O(N__62258),
            .I(N__62226));
    InMux I__12029 (
            .O(N__62255),
            .I(N__62221));
    CascadeMux I__12028 (
            .O(N__62254),
            .I(N__62218));
    InMux I__12027 (
            .O(N__62253),
            .I(N__62215));
    LocalMux I__12026 (
            .O(N__62250),
            .I(N__62212));
    InMux I__12025 (
            .O(N__62247),
            .I(N__62205));
    InMux I__12024 (
            .O(N__62246),
            .I(N__62205));
    InMux I__12023 (
            .O(N__62245),
            .I(N__62205));
    LocalMux I__12022 (
            .O(N__62242),
            .I(N__62202));
    InMux I__12021 (
            .O(N__62241),
            .I(N__62199));
    CascadeMux I__12020 (
            .O(N__62240),
            .I(N__62196));
    CascadeMux I__12019 (
            .O(N__62239),
            .I(N__62193));
    LocalMux I__12018 (
            .O(N__62236),
            .I(N__62188));
    LocalMux I__12017 (
            .O(N__62233),
            .I(N__62188));
    InMux I__12016 (
            .O(N__62230),
            .I(N__62185));
    InMux I__12015 (
            .O(N__62229),
            .I(N__62182));
    LocalMux I__12014 (
            .O(N__62226),
            .I(N__62179));
    CascadeMux I__12013 (
            .O(N__62225),
            .I(N__62174));
    InMux I__12012 (
            .O(N__62224),
            .I(N__62169));
    LocalMux I__12011 (
            .O(N__62221),
            .I(N__62166));
    InMux I__12010 (
            .O(N__62218),
            .I(N__62163));
    LocalMux I__12009 (
            .O(N__62215),
            .I(N__62160));
    Span4Mux_v I__12008 (
            .O(N__62212),
            .I(N__62155));
    LocalMux I__12007 (
            .O(N__62205),
            .I(N__62155));
    Span4Mux_h I__12006 (
            .O(N__62202),
            .I(N__62150));
    LocalMux I__12005 (
            .O(N__62199),
            .I(N__62150));
    InMux I__12004 (
            .O(N__62196),
            .I(N__62144));
    InMux I__12003 (
            .O(N__62193),
            .I(N__62144));
    Span4Mux_v I__12002 (
            .O(N__62188),
            .I(N__62141));
    LocalMux I__12001 (
            .O(N__62185),
            .I(N__62134));
    LocalMux I__12000 (
            .O(N__62182),
            .I(N__62134));
    Span4Mux_v I__11999 (
            .O(N__62179),
            .I(N__62134));
    CascadeMux I__11998 (
            .O(N__62178),
            .I(N__62131));
    InMux I__11997 (
            .O(N__62177),
            .I(N__62127));
    InMux I__11996 (
            .O(N__62174),
            .I(N__62124));
    InMux I__11995 (
            .O(N__62173),
            .I(N__62119));
    InMux I__11994 (
            .O(N__62172),
            .I(N__62119));
    LocalMux I__11993 (
            .O(N__62169),
            .I(N__62114));
    Span4Mux_h I__11992 (
            .O(N__62166),
            .I(N__62114));
    LocalMux I__11991 (
            .O(N__62163),
            .I(N__62109));
    Span4Mux_h I__11990 (
            .O(N__62160),
            .I(N__62109));
    Span4Mux_h I__11989 (
            .O(N__62155),
            .I(N__62106));
    Span4Mux_h I__11988 (
            .O(N__62150),
            .I(N__62103));
    InMux I__11987 (
            .O(N__62149),
            .I(N__62100));
    LocalMux I__11986 (
            .O(N__62144),
            .I(N__62095));
    Span4Mux_h I__11985 (
            .O(N__62141),
            .I(N__62095));
    Span4Mux_v I__11984 (
            .O(N__62134),
            .I(N__62092));
    InMux I__11983 (
            .O(N__62131),
            .I(N__62087));
    InMux I__11982 (
            .O(N__62130),
            .I(N__62087));
    LocalMux I__11981 (
            .O(N__62127),
            .I(N__62072));
    LocalMux I__11980 (
            .O(N__62124),
            .I(N__62072));
    LocalMux I__11979 (
            .O(N__62119),
            .I(N__62072));
    Span4Mux_v I__11978 (
            .O(N__62114),
            .I(N__62072));
    Span4Mux_h I__11977 (
            .O(N__62109),
            .I(N__62072));
    Span4Mux_h I__11976 (
            .O(N__62106),
            .I(N__62072));
    Span4Mux_v I__11975 (
            .O(N__62103),
            .I(N__62072));
    LocalMux I__11974 (
            .O(N__62100),
            .I(N__62066));
    Span4Mux_v I__11973 (
            .O(N__62095),
            .I(N__62066));
    Span4Mux_v I__11972 (
            .O(N__62092),
            .I(N__62063));
    LocalMux I__11971 (
            .O(N__62087),
            .I(N__62058));
    Span4Mux_v I__11970 (
            .O(N__62072),
            .I(N__62058));
    InMux I__11969 (
            .O(N__62071),
            .I(N__62055));
    Span4Mux_v I__11968 (
            .O(N__62066),
            .I(N__62050));
    Span4Mux_v I__11967 (
            .O(N__62063),
            .I(N__62050));
    Span4Mux_v I__11966 (
            .O(N__62058),
            .I(N__62045));
    LocalMux I__11965 (
            .O(N__62055),
            .I(N__62045));
    Odrv4 I__11964 (
            .O(N__62050),
            .I(\c0.n18011 ));
    Odrv4 I__11963 (
            .O(N__62045),
            .I(\c0.n18011 ));
    CascadeMux I__11962 (
            .O(N__62040),
            .I(N__62036));
    InMux I__11961 (
            .O(N__62039),
            .I(N__62033));
    InMux I__11960 (
            .O(N__62036),
            .I(N__62030));
    LocalMux I__11959 (
            .O(N__62033),
            .I(N__62027));
    LocalMux I__11958 (
            .O(N__62030),
            .I(N__62022));
    Span4Mux_h I__11957 (
            .O(N__62027),
            .I(N__62019));
    InMux I__11956 (
            .O(N__62026),
            .I(N__62014));
    InMux I__11955 (
            .O(N__62025),
            .I(N__62014));
    Odrv4 I__11954 (
            .O(N__62022),
            .I(\c0.data_in_frame_23_4 ));
    Odrv4 I__11953 (
            .O(N__62019),
            .I(\c0.data_in_frame_23_4 ));
    LocalMux I__11952 (
            .O(N__62014),
            .I(\c0.data_in_frame_23_4 ));
    InMux I__11951 (
            .O(N__62007),
            .I(N__62004));
    LocalMux I__11950 (
            .O(N__62004),
            .I(N__62000));
    CascadeMux I__11949 (
            .O(N__62003),
            .I(N__61996));
    Span4Mux_h I__11948 (
            .O(N__62000),
            .I(N__61993));
    InMux I__11947 (
            .O(N__61999),
            .I(N__61989));
    InMux I__11946 (
            .O(N__61996),
            .I(N__61986));
    Span4Mux_v I__11945 (
            .O(N__61993),
            .I(N__61983));
    InMux I__11944 (
            .O(N__61992),
            .I(N__61980));
    LocalMux I__11943 (
            .O(N__61989),
            .I(N__61977));
    LocalMux I__11942 (
            .O(N__61986),
            .I(N__61972));
    Span4Mux_h I__11941 (
            .O(N__61983),
            .I(N__61972));
    LocalMux I__11940 (
            .O(N__61980),
            .I(\c0.data_in_frame_16_4 ));
    Odrv12 I__11939 (
            .O(N__61977),
            .I(\c0.data_in_frame_16_4 ));
    Odrv4 I__11938 (
            .O(N__61972),
            .I(\c0.data_in_frame_16_4 ));
    InMux I__11937 (
            .O(N__61965),
            .I(\quad_counter0.n30138 ));
    CascadeMux I__11936 (
            .O(N__61962),
            .I(N__61951));
    CascadeMux I__11935 (
            .O(N__61961),
            .I(N__61947));
    CascadeMux I__11934 (
            .O(N__61960),
            .I(N__61943));
    CascadeMux I__11933 (
            .O(N__61959),
            .I(N__61939));
    CascadeMux I__11932 (
            .O(N__61958),
            .I(N__61934));
    CascadeMux I__11931 (
            .O(N__61957),
            .I(N__61930));
    CascadeMux I__11930 (
            .O(N__61956),
            .I(N__61926));
    CascadeMux I__11929 (
            .O(N__61955),
            .I(N__61922));
    InMux I__11928 (
            .O(N__61954),
            .I(N__61911));
    InMux I__11927 (
            .O(N__61951),
            .I(N__61894));
    InMux I__11926 (
            .O(N__61950),
            .I(N__61894));
    InMux I__11925 (
            .O(N__61947),
            .I(N__61894));
    InMux I__11924 (
            .O(N__61946),
            .I(N__61894));
    InMux I__11923 (
            .O(N__61943),
            .I(N__61894));
    InMux I__11922 (
            .O(N__61942),
            .I(N__61894));
    InMux I__11921 (
            .O(N__61939),
            .I(N__61894));
    InMux I__11920 (
            .O(N__61938),
            .I(N__61894));
    InMux I__11919 (
            .O(N__61937),
            .I(N__61877));
    InMux I__11918 (
            .O(N__61934),
            .I(N__61877));
    InMux I__11917 (
            .O(N__61933),
            .I(N__61877));
    InMux I__11916 (
            .O(N__61930),
            .I(N__61877));
    InMux I__11915 (
            .O(N__61929),
            .I(N__61877));
    InMux I__11914 (
            .O(N__61926),
            .I(N__61877));
    InMux I__11913 (
            .O(N__61925),
            .I(N__61877));
    InMux I__11912 (
            .O(N__61922),
            .I(N__61877));
    CascadeMux I__11911 (
            .O(N__61921),
            .I(N__61874));
    CascadeMux I__11910 (
            .O(N__61920),
            .I(N__61870));
    CascadeMux I__11909 (
            .O(N__61919),
            .I(N__61866));
    CascadeMux I__11908 (
            .O(N__61918),
            .I(N__61862));
    CascadeMux I__11907 (
            .O(N__61917),
            .I(N__61858));
    CascadeMux I__11906 (
            .O(N__61916),
            .I(N__61855));
    CascadeMux I__11905 (
            .O(N__61915),
            .I(N__61851));
    CascadeMux I__11904 (
            .O(N__61914),
            .I(N__61847));
    LocalMux I__11903 (
            .O(N__61911),
            .I(N__61838));
    LocalMux I__11902 (
            .O(N__61894),
            .I(N__61838));
    LocalMux I__11901 (
            .O(N__61877),
            .I(N__61838));
    InMux I__11900 (
            .O(N__61874),
            .I(N__61821));
    InMux I__11899 (
            .O(N__61873),
            .I(N__61821));
    InMux I__11898 (
            .O(N__61870),
            .I(N__61821));
    InMux I__11897 (
            .O(N__61869),
            .I(N__61821));
    InMux I__11896 (
            .O(N__61866),
            .I(N__61821));
    InMux I__11895 (
            .O(N__61865),
            .I(N__61821));
    InMux I__11894 (
            .O(N__61862),
            .I(N__61821));
    InMux I__11893 (
            .O(N__61861),
            .I(N__61821));
    InMux I__11892 (
            .O(N__61858),
            .I(N__61818));
    InMux I__11891 (
            .O(N__61855),
            .I(N__61803));
    InMux I__11890 (
            .O(N__61854),
            .I(N__61803));
    InMux I__11889 (
            .O(N__61851),
            .I(N__61803));
    InMux I__11888 (
            .O(N__61850),
            .I(N__61803));
    InMux I__11887 (
            .O(N__61847),
            .I(N__61803));
    InMux I__11886 (
            .O(N__61846),
            .I(N__61803));
    InMux I__11885 (
            .O(N__61845),
            .I(N__61803));
    Span4Mux_v I__11884 (
            .O(N__61838),
            .I(N__61798));
    LocalMux I__11883 (
            .O(N__61821),
            .I(N__61798));
    LocalMux I__11882 (
            .O(N__61818),
            .I(N__61793));
    LocalMux I__11881 (
            .O(N__61803),
            .I(N__61793));
    Span4Mux_h I__11880 (
            .O(N__61798),
            .I(N__61790));
    Span4Mux_h I__11879 (
            .O(N__61793),
            .I(N__61787));
    Span4Mux_h I__11878 (
            .O(N__61790),
            .I(N__61784));
    Span4Mux_h I__11877 (
            .O(N__61787),
            .I(N__61781));
    Odrv4 I__11876 (
            .O(N__61784),
            .I(\quad_counter0.n2300 ));
    Odrv4 I__11875 (
            .O(N__61781),
            .I(\quad_counter0.n2300 ));
    InMux I__11874 (
            .O(N__61776),
            .I(bfn_17_26_0_));
    InMux I__11873 (
            .O(N__61773),
            .I(N__61770));
    LocalMux I__11872 (
            .O(N__61770),
            .I(\c0.n12_adj_4759 ));
    InMux I__11871 (
            .O(N__61767),
            .I(N__61764));
    LocalMux I__11870 (
            .O(N__61764),
            .I(N__61761));
    Span4Mux_h I__11869 (
            .O(N__61761),
            .I(N__61758));
    Odrv4 I__11868 (
            .O(N__61758),
            .I(\c0.n34841 ));
    CascadeMux I__11867 (
            .O(N__61755),
            .I(N__61752));
    InMux I__11866 (
            .O(N__61752),
            .I(N__61749));
    LocalMux I__11865 (
            .O(N__61749),
            .I(N__61746));
    Span4Mux_h I__11864 (
            .O(N__61746),
            .I(N__61743));
    Odrv4 I__11863 (
            .O(N__61743),
            .I(\c0.n6_adj_4666 ));
    InMux I__11862 (
            .O(N__61740),
            .I(N__61736));
    InMux I__11861 (
            .O(N__61739),
            .I(N__61733));
    LocalMux I__11860 (
            .O(N__61736),
            .I(N__61730));
    LocalMux I__11859 (
            .O(N__61733),
            .I(N__61727));
    Odrv4 I__11858 (
            .O(N__61730),
            .I(\c0.n32366 ));
    Odrv4 I__11857 (
            .O(N__61727),
            .I(\c0.n32366 ));
    InMux I__11856 (
            .O(N__61722),
            .I(N__61716));
    InMux I__11855 (
            .O(N__61721),
            .I(N__61711));
    InMux I__11854 (
            .O(N__61720),
            .I(N__61711));
    InMux I__11853 (
            .O(N__61719),
            .I(N__61708));
    LocalMux I__11852 (
            .O(N__61716),
            .I(\c0.data_in_frame_21_7 ));
    LocalMux I__11851 (
            .O(N__61711),
            .I(\c0.data_in_frame_21_7 ));
    LocalMux I__11850 (
            .O(N__61708),
            .I(\c0.data_in_frame_21_7 ));
    CascadeMux I__11849 (
            .O(N__61701),
            .I(N__61695));
    InMux I__11848 (
            .O(N__61700),
            .I(N__61690));
    InMux I__11847 (
            .O(N__61699),
            .I(N__61690));
    InMux I__11846 (
            .O(N__61698),
            .I(N__61687));
    InMux I__11845 (
            .O(N__61695),
            .I(N__61684));
    LocalMux I__11844 (
            .O(N__61690),
            .I(N__61679));
    LocalMux I__11843 (
            .O(N__61687),
            .I(N__61679));
    LocalMux I__11842 (
            .O(N__61684),
            .I(N__61674));
    Span4Mux_v I__11841 (
            .O(N__61679),
            .I(N__61674));
    Odrv4 I__11840 (
            .O(N__61674),
            .I(\c0.data_in_frame_21_6 ));
    InMux I__11839 (
            .O(N__61671),
            .I(N__61667));
    CascadeMux I__11838 (
            .O(N__61670),
            .I(N__61664));
    LocalMux I__11837 (
            .O(N__61667),
            .I(N__61660));
    InMux I__11836 (
            .O(N__61664),
            .I(N__61656));
    InMux I__11835 (
            .O(N__61663),
            .I(N__61653));
    Span4Mux_v I__11834 (
            .O(N__61660),
            .I(N__61650));
    InMux I__11833 (
            .O(N__61659),
            .I(N__61647));
    LocalMux I__11832 (
            .O(N__61656),
            .I(\c0.data_in_frame_24_1 ));
    LocalMux I__11831 (
            .O(N__61653),
            .I(\c0.data_in_frame_24_1 ));
    Odrv4 I__11830 (
            .O(N__61650),
            .I(\c0.data_in_frame_24_1 ));
    LocalMux I__11829 (
            .O(N__61647),
            .I(\c0.data_in_frame_24_1 ));
    InMux I__11828 (
            .O(N__61638),
            .I(N__61635));
    LocalMux I__11827 (
            .O(N__61635),
            .I(N__61632));
    Span4Mux_h I__11826 (
            .O(N__61632),
            .I(N__61628));
    InMux I__11825 (
            .O(N__61631),
            .I(N__61625));
    Odrv4 I__11824 (
            .O(N__61628),
            .I(\c0.n33662 ));
    LocalMux I__11823 (
            .O(N__61625),
            .I(\c0.n33662 ));
    CascadeMux I__11822 (
            .O(N__61620),
            .I(\c0.n36530_cascade_ ));
    InMux I__11821 (
            .O(N__61617),
            .I(N__61612));
    InMux I__11820 (
            .O(N__61616),
            .I(N__61609));
    InMux I__11819 (
            .O(N__61615),
            .I(N__61605));
    LocalMux I__11818 (
            .O(N__61612),
            .I(N__61600));
    LocalMux I__11817 (
            .O(N__61609),
            .I(N__61600));
    InMux I__11816 (
            .O(N__61608),
            .I(N__61597));
    LocalMux I__11815 (
            .O(N__61605),
            .I(N__61592));
    Span4Mux_h I__11814 (
            .O(N__61600),
            .I(N__61592));
    LocalMux I__11813 (
            .O(N__61597),
            .I(encoder0_position_21));
    Odrv4 I__11812 (
            .O(N__61592),
            .I(encoder0_position_21));
    InMux I__11811 (
            .O(N__61587),
            .I(N__61584));
    LocalMux I__11810 (
            .O(N__61584),
            .I(n2324));
    InMux I__11809 (
            .O(N__61581),
            .I(\quad_counter0.n30129 ));
    InMux I__11808 (
            .O(N__61578),
            .I(N__61575));
    LocalMux I__11807 (
            .O(N__61575),
            .I(N__61572));
    Span4Mux_h I__11806 (
            .O(N__61572),
            .I(N__61569));
    Odrv4 I__11805 (
            .O(N__61569),
            .I(n2323));
    InMux I__11804 (
            .O(N__61566),
            .I(\quad_counter0.n30130 ));
    InMux I__11803 (
            .O(N__61563),
            .I(bfn_17_25_0_));
    InMux I__11802 (
            .O(N__61560),
            .I(\quad_counter0.n30132 ));
    InMux I__11801 (
            .O(N__61557),
            .I(\quad_counter0.n30133 ));
    InMux I__11800 (
            .O(N__61554),
            .I(\quad_counter0.n30134 ));
    InMux I__11799 (
            .O(N__61551),
            .I(N__61548));
    LocalMux I__11798 (
            .O(N__61548),
            .I(n2318));
    InMux I__11797 (
            .O(N__61545),
            .I(\quad_counter0.n30135 ));
    InMux I__11796 (
            .O(N__61542),
            .I(\quad_counter0.n30136 ));
    InMux I__11795 (
            .O(N__61539),
            .I(N__61536));
    LocalMux I__11794 (
            .O(N__61536),
            .I(N__61533));
    Span4Mux_h I__11793 (
            .O(N__61533),
            .I(N__61530));
    Odrv4 I__11792 (
            .O(N__61530),
            .I(n2316));
    InMux I__11791 (
            .O(N__61527),
            .I(\quad_counter0.n30137 ));
    InMux I__11790 (
            .O(N__61524),
            .I(\quad_counter0.n30120 ));
    InMux I__11789 (
            .O(N__61521),
            .I(\quad_counter0.n30121 ));
    InMux I__11788 (
            .O(N__61518),
            .I(\quad_counter0.n30122 ));
    InMux I__11787 (
            .O(N__61515),
            .I(bfn_17_24_0_));
    InMux I__11786 (
            .O(N__61512),
            .I(\quad_counter0.n30124 ));
    InMux I__11785 (
            .O(N__61509),
            .I(\quad_counter0.n30125 ));
    InMux I__11784 (
            .O(N__61506),
            .I(\quad_counter0.n30126 ));
    InMux I__11783 (
            .O(N__61503),
            .I(N__61500));
    LocalMux I__11782 (
            .O(N__61500),
            .I(N__61497));
    Span4Mux_h I__11781 (
            .O(N__61497),
            .I(N__61494));
    Odrv4 I__11780 (
            .O(N__61494),
            .I(n2326));
    InMux I__11779 (
            .O(N__61491),
            .I(\quad_counter0.n30127 ));
    InMux I__11778 (
            .O(N__61488),
            .I(\quad_counter0.n30128 ));
    InMux I__11777 (
            .O(N__61485),
            .I(\quad_counter0.n30111 ));
    InMux I__11776 (
            .O(N__61482),
            .I(\quad_counter0.n30112 ));
    InMux I__11775 (
            .O(N__61479),
            .I(\quad_counter0.n30113 ));
    InMux I__11774 (
            .O(N__61476),
            .I(\quad_counter0.n30114 ));
    InMux I__11773 (
            .O(N__61473),
            .I(bfn_17_23_0_));
    InMux I__11772 (
            .O(N__61470),
            .I(\quad_counter0.n30116 ));
    InMux I__11771 (
            .O(N__61467),
            .I(\quad_counter0.n30117 ));
    InMux I__11770 (
            .O(N__61464),
            .I(\quad_counter0.n30118 ));
    InMux I__11769 (
            .O(N__61461),
            .I(\quad_counter0.n30119 ));
    CascadeMux I__11768 (
            .O(N__61458),
            .I(N__61454));
    InMux I__11767 (
            .O(N__61457),
            .I(N__61449));
    InMux I__11766 (
            .O(N__61454),
            .I(N__61444));
    InMux I__11765 (
            .O(N__61453),
            .I(N__61444));
    InMux I__11764 (
            .O(N__61452),
            .I(N__61441));
    LocalMux I__11763 (
            .O(N__61449),
            .I(N__61430));
    LocalMux I__11762 (
            .O(N__61444),
            .I(N__61430));
    LocalMux I__11761 (
            .O(N__61441),
            .I(N__61430));
    InMux I__11760 (
            .O(N__61440),
            .I(N__61425));
    InMux I__11759 (
            .O(N__61439),
            .I(N__61425));
    InMux I__11758 (
            .O(N__61438),
            .I(N__61422));
    CascadeMux I__11757 (
            .O(N__61437),
            .I(N__61419));
    Span4Mux_h I__11756 (
            .O(N__61430),
            .I(N__61416));
    LocalMux I__11755 (
            .O(N__61425),
            .I(N__61411));
    LocalMux I__11754 (
            .O(N__61422),
            .I(N__61411));
    InMux I__11753 (
            .O(N__61419),
            .I(N__61408));
    Span4Mux_h I__11752 (
            .O(N__61416),
            .I(N__61405));
    Span12Mux_h I__11751 (
            .O(N__61411),
            .I(N__61402));
    LocalMux I__11750 (
            .O(N__61408),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__11749 (
            .O(N__61405),
            .I(\c0.data_in_frame_0_7 ));
    Odrv12 I__11748 (
            .O(N__61402),
            .I(\c0.data_in_frame_0_7 ));
    InMux I__11747 (
            .O(N__61395),
            .I(N__61392));
    LocalMux I__11746 (
            .O(N__61392),
            .I(N__61388));
    InMux I__11745 (
            .O(N__61391),
            .I(N__61385));
    Span4Mux_v I__11744 (
            .O(N__61388),
            .I(N__61382));
    LocalMux I__11743 (
            .O(N__61385),
            .I(data_out_frame_8_6));
    Odrv4 I__11742 (
            .O(N__61382),
            .I(data_out_frame_8_6));
    InMux I__11741 (
            .O(N__61377),
            .I(N__61373));
    InMux I__11740 (
            .O(N__61376),
            .I(N__61370));
    LocalMux I__11739 (
            .O(N__61373),
            .I(N__61367));
    LocalMux I__11738 (
            .O(N__61370),
            .I(data_out_frame_5_6));
    Odrv4 I__11737 (
            .O(N__61367),
            .I(data_out_frame_5_6));
    InMux I__11736 (
            .O(N__61362),
            .I(N__61359));
    LocalMux I__11735 (
            .O(N__61359),
            .I(N__61356));
    Sp12to4 I__11734 (
            .O(N__61356),
            .I(N__61353));
    Odrv12 I__11733 (
            .O(N__61353),
            .I(\quad_counter0.count_direction ));
    InMux I__11732 (
            .O(N__61350),
            .I(\quad_counter0.n30108 ));
    InMux I__11731 (
            .O(N__61347),
            .I(\quad_counter0.n30109 ));
    InMux I__11730 (
            .O(N__61344),
            .I(\quad_counter0.n30110 ));
    InMux I__11729 (
            .O(N__61341),
            .I(N__61337));
    CascadeMux I__11728 (
            .O(N__61340),
            .I(N__61334));
    LocalMux I__11727 (
            .O(N__61337),
            .I(N__61331));
    InMux I__11726 (
            .O(N__61334),
            .I(N__61328));
    Span4Mux_h I__11725 (
            .O(N__61331),
            .I(N__61325));
    LocalMux I__11724 (
            .O(N__61328),
            .I(\c0.data_in_frame_6_4 ));
    Odrv4 I__11723 (
            .O(N__61325),
            .I(\c0.data_in_frame_6_4 ));
    InMux I__11722 (
            .O(N__61320),
            .I(N__61314));
    InMux I__11721 (
            .O(N__61319),
            .I(N__61314));
    LocalMux I__11720 (
            .O(N__61314),
            .I(N__61311));
    Odrv4 I__11719 (
            .O(N__61311),
            .I(data_out_frame_6_5));
    CascadeMux I__11718 (
            .O(N__61308),
            .I(N__61305));
    InMux I__11717 (
            .O(N__61305),
            .I(N__61299));
    InMux I__11716 (
            .O(N__61304),
            .I(N__61299));
    LocalMux I__11715 (
            .O(N__61299),
            .I(data_out_frame_7_5));
    InMux I__11714 (
            .O(N__61296),
            .I(N__61293));
    LocalMux I__11713 (
            .O(N__61293),
            .I(\c0.n36086 ));
    CascadeMux I__11712 (
            .O(N__61290),
            .I(\c0.n5_adj_4619_cascade_ ));
    InMux I__11711 (
            .O(N__61287),
            .I(N__61283));
    InMux I__11710 (
            .O(N__61286),
            .I(N__61280));
    LocalMux I__11709 (
            .O(N__61283),
            .I(N__61277));
    LocalMux I__11708 (
            .O(N__61280),
            .I(data_out_frame_6_6));
    Odrv4 I__11707 (
            .O(N__61277),
            .I(data_out_frame_6_6));
    InMux I__11706 (
            .O(N__61272),
            .I(N__61269));
    LocalMux I__11705 (
            .O(N__61269),
            .I(N__61266));
    Odrv4 I__11704 (
            .O(N__61266),
            .I(\c0.n36012 ));
    InMux I__11703 (
            .O(N__61263),
            .I(N__61260));
    LocalMux I__11702 (
            .O(N__61260),
            .I(N__61257));
    Span4Mux_v I__11701 (
            .O(N__61257),
            .I(N__61254));
    Odrv4 I__11700 (
            .O(N__61254),
            .I(\c0.n5_adj_4624 ));
    InMux I__11699 (
            .O(N__61251),
            .I(N__61248));
    LocalMux I__11698 (
            .O(N__61248),
            .I(N__61244));
    InMux I__11697 (
            .O(N__61247),
            .I(N__61241));
    Span4Mux_h I__11696 (
            .O(N__61244),
            .I(N__61238));
    LocalMux I__11695 (
            .O(N__61241),
            .I(data_out_frame_9_1));
    Odrv4 I__11694 (
            .O(N__61238),
            .I(data_out_frame_9_1));
    InMux I__11693 (
            .O(N__61233),
            .I(N__61230));
    LocalMux I__11692 (
            .O(N__61230),
            .I(N__61227));
    Span4Mux_h I__11691 (
            .O(N__61227),
            .I(N__61223));
    InMux I__11690 (
            .O(N__61226),
            .I(N__61220));
    Odrv4 I__11689 (
            .O(N__61223),
            .I(\c0.n33500 ));
    LocalMux I__11688 (
            .O(N__61220),
            .I(\c0.n33500 ));
    InMux I__11687 (
            .O(N__61215),
            .I(N__61211));
    InMux I__11686 (
            .O(N__61214),
            .I(N__61206));
    LocalMux I__11685 (
            .O(N__61211),
            .I(N__61203));
    InMux I__11684 (
            .O(N__61210),
            .I(N__61200));
    InMux I__11683 (
            .O(N__61209),
            .I(N__61197));
    LocalMux I__11682 (
            .O(N__61206),
            .I(N__61190));
    Sp12to4 I__11681 (
            .O(N__61203),
            .I(N__61190));
    LocalMux I__11680 (
            .O(N__61200),
            .I(N__61190));
    LocalMux I__11679 (
            .O(N__61197),
            .I(\c0.n18627 ));
    Odrv12 I__11678 (
            .O(N__61190),
            .I(\c0.n18627 ));
    InMux I__11677 (
            .O(N__61185),
            .I(N__61181));
    InMux I__11676 (
            .O(N__61184),
            .I(N__61178));
    LocalMux I__11675 (
            .O(N__61181),
            .I(N__61173));
    LocalMux I__11674 (
            .O(N__61178),
            .I(N__61170));
    InMux I__11673 (
            .O(N__61177),
            .I(N__61167));
    InMux I__11672 (
            .O(N__61176),
            .I(N__61164));
    Span4Mux_h I__11671 (
            .O(N__61173),
            .I(N__61161));
    Span4Mux_v I__11670 (
            .O(N__61170),
            .I(N__61158));
    LocalMux I__11669 (
            .O(N__61167),
            .I(N__61155));
    LocalMux I__11668 (
            .O(N__61164),
            .I(N__61152));
    Span4Mux_h I__11667 (
            .O(N__61161),
            .I(N__61149));
    Span4Mux_h I__11666 (
            .O(N__61158),
            .I(N__61146));
    Span4Mux_h I__11665 (
            .O(N__61155),
            .I(N__61143));
    Span4Mux_h I__11664 (
            .O(N__61152),
            .I(N__61140));
    Span4Mux_v I__11663 (
            .O(N__61149),
            .I(N__61137));
    Span4Mux_h I__11662 (
            .O(N__61146),
            .I(N__61134));
    Span4Mux_h I__11661 (
            .O(N__61143),
            .I(N__61129));
    Span4Mux_h I__11660 (
            .O(N__61140),
            .I(N__61129));
    Odrv4 I__11659 (
            .O(N__61137),
            .I(\c0.n18479 ));
    Odrv4 I__11658 (
            .O(N__61134),
            .I(\c0.n18479 ));
    Odrv4 I__11657 (
            .O(N__61129),
            .I(\c0.n18479 ));
    InMux I__11656 (
            .O(N__61122),
            .I(N__61119));
    LocalMux I__11655 (
            .O(N__61119),
            .I(N__61115));
    InMux I__11654 (
            .O(N__61118),
            .I(N__61112));
    Odrv4 I__11653 (
            .O(N__61115),
            .I(data_out_frame_11_7));
    LocalMux I__11652 (
            .O(N__61112),
            .I(data_out_frame_11_7));
    InMux I__11651 (
            .O(N__61107),
            .I(N__61103));
    InMux I__11650 (
            .O(N__61106),
            .I(N__61100));
    LocalMux I__11649 (
            .O(N__61103),
            .I(data_out_frame_5_5));
    LocalMux I__11648 (
            .O(N__61100),
            .I(data_out_frame_5_5));
    InMux I__11647 (
            .O(N__61095),
            .I(N__61092));
    LocalMux I__11646 (
            .O(N__61092),
            .I(N__61088));
    InMux I__11645 (
            .O(N__61091),
            .I(N__61085));
    Span4Mux_h I__11644 (
            .O(N__61088),
            .I(N__61082));
    LocalMux I__11643 (
            .O(N__61085),
            .I(data_out_frame_7_2));
    Odrv4 I__11642 (
            .O(N__61082),
            .I(data_out_frame_7_2));
    InMux I__11641 (
            .O(N__61077),
            .I(N__61074));
    LocalMux I__11640 (
            .O(N__61074),
            .I(\c0.n36021 ));
    InMux I__11639 (
            .O(N__61071),
            .I(N__61067));
    InMux I__11638 (
            .O(N__61070),
            .I(N__61064));
    LocalMux I__11637 (
            .O(N__61067),
            .I(data_out_frame_11_0));
    LocalMux I__11636 (
            .O(N__61064),
            .I(data_out_frame_11_0));
    InMux I__11635 (
            .O(N__61059),
            .I(N__61055));
    InMux I__11634 (
            .O(N__61058),
            .I(N__61052));
    LocalMux I__11633 (
            .O(N__61055),
            .I(data_out_frame_10_0));
    LocalMux I__11632 (
            .O(N__61052),
            .I(data_out_frame_10_0));
    InMux I__11631 (
            .O(N__61047),
            .I(N__61044));
    LocalMux I__11630 (
            .O(N__61044),
            .I(N__61041));
    Span4Mux_h I__11629 (
            .O(N__61041),
            .I(N__61038));
    Odrv4 I__11628 (
            .O(N__61038),
            .I(\c0.n36197 ));
    InMux I__11627 (
            .O(N__61035),
            .I(N__61031));
    InMux I__11626 (
            .O(N__61034),
            .I(N__61028));
    LocalMux I__11625 (
            .O(N__61031),
            .I(data_out_frame_13_7));
    LocalMux I__11624 (
            .O(N__61028),
            .I(data_out_frame_13_7));
    InMux I__11623 (
            .O(N__61023),
            .I(N__61020));
    LocalMux I__11622 (
            .O(N__61020),
            .I(\c0.n36191 ));
    InMux I__11621 (
            .O(N__61017),
            .I(N__61013));
    InMux I__11620 (
            .O(N__61016),
            .I(N__61010));
    LocalMux I__11619 (
            .O(N__61013),
            .I(data_out_frame_10_6));
    LocalMux I__11618 (
            .O(N__61010),
            .I(data_out_frame_10_6));
    InMux I__11617 (
            .O(N__61005),
            .I(N__60999));
    InMux I__11616 (
            .O(N__61004),
            .I(N__60999));
    LocalMux I__11615 (
            .O(N__60999),
            .I(data_out_frame_11_6));
    CascadeMux I__11614 (
            .O(N__60996),
            .I(N__60993));
    InMux I__11613 (
            .O(N__60993),
            .I(N__60987));
    InMux I__11612 (
            .O(N__60992),
            .I(N__60987));
    LocalMux I__11611 (
            .O(N__60987),
            .I(data_out_frame_9_6));
    CascadeMux I__11610 (
            .O(N__60984),
            .I(\c0.n36185_cascade_ ));
    InMux I__11609 (
            .O(N__60981),
            .I(N__60978));
    LocalMux I__11608 (
            .O(N__60978),
            .I(N__60975));
    Span4Mux_v I__11607 (
            .O(N__60975),
            .I(N__60972));
    Odrv4 I__11606 (
            .O(N__60972),
            .I(\c0.n36188 ));
    InMux I__11605 (
            .O(N__60969),
            .I(N__60966));
    LocalMux I__11604 (
            .O(N__60966),
            .I(\c0.n5_adj_4515 ));
    InMux I__11603 (
            .O(N__60963),
            .I(N__60960));
    LocalMux I__11602 (
            .O(N__60960),
            .I(\c0.n6_adj_4514 ));
    CascadeMux I__11601 (
            .O(N__60957),
            .I(\c0.n35836_cascade_ ));
    InMux I__11600 (
            .O(N__60954),
            .I(N__60951));
    LocalMux I__11599 (
            .O(N__60951),
            .I(n35838));
    InMux I__11598 (
            .O(N__60948),
            .I(N__60944));
    InMux I__11597 (
            .O(N__60947),
            .I(N__60941));
    LocalMux I__11596 (
            .O(N__60944),
            .I(data_out_frame_10_3));
    LocalMux I__11595 (
            .O(N__60941),
            .I(data_out_frame_10_3));
    InMux I__11594 (
            .O(N__60936),
            .I(N__60932));
    InMux I__11593 (
            .O(N__60935),
            .I(N__60929));
    LocalMux I__11592 (
            .O(N__60932),
            .I(data_out_frame_8_3));
    LocalMux I__11591 (
            .O(N__60929),
            .I(data_out_frame_8_3));
    InMux I__11590 (
            .O(N__60924),
            .I(N__60920));
    InMux I__11589 (
            .O(N__60923),
            .I(N__60917));
    LocalMux I__11588 (
            .O(N__60920),
            .I(data_out_frame_12_7));
    LocalMux I__11587 (
            .O(N__60917),
            .I(data_out_frame_12_7));
    InMux I__11586 (
            .O(N__60912),
            .I(N__60908));
    InMux I__11585 (
            .O(N__60911),
            .I(N__60905));
    LocalMux I__11584 (
            .O(N__60908),
            .I(N__60899));
    LocalMux I__11583 (
            .O(N__60905),
            .I(N__60899));
    InMux I__11582 (
            .O(N__60904),
            .I(N__60896));
    Span4Mux_h I__11581 (
            .O(N__60899),
            .I(N__60893));
    LocalMux I__11580 (
            .O(N__60896),
            .I(N__60890));
    Odrv4 I__11579 (
            .O(N__60893),
            .I(\quad_counter0.n2610 ));
    Odrv4 I__11578 (
            .O(N__60890),
            .I(\quad_counter0.n2610 ));
    InMux I__11577 (
            .O(N__60885),
            .I(\quad_counter0.n30280 ));
    InMux I__11576 (
            .O(N__60882),
            .I(N__60878));
    InMux I__11575 (
            .O(N__60881),
            .I(N__60875));
    LocalMux I__11574 (
            .O(N__60878),
            .I(N__60870));
    LocalMux I__11573 (
            .O(N__60875),
            .I(N__60870));
    Span4Mux_v I__11572 (
            .O(N__60870),
            .I(N__60866));
    InMux I__11571 (
            .O(N__60869),
            .I(N__60863));
    Odrv4 I__11570 (
            .O(N__60866),
            .I(\quad_counter0.n2609 ));
    LocalMux I__11569 (
            .O(N__60863),
            .I(\quad_counter0.n2609 ));
    InMux I__11568 (
            .O(N__60858),
            .I(\quad_counter0.n30281 ));
    InMux I__11567 (
            .O(N__60855),
            .I(N__60851));
    InMux I__11566 (
            .O(N__60854),
            .I(N__60848));
    LocalMux I__11565 (
            .O(N__60851),
            .I(N__60843));
    LocalMux I__11564 (
            .O(N__60848),
            .I(N__60843));
    Span4Mux_v I__11563 (
            .O(N__60843),
            .I(N__60839));
    InMux I__11562 (
            .O(N__60842),
            .I(N__60836));
    Odrv4 I__11561 (
            .O(N__60839),
            .I(\quad_counter0.n2608 ));
    LocalMux I__11560 (
            .O(N__60836),
            .I(\quad_counter0.n2608 ));
    InMux I__11559 (
            .O(N__60831),
            .I(\quad_counter0.n30282 ));
    InMux I__11558 (
            .O(N__60828),
            .I(N__60823));
    InMux I__11557 (
            .O(N__60827),
            .I(N__60820));
    InMux I__11556 (
            .O(N__60826),
            .I(N__60817));
    LocalMux I__11555 (
            .O(N__60823),
            .I(N__60810));
    LocalMux I__11554 (
            .O(N__60820),
            .I(N__60810));
    LocalMux I__11553 (
            .O(N__60817),
            .I(N__60810));
    Span4Mux_h I__11552 (
            .O(N__60810),
            .I(N__60807));
    Odrv4 I__11551 (
            .O(N__60807),
            .I(\quad_counter0.n2607 ));
    InMux I__11550 (
            .O(N__60804),
            .I(\quad_counter0.n30283 ));
    InMux I__11549 (
            .O(N__60801),
            .I(\quad_counter0.n30284 ));
    InMux I__11548 (
            .O(N__60798),
            .I(N__60794));
    InMux I__11547 (
            .O(N__60797),
            .I(N__60791));
    LocalMux I__11546 (
            .O(N__60794),
            .I(N__60786));
    LocalMux I__11545 (
            .O(N__60791),
            .I(N__60786));
    Span4Mux_h I__11544 (
            .O(N__60786),
            .I(N__60782));
    InMux I__11543 (
            .O(N__60785),
            .I(N__60779));
    Odrv4 I__11542 (
            .O(N__60782),
            .I(\quad_counter0.n2606 ));
    LocalMux I__11541 (
            .O(N__60779),
            .I(\quad_counter0.n2606 ));
    InMux I__11540 (
            .O(N__60774),
            .I(N__60768));
    InMux I__11539 (
            .O(N__60773),
            .I(N__60768));
    LocalMux I__11538 (
            .O(N__60768),
            .I(data_out_frame_9_3));
    CascadeMux I__11537 (
            .O(N__60765),
            .I(\c0.n36161_cascade_ ));
    CascadeMux I__11536 (
            .O(N__60762),
            .I(\c0.n36164_cascade_ ));
    InMux I__11535 (
            .O(N__60759),
            .I(N__60756));
    LocalMux I__11534 (
            .O(N__60756),
            .I(n36082));
    InMux I__11533 (
            .O(N__60753),
            .I(N__60749));
    InMux I__11532 (
            .O(N__60752),
            .I(N__60746));
    LocalMux I__11531 (
            .O(N__60749),
            .I(N__60741));
    LocalMux I__11530 (
            .O(N__60746),
            .I(N__60741));
    Span4Mux_h I__11529 (
            .O(N__60741),
            .I(N__60737));
    InMux I__11528 (
            .O(N__60740),
            .I(N__60734));
    Odrv4 I__11527 (
            .O(N__60737),
            .I(\quad_counter0.n2618 ));
    LocalMux I__11526 (
            .O(N__60734),
            .I(\quad_counter0.n2618 ));
    InMux I__11525 (
            .O(N__60729),
            .I(\quad_counter0.n30272 ));
    InMux I__11524 (
            .O(N__60726),
            .I(N__60722));
    InMux I__11523 (
            .O(N__60725),
            .I(N__60719));
    LocalMux I__11522 (
            .O(N__60722),
            .I(N__60716));
    LocalMux I__11521 (
            .O(N__60719),
            .I(N__60713));
    Span4Mux_v I__11520 (
            .O(N__60716),
            .I(N__60707));
    Span4Mux_v I__11519 (
            .O(N__60713),
            .I(N__60707));
    InMux I__11518 (
            .O(N__60712),
            .I(N__60704));
    Odrv4 I__11517 (
            .O(N__60707),
            .I(\quad_counter0.n2617 ));
    LocalMux I__11516 (
            .O(N__60704),
            .I(\quad_counter0.n2617 ));
    InMux I__11515 (
            .O(N__60699),
            .I(\quad_counter0.n30273 ));
    InMux I__11514 (
            .O(N__60696),
            .I(N__60692));
    InMux I__11513 (
            .O(N__60695),
            .I(N__60689));
    LocalMux I__11512 (
            .O(N__60692),
            .I(N__60684));
    LocalMux I__11511 (
            .O(N__60689),
            .I(N__60684));
    Span4Mux_v I__11510 (
            .O(N__60684),
            .I(N__60680));
    InMux I__11509 (
            .O(N__60683),
            .I(N__60677));
    Odrv4 I__11508 (
            .O(N__60680),
            .I(\quad_counter0.n2616 ));
    LocalMux I__11507 (
            .O(N__60677),
            .I(\quad_counter0.n2616 ));
    InMux I__11506 (
            .O(N__60672),
            .I(\quad_counter0.n30274 ));
    InMux I__11505 (
            .O(N__60669),
            .I(N__60665));
    InMux I__11504 (
            .O(N__60668),
            .I(N__60662));
    LocalMux I__11503 (
            .O(N__60665),
            .I(N__60656));
    LocalMux I__11502 (
            .O(N__60662),
            .I(N__60656));
    CascadeMux I__11501 (
            .O(N__60661),
            .I(N__60653));
    Span4Mux_h I__11500 (
            .O(N__60656),
            .I(N__60650));
    InMux I__11499 (
            .O(N__60653),
            .I(N__60647));
    Odrv4 I__11498 (
            .O(N__60650),
            .I(\quad_counter0.n2615 ));
    LocalMux I__11497 (
            .O(N__60647),
            .I(\quad_counter0.n2615 ));
    InMux I__11496 (
            .O(N__60642),
            .I(\quad_counter0.n30275 ));
    InMux I__11495 (
            .O(N__60639),
            .I(N__60635));
    InMux I__11494 (
            .O(N__60638),
            .I(N__60632));
    LocalMux I__11493 (
            .O(N__60635),
            .I(N__60627));
    LocalMux I__11492 (
            .O(N__60632),
            .I(N__60627));
    Span4Mux_h I__11491 (
            .O(N__60627),
            .I(N__60623));
    InMux I__11490 (
            .O(N__60626),
            .I(N__60620));
    Odrv4 I__11489 (
            .O(N__60623),
            .I(\quad_counter0.n2614 ));
    LocalMux I__11488 (
            .O(N__60620),
            .I(\quad_counter0.n2614 ));
    InMux I__11487 (
            .O(N__60615),
            .I(\quad_counter0.n30276 ));
    InMux I__11486 (
            .O(N__60612),
            .I(N__60607));
    InMux I__11485 (
            .O(N__60611),
            .I(N__60604));
    InMux I__11484 (
            .O(N__60610),
            .I(N__60601));
    LocalMux I__11483 (
            .O(N__60607),
            .I(N__60596));
    LocalMux I__11482 (
            .O(N__60604),
            .I(N__60596));
    LocalMux I__11481 (
            .O(N__60601),
            .I(N__60593));
    Span4Mux_v I__11480 (
            .O(N__60596),
            .I(N__60590));
    Span4Mux_h I__11479 (
            .O(N__60593),
            .I(N__60587));
    Odrv4 I__11478 (
            .O(N__60590),
            .I(\quad_counter0.n2613 ));
    Odrv4 I__11477 (
            .O(N__60587),
            .I(\quad_counter0.n2613 ));
    InMux I__11476 (
            .O(N__60582),
            .I(\quad_counter0.n30277 ));
    InMux I__11475 (
            .O(N__60579),
            .I(N__60575));
    InMux I__11474 (
            .O(N__60578),
            .I(N__60572));
    LocalMux I__11473 (
            .O(N__60575),
            .I(N__60566));
    LocalMux I__11472 (
            .O(N__60572),
            .I(N__60566));
    CascadeMux I__11471 (
            .O(N__60571),
            .I(N__60563));
    Span4Mux_h I__11470 (
            .O(N__60566),
            .I(N__60560));
    InMux I__11469 (
            .O(N__60563),
            .I(N__60557));
    Odrv4 I__11468 (
            .O(N__60560),
            .I(\quad_counter0.n2612 ));
    LocalMux I__11467 (
            .O(N__60557),
            .I(\quad_counter0.n2612 ));
    InMux I__11466 (
            .O(N__60552),
            .I(\quad_counter0.n30278 ));
    InMux I__11465 (
            .O(N__60549),
            .I(N__60545));
    InMux I__11464 (
            .O(N__60548),
            .I(N__60542));
    LocalMux I__11463 (
            .O(N__60545),
            .I(N__60537));
    LocalMux I__11462 (
            .O(N__60542),
            .I(N__60537));
    Span4Mux_h I__11461 (
            .O(N__60537),
            .I(N__60533));
    InMux I__11460 (
            .O(N__60536),
            .I(N__60530));
    Odrv4 I__11459 (
            .O(N__60533),
            .I(\quad_counter0.n2611 ));
    LocalMux I__11458 (
            .O(N__60530),
            .I(\quad_counter0.n2611 ));
    InMux I__11457 (
            .O(N__60525),
            .I(bfn_17_14_0_));
    InMux I__11456 (
            .O(N__60522),
            .I(\quad_counter0.n30164 ));
    InMux I__11455 (
            .O(N__60519),
            .I(N__60515));
    InMux I__11454 (
            .O(N__60518),
            .I(N__60512));
    LocalMux I__11453 (
            .O(N__60515),
            .I(N__60506));
    LocalMux I__11452 (
            .O(N__60512),
            .I(N__60506));
    InMux I__11451 (
            .O(N__60511),
            .I(N__60503));
    Span4Mux_h I__11450 (
            .O(N__60506),
            .I(N__60499));
    LocalMux I__11449 (
            .O(N__60503),
            .I(N__60496));
    InMux I__11448 (
            .O(N__60502),
            .I(N__60493));
    Span4Mux_h I__11447 (
            .O(N__60499),
            .I(N__60490));
    Span12Mux_h I__11446 (
            .O(N__60496),
            .I(N__60487));
    LocalMux I__11445 (
            .O(N__60493),
            .I(\quad_counter0.millisecond_counter_26 ));
    Odrv4 I__11444 (
            .O(N__60490),
            .I(\quad_counter0.millisecond_counter_26 ));
    Odrv12 I__11443 (
            .O(N__60487),
            .I(\quad_counter0.millisecond_counter_26 ));
    InMux I__11442 (
            .O(N__60480),
            .I(\quad_counter0.n30165 ));
    InMux I__11441 (
            .O(N__60477),
            .I(N__60472));
    InMux I__11440 (
            .O(N__60476),
            .I(N__60469));
    InMux I__11439 (
            .O(N__60475),
            .I(N__60466));
    LocalMux I__11438 (
            .O(N__60472),
            .I(N__60461));
    LocalMux I__11437 (
            .O(N__60469),
            .I(N__60461));
    LocalMux I__11436 (
            .O(N__60466),
            .I(N__60458));
    Span4Mux_h I__11435 (
            .O(N__60461),
            .I(N__60454));
    Span4Mux_v I__11434 (
            .O(N__60458),
            .I(N__60451));
    InMux I__11433 (
            .O(N__60457),
            .I(N__60448));
    Span4Mux_v I__11432 (
            .O(N__60454),
            .I(N__60443));
    Span4Mux_h I__11431 (
            .O(N__60451),
            .I(N__60443));
    LocalMux I__11430 (
            .O(N__60448),
            .I(\quad_counter0.millisecond_counter_27 ));
    Odrv4 I__11429 (
            .O(N__60443),
            .I(\quad_counter0.millisecond_counter_27 ));
    InMux I__11428 (
            .O(N__60438),
            .I(\quad_counter0.n30166 ));
    CascadeMux I__11427 (
            .O(N__60435),
            .I(N__60430));
    InMux I__11426 (
            .O(N__60434),
            .I(N__60427));
    InMux I__11425 (
            .O(N__60433),
            .I(N__60424));
    InMux I__11424 (
            .O(N__60430),
            .I(N__60421));
    LocalMux I__11423 (
            .O(N__60427),
            .I(N__60416));
    LocalMux I__11422 (
            .O(N__60424),
            .I(N__60416));
    LocalMux I__11421 (
            .O(N__60421),
            .I(N__60413));
    Span4Mux_v I__11420 (
            .O(N__60416),
            .I(N__60407));
    Span4Mux_h I__11419 (
            .O(N__60413),
            .I(N__60407));
    InMux I__11418 (
            .O(N__60412),
            .I(N__60404));
    Span4Mux_h I__11417 (
            .O(N__60407),
            .I(N__60401));
    LocalMux I__11416 (
            .O(N__60404),
            .I(\quad_counter0.millisecond_counter_28 ));
    Odrv4 I__11415 (
            .O(N__60401),
            .I(\quad_counter0.millisecond_counter_28 ));
    InMux I__11414 (
            .O(N__60396),
            .I(\quad_counter0.n30167 ));
    InMux I__11413 (
            .O(N__60393),
            .I(N__60388));
    InMux I__11412 (
            .O(N__60392),
            .I(N__60385));
    InMux I__11411 (
            .O(N__60391),
            .I(N__60382));
    LocalMux I__11410 (
            .O(N__60388),
            .I(N__60379));
    LocalMux I__11409 (
            .O(N__60385),
            .I(N__60376));
    LocalMux I__11408 (
            .O(N__60382),
            .I(N__60373));
    Span4Mux_v I__11407 (
            .O(N__60379),
            .I(N__60365));
    Span4Mux_v I__11406 (
            .O(N__60376),
            .I(N__60365));
    Span4Mux_h I__11405 (
            .O(N__60373),
            .I(N__60365));
    InMux I__11404 (
            .O(N__60372),
            .I(N__60362));
    Span4Mux_h I__11403 (
            .O(N__60365),
            .I(N__60359));
    LocalMux I__11402 (
            .O(N__60362),
            .I(\quad_counter0.millisecond_counter_29 ));
    Odrv4 I__11401 (
            .O(N__60359),
            .I(\quad_counter0.millisecond_counter_29 ));
    InMux I__11400 (
            .O(N__60354),
            .I(\quad_counter0.n30168 ));
    InMux I__11399 (
            .O(N__60351),
            .I(N__60346));
    InMux I__11398 (
            .O(N__60350),
            .I(N__60343));
    InMux I__11397 (
            .O(N__60349),
            .I(N__60340));
    LocalMux I__11396 (
            .O(N__60346),
            .I(N__60335));
    LocalMux I__11395 (
            .O(N__60343),
            .I(N__60335));
    LocalMux I__11394 (
            .O(N__60340),
            .I(N__60332));
    Span4Mux_v I__11393 (
            .O(N__60335),
            .I(N__60326));
    Span4Mux_h I__11392 (
            .O(N__60332),
            .I(N__60326));
    InMux I__11391 (
            .O(N__60331),
            .I(N__60323));
    Span4Mux_h I__11390 (
            .O(N__60326),
            .I(N__60320));
    LocalMux I__11389 (
            .O(N__60323),
            .I(\quad_counter0.millisecond_counter_30 ));
    Odrv4 I__11388 (
            .O(N__60320),
            .I(\quad_counter0.millisecond_counter_30 ));
    InMux I__11387 (
            .O(N__60315),
            .I(\quad_counter0.n30169 ));
    InMux I__11386 (
            .O(N__60312),
            .I(\quad_counter0.n30170 ));
    InMux I__11385 (
            .O(N__60309),
            .I(N__60304));
    InMux I__11384 (
            .O(N__60308),
            .I(N__60301));
    InMux I__11383 (
            .O(N__60307),
            .I(N__60298));
    LocalMux I__11382 (
            .O(N__60304),
            .I(N__60293));
    LocalMux I__11381 (
            .O(N__60301),
            .I(N__60293));
    LocalMux I__11380 (
            .O(N__60298),
            .I(N__60290));
    Span4Mux_v I__11379 (
            .O(N__60293),
            .I(N__60284));
    Span4Mux_h I__11378 (
            .O(N__60290),
            .I(N__60284));
    InMux I__11377 (
            .O(N__60289),
            .I(N__60281));
    Span4Mux_h I__11376 (
            .O(N__60284),
            .I(N__60278));
    LocalMux I__11375 (
            .O(N__60281),
            .I(\quad_counter0.millisecond_counter_31 ));
    Odrv4 I__11374 (
            .O(N__60278),
            .I(\quad_counter0.millisecond_counter_31 ));
    InMux I__11373 (
            .O(N__60273),
            .I(N__60269));
    InMux I__11372 (
            .O(N__60272),
            .I(N__60266));
    LocalMux I__11371 (
            .O(N__60269),
            .I(N__60263));
    LocalMux I__11370 (
            .O(N__60266),
            .I(N__60260));
    Span12Mux_v I__11369 (
            .O(N__60263),
            .I(N__60257));
    Odrv4 I__11368 (
            .O(N__60260),
            .I(n34523));
    Odrv12 I__11367 (
            .O(N__60257),
            .I(n34523));
    InMux I__11366 (
            .O(N__60252),
            .I(N__60249));
    LocalMux I__11365 (
            .O(N__60249),
            .I(N__60245));
    InMux I__11364 (
            .O(N__60248),
            .I(N__60242));
    Span12Mux_v I__11363 (
            .O(N__60245),
            .I(N__60239));
    LocalMux I__11362 (
            .O(N__60242),
            .I(count_prev_0));
    Odrv12 I__11361 (
            .O(N__60239),
            .I(count_prev_0));
    InMux I__11360 (
            .O(N__60234),
            .I(N__60230));
    InMux I__11359 (
            .O(N__60233),
            .I(N__60227));
    LocalMux I__11358 (
            .O(N__60230),
            .I(N__60221));
    LocalMux I__11357 (
            .O(N__60227),
            .I(N__60221));
    CascadeMux I__11356 (
            .O(N__60226),
            .I(N__60218));
    Span4Mux_h I__11355 (
            .O(N__60221),
            .I(N__60215));
    InMux I__11354 (
            .O(N__60218),
            .I(N__60212));
    Odrv4 I__11353 (
            .O(N__60215),
            .I(\quad_counter0.n2619 ));
    LocalMux I__11352 (
            .O(N__60212),
            .I(\quad_counter0.n2619 ));
    InMux I__11351 (
            .O(N__60207),
            .I(bfn_17_13_0_));
    InMux I__11350 (
            .O(N__60204),
            .I(N__60199));
    InMux I__11349 (
            .O(N__60203),
            .I(N__60196));
    InMux I__11348 (
            .O(N__60202),
            .I(N__60192));
    LocalMux I__11347 (
            .O(N__60199),
            .I(N__60189));
    LocalMux I__11346 (
            .O(N__60196),
            .I(N__60186));
    InMux I__11345 (
            .O(N__60195),
            .I(N__60183));
    LocalMux I__11344 (
            .O(N__60192),
            .I(N__60180));
    Span4Mux_h I__11343 (
            .O(N__60189),
            .I(N__60177));
    Span4Mux_h I__11342 (
            .O(N__60186),
            .I(N__60174));
    LocalMux I__11341 (
            .O(N__60183),
            .I(N__60169));
    Span4Mux_v I__11340 (
            .O(N__60180),
            .I(N__60169));
    Odrv4 I__11339 (
            .O(N__60177),
            .I(\quad_counter0.millisecond_counter_17 ));
    Odrv4 I__11338 (
            .O(N__60174),
            .I(\quad_counter0.millisecond_counter_17 ));
    Odrv4 I__11337 (
            .O(N__60169),
            .I(\quad_counter0.millisecond_counter_17 ));
    InMux I__11336 (
            .O(N__60162),
            .I(\quad_counter0.n30156 ));
    InMux I__11335 (
            .O(N__60159),
            .I(\quad_counter0.n30157 ));
    InMux I__11334 (
            .O(N__60156),
            .I(\quad_counter0.n30158 ));
    InMux I__11333 (
            .O(N__60153),
            .I(\quad_counter0.n30159 ));
    InMux I__11332 (
            .O(N__60150),
            .I(\quad_counter0.n30160 ));
    InMux I__11331 (
            .O(N__60147),
            .I(N__60142));
    InMux I__11330 (
            .O(N__60146),
            .I(N__60139));
    InMux I__11329 (
            .O(N__60145),
            .I(N__60136));
    LocalMux I__11328 (
            .O(N__60142),
            .I(N__60130));
    LocalMux I__11327 (
            .O(N__60139),
            .I(N__60130));
    LocalMux I__11326 (
            .O(N__60136),
            .I(N__60127));
    InMux I__11325 (
            .O(N__60135),
            .I(N__60124));
    Span4Mux_h I__11324 (
            .O(N__60130),
            .I(N__60119));
    Span4Mux_h I__11323 (
            .O(N__60127),
            .I(N__60119));
    LocalMux I__11322 (
            .O(N__60124),
            .I(N__60114));
    Span4Mux_v I__11321 (
            .O(N__60119),
            .I(N__60114));
    Odrv4 I__11320 (
            .O(N__60114),
            .I(\quad_counter0.millisecond_counter_22 ));
    InMux I__11319 (
            .O(N__60111),
            .I(\quad_counter0.n30161 ));
    CascadeMux I__11318 (
            .O(N__60108),
            .I(N__60103));
    InMux I__11317 (
            .O(N__60107),
            .I(N__60100));
    InMux I__11316 (
            .O(N__60106),
            .I(N__60097));
    InMux I__11315 (
            .O(N__60103),
            .I(N__60094));
    LocalMux I__11314 (
            .O(N__60100),
            .I(N__60088));
    LocalMux I__11313 (
            .O(N__60097),
            .I(N__60088));
    LocalMux I__11312 (
            .O(N__60094),
            .I(N__60085));
    InMux I__11311 (
            .O(N__60093),
            .I(N__60082));
    Span4Mux_h I__11310 (
            .O(N__60088),
            .I(N__60079));
    Span12Mux_s9_v I__11309 (
            .O(N__60085),
            .I(N__60076));
    LocalMux I__11308 (
            .O(N__60082),
            .I(N__60071));
    Span4Mux_v I__11307 (
            .O(N__60079),
            .I(N__60071));
    Odrv12 I__11306 (
            .O(N__60076),
            .I(\quad_counter0.millisecond_counter_23 ));
    Odrv4 I__11305 (
            .O(N__60071),
            .I(\quad_counter0.millisecond_counter_23 ));
    InMux I__11304 (
            .O(N__60066),
            .I(\quad_counter0.n30162 ));
    InMux I__11303 (
            .O(N__60063),
            .I(N__60058));
    InMux I__11302 (
            .O(N__60062),
            .I(N__60055));
    InMux I__11301 (
            .O(N__60061),
            .I(N__60052));
    LocalMux I__11300 (
            .O(N__60058),
            .I(N__60045));
    LocalMux I__11299 (
            .O(N__60055),
            .I(N__60045));
    LocalMux I__11298 (
            .O(N__60052),
            .I(N__60045));
    Span4Mux_v I__11297 (
            .O(N__60045),
            .I(N__60041));
    InMux I__11296 (
            .O(N__60044),
            .I(N__60038));
    Span4Mux_h I__11295 (
            .O(N__60041),
            .I(N__60035));
    LocalMux I__11294 (
            .O(N__60038),
            .I(\quad_counter0.millisecond_counter_24 ));
    Odrv4 I__11293 (
            .O(N__60035),
            .I(\quad_counter0.millisecond_counter_24 ));
    InMux I__11292 (
            .O(N__60030),
            .I(bfn_17_11_0_));
    InMux I__11291 (
            .O(N__60027),
            .I(N__60022));
    InMux I__11290 (
            .O(N__60026),
            .I(N__60019));
    InMux I__11289 (
            .O(N__60025),
            .I(N__60016));
    LocalMux I__11288 (
            .O(N__60022),
            .I(N__60011));
    LocalMux I__11287 (
            .O(N__60019),
            .I(N__60011));
    LocalMux I__11286 (
            .O(N__60016),
            .I(N__60008));
    Span4Mux_h I__11285 (
            .O(N__60011),
            .I(N__60004));
    Span4Mux_h I__11284 (
            .O(N__60008),
            .I(N__60001));
    InMux I__11283 (
            .O(N__60007),
            .I(N__59998));
    Span4Mux_h I__11282 (
            .O(N__60004),
            .I(N__59995));
    Span4Mux_h I__11281 (
            .O(N__60001),
            .I(N__59992));
    LocalMux I__11280 (
            .O(N__59998),
            .I(\quad_counter0.millisecond_counter_25 ));
    Odrv4 I__11279 (
            .O(N__59995),
            .I(\quad_counter0.millisecond_counter_25 ));
    Odrv4 I__11278 (
            .O(N__59992),
            .I(\quad_counter0.millisecond_counter_25 ));
    InMux I__11277 (
            .O(N__59985),
            .I(N__59980));
    InMux I__11276 (
            .O(N__59984),
            .I(N__59976));
    InMux I__11275 (
            .O(N__59983),
            .I(N__59973));
    LocalMux I__11274 (
            .O(N__59980),
            .I(N__59970));
    InMux I__11273 (
            .O(N__59979),
            .I(N__59967));
    LocalMux I__11272 (
            .O(N__59976),
            .I(N__59962));
    LocalMux I__11271 (
            .O(N__59973),
            .I(N__59962));
    Span4Mux_v I__11270 (
            .O(N__59970),
            .I(N__59959));
    LocalMux I__11269 (
            .O(N__59967),
            .I(\quad_counter0.millisecond_counter_8 ));
    Odrv12 I__11268 (
            .O(N__59962),
            .I(\quad_counter0.millisecond_counter_8 ));
    Odrv4 I__11267 (
            .O(N__59959),
            .I(\quad_counter0.millisecond_counter_8 ));
    InMux I__11266 (
            .O(N__59952),
            .I(bfn_17_9_0_));
    InMux I__11265 (
            .O(N__59949),
            .I(N__59943));
    InMux I__11264 (
            .O(N__59948),
            .I(N__59940));
    InMux I__11263 (
            .O(N__59947),
            .I(N__59937));
    InMux I__11262 (
            .O(N__59946),
            .I(N__59934));
    LocalMux I__11261 (
            .O(N__59943),
            .I(N__59929));
    LocalMux I__11260 (
            .O(N__59940),
            .I(N__59929));
    LocalMux I__11259 (
            .O(N__59937),
            .I(N__59926));
    LocalMux I__11258 (
            .O(N__59934),
            .I(\quad_counter0.millisecond_counter_9 ));
    Odrv4 I__11257 (
            .O(N__59929),
            .I(\quad_counter0.millisecond_counter_9 ));
    Odrv12 I__11256 (
            .O(N__59926),
            .I(\quad_counter0.millisecond_counter_9 ));
    InMux I__11255 (
            .O(N__59919),
            .I(\quad_counter0.n30148 ));
    InMux I__11254 (
            .O(N__59916),
            .I(N__59910));
    InMux I__11253 (
            .O(N__59915),
            .I(N__59907));
    InMux I__11252 (
            .O(N__59914),
            .I(N__59904));
    InMux I__11251 (
            .O(N__59913),
            .I(N__59901));
    LocalMux I__11250 (
            .O(N__59910),
            .I(N__59894));
    LocalMux I__11249 (
            .O(N__59907),
            .I(N__59894));
    LocalMux I__11248 (
            .O(N__59904),
            .I(N__59894));
    LocalMux I__11247 (
            .O(N__59901),
            .I(N__59889));
    Span4Mux_h I__11246 (
            .O(N__59894),
            .I(N__59889));
    Odrv4 I__11245 (
            .O(N__59889),
            .I(\quad_counter0.millisecond_counter_10 ));
    InMux I__11244 (
            .O(N__59886),
            .I(\quad_counter0.n30149 ));
    InMux I__11243 (
            .O(N__59883),
            .I(N__59877));
    InMux I__11242 (
            .O(N__59882),
            .I(N__59874));
    InMux I__11241 (
            .O(N__59881),
            .I(N__59871));
    InMux I__11240 (
            .O(N__59880),
            .I(N__59868));
    LocalMux I__11239 (
            .O(N__59877),
            .I(N__59861));
    LocalMux I__11238 (
            .O(N__59874),
            .I(N__59861));
    LocalMux I__11237 (
            .O(N__59871),
            .I(N__59861));
    LocalMux I__11236 (
            .O(N__59868),
            .I(\quad_counter0.millisecond_counter_11 ));
    Odrv12 I__11235 (
            .O(N__59861),
            .I(\quad_counter0.millisecond_counter_11 ));
    InMux I__11234 (
            .O(N__59856),
            .I(\quad_counter0.n30150 ));
    InMux I__11233 (
            .O(N__59853),
            .I(N__59849));
    InMux I__11232 (
            .O(N__59852),
            .I(N__59846));
    LocalMux I__11231 (
            .O(N__59849),
            .I(N__59840));
    LocalMux I__11230 (
            .O(N__59846),
            .I(N__59840));
    InMux I__11229 (
            .O(N__59845),
            .I(N__59837));
    Span4Mux_h I__11228 (
            .O(N__59840),
            .I(N__59833));
    LocalMux I__11227 (
            .O(N__59837),
            .I(N__59830));
    InMux I__11226 (
            .O(N__59836),
            .I(N__59827));
    Span4Mux_h I__11225 (
            .O(N__59833),
            .I(N__59824));
    Span12Mux_v I__11224 (
            .O(N__59830),
            .I(N__59821));
    LocalMux I__11223 (
            .O(N__59827),
            .I(\quad_counter0.millisecond_counter_12 ));
    Odrv4 I__11222 (
            .O(N__59824),
            .I(\quad_counter0.millisecond_counter_12 ));
    Odrv12 I__11221 (
            .O(N__59821),
            .I(\quad_counter0.millisecond_counter_12 ));
    InMux I__11220 (
            .O(N__59814),
            .I(\quad_counter0.n30151 ));
    InMux I__11219 (
            .O(N__59811),
            .I(N__59807));
    InMux I__11218 (
            .O(N__59810),
            .I(N__59804));
    LocalMux I__11217 (
            .O(N__59807),
            .I(N__59799));
    LocalMux I__11216 (
            .O(N__59804),
            .I(N__59799));
    Span4Mux_h I__11215 (
            .O(N__59799),
            .I(N__59796));
    Span4Mux_v I__11214 (
            .O(N__59796),
            .I(N__59791));
    InMux I__11213 (
            .O(N__59795),
            .I(N__59788));
    InMux I__11212 (
            .O(N__59794),
            .I(N__59785));
    Span4Mux_h I__11211 (
            .O(N__59791),
            .I(N__59782));
    LocalMux I__11210 (
            .O(N__59788),
            .I(N__59779));
    LocalMux I__11209 (
            .O(N__59785),
            .I(\quad_counter0.millisecond_counter_13 ));
    Odrv4 I__11208 (
            .O(N__59782),
            .I(\quad_counter0.millisecond_counter_13 ));
    Odrv12 I__11207 (
            .O(N__59779),
            .I(\quad_counter0.millisecond_counter_13 ));
    InMux I__11206 (
            .O(N__59772),
            .I(\quad_counter0.n30152 ));
    InMux I__11205 (
            .O(N__59769),
            .I(N__59764));
    InMux I__11204 (
            .O(N__59768),
            .I(N__59761));
    InMux I__11203 (
            .O(N__59767),
            .I(N__59758));
    LocalMux I__11202 (
            .O(N__59764),
            .I(N__59755));
    LocalMux I__11201 (
            .O(N__59761),
            .I(N__59750));
    LocalMux I__11200 (
            .O(N__59758),
            .I(N__59750));
    Span4Mux_h I__11199 (
            .O(N__59755),
            .I(N__59747));
    Sp12to4 I__11198 (
            .O(N__59750),
            .I(N__59743));
    Span4Mux_h I__11197 (
            .O(N__59747),
            .I(N__59740));
    InMux I__11196 (
            .O(N__59746),
            .I(N__59737));
    Span12Mux_h I__11195 (
            .O(N__59743),
            .I(N__59734));
    Span4Mux_v I__11194 (
            .O(N__59740),
            .I(N__59731));
    LocalMux I__11193 (
            .O(N__59737),
            .I(\quad_counter0.millisecond_counter_14 ));
    Odrv12 I__11192 (
            .O(N__59734),
            .I(\quad_counter0.millisecond_counter_14 ));
    Odrv4 I__11191 (
            .O(N__59731),
            .I(\quad_counter0.millisecond_counter_14 ));
    InMux I__11190 (
            .O(N__59724),
            .I(\quad_counter0.n30153 ));
    InMux I__11189 (
            .O(N__59721),
            .I(N__59716));
    InMux I__11188 (
            .O(N__59720),
            .I(N__59713));
    InMux I__11187 (
            .O(N__59719),
            .I(N__59710));
    LocalMux I__11186 (
            .O(N__59716),
            .I(N__59705));
    LocalMux I__11185 (
            .O(N__59713),
            .I(N__59705));
    LocalMux I__11184 (
            .O(N__59710),
            .I(N__59702));
    Span4Mux_h I__11183 (
            .O(N__59705),
            .I(N__59699));
    Span4Mux_h I__11182 (
            .O(N__59702),
            .I(N__59696));
    Span4Mux_h I__11181 (
            .O(N__59699),
            .I(N__59692));
    Span4Mux_h I__11180 (
            .O(N__59696),
            .I(N__59689));
    InMux I__11179 (
            .O(N__59695),
            .I(N__59686));
    Span4Mux_v I__11178 (
            .O(N__59692),
            .I(N__59683));
    Span4Mux_v I__11177 (
            .O(N__59689),
            .I(N__59680));
    LocalMux I__11176 (
            .O(N__59686),
            .I(\quad_counter0.millisecond_counter_15 ));
    Odrv4 I__11175 (
            .O(N__59683),
            .I(\quad_counter0.millisecond_counter_15 ));
    Odrv4 I__11174 (
            .O(N__59680),
            .I(\quad_counter0.millisecond_counter_15 ));
    InMux I__11173 (
            .O(N__59673),
            .I(\quad_counter0.n30154 ));
    InMux I__11172 (
            .O(N__59670),
            .I(N__59666));
    InMux I__11171 (
            .O(N__59669),
            .I(N__59663));
    LocalMux I__11170 (
            .O(N__59666),
            .I(N__59656));
    LocalMux I__11169 (
            .O(N__59663),
            .I(N__59656));
    InMux I__11168 (
            .O(N__59662),
            .I(N__59653));
    InMux I__11167 (
            .O(N__59661),
            .I(N__59650));
    Span4Mux_v I__11166 (
            .O(N__59656),
            .I(N__59647));
    LocalMux I__11165 (
            .O(N__59653),
            .I(N__59644));
    LocalMux I__11164 (
            .O(N__59650),
            .I(N__59639));
    Span4Mux_h I__11163 (
            .O(N__59647),
            .I(N__59639));
    Span4Mux_h I__11162 (
            .O(N__59644),
            .I(N__59636));
    Odrv4 I__11161 (
            .O(N__59639),
            .I(\quad_counter0.millisecond_counter_16 ));
    Odrv4 I__11160 (
            .O(N__59636),
            .I(\quad_counter0.millisecond_counter_16 ));
    InMux I__11159 (
            .O(N__59631),
            .I(bfn_17_10_0_));
    InMux I__11158 (
            .O(N__59628),
            .I(N__59624));
    InMux I__11157 (
            .O(N__59627),
            .I(N__59621));
    LocalMux I__11156 (
            .O(N__59624),
            .I(\quad_counter0.millisecond_counter_0 ));
    LocalMux I__11155 (
            .O(N__59621),
            .I(\quad_counter0.millisecond_counter_0 ));
    InMux I__11154 (
            .O(N__59616),
            .I(bfn_17_8_0_));
    CascadeMux I__11153 (
            .O(N__59613),
            .I(N__59610));
    InMux I__11152 (
            .O(N__59610),
            .I(N__59607));
    LocalMux I__11151 (
            .O(N__59607),
            .I(N__59604));
    Span4Mux_v I__11150 (
            .O(N__59604),
            .I(N__59600));
    InMux I__11149 (
            .O(N__59603),
            .I(N__59597));
    Odrv4 I__11148 (
            .O(N__59600),
            .I(\quad_counter0.millisecond_counter_1 ));
    LocalMux I__11147 (
            .O(N__59597),
            .I(\quad_counter0.millisecond_counter_1 ));
    InMux I__11146 (
            .O(N__59592),
            .I(\quad_counter0.n30140 ));
    InMux I__11145 (
            .O(N__59589),
            .I(N__59585));
    InMux I__11144 (
            .O(N__59588),
            .I(N__59582));
    LocalMux I__11143 (
            .O(N__59585),
            .I(\quad_counter0.millisecond_counter_2 ));
    LocalMux I__11142 (
            .O(N__59582),
            .I(\quad_counter0.millisecond_counter_2 ));
    InMux I__11141 (
            .O(N__59577),
            .I(\quad_counter0.n30141 ));
    InMux I__11140 (
            .O(N__59574),
            .I(N__59570));
    InMux I__11139 (
            .O(N__59573),
            .I(N__59567));
    LocalMux I__11138 (
            .O(N__59570),
            .I(N__59564));
    LocalMux I__11137 (
            .O(N__59567),
            .I(\quad_counter0.millisecond_counter_3 ));
    Odrv4 I__11136 (
            .O(N__59564),
            .I(\quad_counter0.millisecond_counter_3 ));
    InMux I__11135 (
            .O(N__59559),
            .I(\quad_counter0.n30142 ));
    InMux I__11134 (
            .O(N__59556),
            .I(N__59552));
    InMux I__11133 (
            .O(N__59555),
            .I(N__59549));
    LocalMux I__11132 (
            .O(N__59552),
            .I(\quad_counter0.millisecond_counter_4 ));
    LocalMux I__11131 (
            .O(N__59549),
            .I(\quad_counter0.millisecond_counter_4 ));
    InMux I__11130 (
            .O(N__59544),
            .I(\quad_counter0.n30143 ));
    InMux I__11129 (
            .O(N__59541),
            .I(N__59538));
    LocalMux I__11128 (
            .O(N__59538),
            .I(N__59535));
    Span4Mux_h I__11127 (
            .O(N__59535),
            .I(N__59531));
    InMux I__11126 (
            .O(N__59534),
            .I(N__59528));
    Odrv4 I__11125 (
            .O(N__59531),
            .I(\quad_counter0.millisecond_counter_5 ));
    LocalMux I__11124 (
            .O(N__59528),
            .I(\quad_counter0.millisecond_counter_5 ));
    InMux I__11123 (
            .O(N__59523),
            .I(\quad_counter0.n30144 ));
    InMux I__11122 (
            .O(N__59520),
            .I(N__59517));
    LocalMux I__11121 (
            .O(N__59517),
            .I(N__59514));
    Span4Mux_v I__11120 (
            .O(N__59514),
            .I(N__59510));
    InMux I__11119 (
            .O(N__59513),
            .I(N__59507));
    Odrv4 I__11118 (
            .O(N__59510),
            .I(\quad_counter0.millisecond_counter_6 ));
    LocalMux I__11117 (
            .O(N__59507),
            .I(\quad_counter0.millisecond_counter_6 ));
    InMux I__11116 (
            .O(N__59502),
            .I(\quad_counter0.n30145 ));
    InMux I__11115 (
            .O(N__59499),
            .I(N__59496));
    LocalMux I__11114 (
            .O(N__59496),
            .I(N__59493));
    Sp12to4 I__11113 (
            .O(N__59493),
            .I(N__59489));
    InMux I__11112 (
            .O(N__59492),
            .I(N__59486));
    Odrv12 I__11111 (
            .O(N__59489),
            .I(\quad_counter0.millisecond_counter_7 ));
    LocalMux I__11110 (
            .O(N__59486),
            .I(\quad_counter0.millisecond_counter_7 ));
    InMux I__11109 (
            .O(N__59481),
            .I(\quad_counter0.n30146 ));
    CascadeMux I__11108 (
            .O(N__59478),
            .I(\quad_counter1.n28257_cascade_ ));
    CascadeMux I__11107 (
            .O(N__59475),
            .I(\quad_counter1.n10_adj_4472_cascade_ ));
    InMux I__11106 (
            .O(N__59472),
            .I(N__59469));
    LocalMux I__11105 (
            .O(N__59469),
            .I(N__59464));
    InMux I__11104 (
            .O(N__59468),
            .I(N__59459));
    InMux I__11103 (
            .O(N__59467),
            .I(N__59459));
    Odrv4 I__11102 (
            .O(N__59464),
            .I(\quad_counter1.B_delayed ));
    LocalMux I__11101 (
            .O(N__59459),
            .I(\quad_counter1.B_delayed ));
    InMux I__11100 (
            .O(N__59454),
            .I(N__59451));
    LocalMux I__11099 (
            .O(N__59451),
            .I(\quad_counter1.A_delayed ));
    CascadeMux I__11098 (
            .O(N__59448),
            .I(N__59443));
    CascadeMux I__11097 (
            .O(N__59447),
            .I(N__59440));
    InMux I__11096 (
            .O(N__59446),
            .I(N__59436));
    InMux I__11095 (
            .O(N__59443),
            .I(N__59433));
    InMux I__11094 (
            .O(N__59440),
            .I(N__59428));
    InMux I__11093 (
            .O(N__59439),
            .I(N__59428));
    LocalMux I__11092 (
            .O(N__59436),
            .I(N__59423));
    LocalMux I__11091 (
            .O(N__59433),
            .I(N__59423));
    LocalMux I__11090 (
            .O(N__59428),
            .I(N__59420));
    Span4Mux_h I__11089 (
            .O(N__59423),
            .I(N__59416));
    Span4Mux_h I__11088 (
            .O(N__59420),
            .I(N__59413));
    InMux I__11087 (
            .O(N__59419),
            .I(N__59410));
    Span4Mux_h I__11086 (
            .O(N__59416),
            .I(N__59407));
    Span4Mux_h I__11085 (
            .O(N__59413),
            .I(N__59404));
    LocalMux I__11084 (
            .O(N__59410),
            .I(A_filtered_adj_4809));
    Odrv4 I__11083 (
            .O(N__59407),
            .I(A_filtered_adj_4809));
    Odrv4 I__11082 (
            .O(N__59404),
            .I(A_filtered_adj_4809));
    InMux I__11081 (
            .O(N__59397),
            .I(N__59394));
    LocalMux I__11080 (
            .O(N__59394),
            .I(N__59390));
    InMux I__11079 (
            .O(N__59393),
            .I(N__59387));
    Span4Mux_h I__11078 (
            .O(N__59390),
            .I(N__59383));
    LocalMux I__11077 (
            .O(N__59387),
            .I(N__59380));
    InMux I__11076 (
            .O(N__59386),
            .I(N__59377));
    Span4Mux_h I__11075 (
            .O(N__59383),
            .I(N__59374));
    Odrv12 I__11074 (
            .O(N__59380),
            .I(B_filtered_adj_4810));
    LocalMux I__11073 (
            .O(N__59377),
            .I(B_filtered_adj_4810));
    Odrv4 I__11072 (
            .O(N__59374),
            .I(B_filtered_adj_4810));
    InMux I__11071 (
            .O(N__59367),
            .I(N__59363));
    InMux I__11070 (
            .O(N__59366),
            .I(N__59359));
    LocalMux I__11069 (
            .O(N__59363),
            .I(N__59356));
    InMux I__11068 (
            .O(N__59362),
            .I(N__59353));
    LocalMux I__11067 (
            .O(N__59359),
            .I(N__59349));
    Span4Mux_h I__11066 (
            .O(N__59356),
            .I(N__59343));
    LocalMux I__11065 (
            .O(N__59353),
            .I(N__59340));
    InMux I__11064 (
            .O(N__59352),
            .I(N__59337));
    Span12Mux_s7_v I__11063 (
            .O(N__59349),
            .I(N__59334));
    InMux I__11062 (
            .O(N__59348),
            .I(N__59327));
    InMux I__11061 (
            .O(N__59347),
            .I(N__59327));
    InMux I__11060 (
            .O(N__59346),
            .I(N__59327));
    Odrv4 I__11059 (
            .O(N__59343),
            .I(\c0.data_in_frame_19_6 ));
    Odrv12 I__11058 (
            .O(N__59340),
            .I(\c0.data_in_frame_19_6 ));
    LocalMux I__11057 (
            .O(N__59337),
            .I(\c0.data_in_frame_19_6 ));
    Odrv12 I__11056 (
            .O(N__59334),
            .I(\c0.data_in_frame_19_6 ));
    LocalMux I__11055 (
            .O(N__59327),
            .I(\c0.data_in_frame_19_6 ));
    InMux I__11054 (
            .O(N__59316),
            .I(N__59312));
    InMux I__11053 (
            .O(N__59315),
            .I(N__59309));
    LocalMux I__11052 (
            .O(N__59312),
            .I(N__59302));
    LocalMux I__11051 (
            .O(N__59309),
            .I(N__59302));
    InMux I__11050 (
            .O(N__59308),
            .I(N__59299));
    InMux I__11049 (
            .O(N__59307),
            .I(N__59296));
    Span4Mux_v I__11048 (
            .O(N__59302),
            .I(N__59293));
    LocalMux I__11047 (
            .O(N__59299),
            .I(N__59288));
    LocalMux I__11046 (
            .O(N__59296),
            .I(N__59288));
    Span4Mux_h I__11045 (
            .O(N__59293),
            .I(N__59283));
    Span4Mux_v I__11044 (
            .O(N__59288),
            .I(N__59283));
    Odrv4 I__11043 (
            .O(N__59283),
            .I(\c0.n6227 ));
    InMux I__11042 (
            .O(N__59280),
            .I(N__59277));
    LocalMux I__11041 (
            .O(N__59277),
            .I(N__59273));
    InMux I__11040 (
            .O(N__59276),
            .I(N__59270));
    Span4Mux_h I__11039 (
            .O(N__59273),
            .I(N__59267));
    LocalMux I__11038 (
            .O(N__59270),
            .I(N__59264));
    Odrv4 I__11037 (
            .O(N__59267),
            .I(\c0.n31444 ));
    Odrv4 I__11036 (
            .O(N__59264),
            .I(\c0.n31444 ));
    InMux I__11035 (
            .O(N__59259),
            .I(N__59256));
    LocalMux I__11034 (
            .O(N__59256),
            .I(\c0.n41_adj_4704 ));
    InMux I__11033 (
            .O(N__59253),
            .I(N__59250));
    LocalMux I__11032 (
            .O(N__59250),
            .I(N__59247));
    Odrv4 I__11031 (
            .O(N__59247),
            .I(\c0.n42_adj_4703 ));
    CascadeMux I__11030 (
            .O(N__59244),
            .I(\c0.n33490_cascade_ ));
    InMux I__11029 (
            .O(N__59241),
            .I(N__59238));
    LocalMux I__11028 (
            .O(N__59238),
            .I(\c0.n46 ));
    CascadeMux I__11027 (
            .O(N__59235),
            .I(\c0.n25_cascade_ ));
    CascadeMux I__11026 (
            .O(N__59232),
            .I(\c0.n31_cascade_ ));
    InMux I__11025 (
            .O(N__59229),
            .I(N__59225));
    InMux I__11024 (
            .O(N__59228),
            .I(N__59221));
    LocalMux I__11023 (
            .O(N__59225),
            .I(N__59217));
    InMux I__11022 (
            .O(N__59224),
            .I(N__59214));
    LocalMux I__11021 (
            .O(N__59221),
            .I(N__59211));
    InMux I__11020 (
            .O(N__59220),
            .I(N__59208));
    Span4Mux_v I__11019 (
            .O(N__59217),
            .I(N__59203));
    LocalMux I__11018 (
            .O(N__59214),
            .I(N__59203));
    Span4Mux_h I__11017 (
            .O(N__59211),
            .I(N__59198));
    LocalMux I__11016 (
            .O(N__59208),
            .I(N__59198));
    Span4Mux_h I__11015 (
            .O(N__59203),
            .I(N__59195));
    Span4Mux_h I__11014 (
            .O(N__59198),
            .I(N__59192));
    Span4Mux_h I__11013 (
            .O(N__59195),
            .I(N__59189));
    Odrv4 I__11012 (
            .O(N__59192),
            .I(\c0.n18861 ));
    Odrv4 I__11011 (
            .O(N__59189),
            .I(\c0.n18861 ));
    InMux I__11010 (
            .O(N__59184),
            .I(N__59181));
    LocalMux I__11009 (
            .O(N__59181),
            .I(N__59178));
    Span4Mux_v I__11008 (
            .O(N__59178),
            .I(N__59174));
    InMux I__11007 (
            .O(N__59177),
            .I(N__59171));
    Span4Mux_v I__11006 (
            .O(N__59174),
            .I(N__59168));
    LocalMux I__11005 (
            .O(N__59171),
            .I(N__59165));
    Odrv4 I__11004 (
            .O(N__59168),
            .I(\c0.n33913 ));
    Odrv4 I__11003 (
            .O(N__59165),
            .I(\c0.n33913 ));
    InMux I__11002 (
            .O(N__59160),
            .I(N__59157));
    LocalMux I__11001 (
            .O(N__59157),
            .I(N__59154));
    Odrv4 I__11000 (
            .O(N__59154),
            .I(\c0.n33969 ));
    CascadeMux I__10999 (
            .O(N__59151),
            .I(N__59147));
    InMux I__10998 (
            .O(N__59150),
            .I(N__59144));
    InMux I__10997 (
            .O(N__59147),
            .I(N__59141));
    LocalMux I__10996 (
            .O(N__59144),
            .I(N__59138));
    LocalMux I__10995 (
            .O(N__59141),
            .I(N__59134));
    Span4Mux_h I__10994 (
            .O(N__59138),
            .I(N__59131));
    InMux I__10993 (
            .O(N__59137),
            .I(N__59128));
    Odrv4 I__10992 (
            .O(N__59134),
            .I(\c0.data_in_frame_16_5 ));
    Odrv4 I__10991 (
            .O(N__59131),
            .I(\c0.data_in_frame_16_5 ));
    LocalMux I__10990 (
            .O(N__59128),
            .I(\c0.data_in_frame_16_5 ));
    InMux I__10989 (
            .O(N__59121),
            .I(N__59118));
    LocalMux I__10988 (
            .O(N__59118),
            .I(N__59115));
    Span4Mux_h I__10987 (
            .O(N__59115),
            .I(N__59112));
    Odrv4 I__10986 (
            .O(N__59112),
            .I(\c0.n18228 ));
    InMux I__10985 (
            .O(N__59109),
            .I(N__59105));
    InMux I__10984 (
            .O(N__59108),
            .I(N__59102));
    LocalMux I__10983 (
            .O(N__59105),
            .I(N__59099));
    LocalMux I__10982 (
            .O(N__59102),
            .I(N__59096));
    Odrv4 I__10981 (
            .O(N__59099),
            .I(\c0.n33957 ));
    Odrv4 I__10980 (
            .O(N__59096),
            .I(\c0.n33957 ));
    InMux I__10979 (
            .O(N__59091),
            .I(N__59087));
    InMux I__10978 (
            .O(N__59090),
            .I(N__59084));
    LocalMux I__10977 (
            .O(N__59087),
            .I(N__59081));
    LocalMux I__10976 (
            .O(N__59084),
            .I(\c0.data_in_frame_21_0 ));
    Odrv4 I__10975 (
            .O(N__59081),
            .I(\c0.data_in_frame_21_0 ));
    InMux I__10974 (
            .O(N__59076),
            .I(N__59070));
    InMux I__10973 (
            .O(N__59075),
            .I(N__59070));
    LocalMux I__10972 (
            .O(N__59070),
            .I(\c0.data_in_frame_29_0 ));
    InMux I__10971 (
            .O(N__59067),
            .I(N__59064));
    LocalMux I__10970 (
            .O(N__59064),
            .I(\c0.n35181 ));
    CascadeMux I__10969 (
            .O(N__59061),
            .I(N__59058));
    InMux I__10968 (
            .O(N__59058),
            .I(N__59053));
    InMux I__10967 (
            .O(N__59057),
            .I(N__59048));
    InMux I__10966 (
            .O(N__59056),
            .I(N__59048));
    LocalMux I__10965 (
            .O(N__59053),
            .I(\c0.data_in_frame_22_1 ));
    LocalMux I__10964 (
            .O(N__59048),
            .I(\c0.data_in_frame_22_1 ));
    InMux I__10963 (
            .O(N__59043),
            .I(N__59039));
    InMux I__10962 (
            .O(N__59042),
            .I(N__59036));
    LocalMux I__10961 (
            .O(N__59039),
            .I(N__59033));
    LocalMux I__10960 (
            .O(N__59036),
            .I(N__59030));
    Odrv4 I__10959 (
            .O(N__59033),
            .I(\c0.n33598 ));
    Odrv4 I__10958 (
            .O(N__59030),
            .I(\c0.n33598 ));
    CascadeMux I__10957 (
            .O(N__59025),
            .I(\c0.n33374_cascade_ ));
    InMux I__10956 (
            .O(N__59022),
            .I(N__59018));
    CascadeMux I__10955 (
            .O(N__59021),
            .I(N__59015));
    LocalMux I__10954 (
            .O(N__59018),
            .I(N__59012));
    InMux I__10953 (
            .O(N__59015),
            .I(N__59009));
    Span4Mux_h I__10952 (
            .O(N__59012),
            .I(N__59006));
    LocalMux I__10951 (
            .O(N__59009),
            .I(\c0.data_in_frame_28_6 ));
    Odrv4 I__10950 (
            .O(N__59006),
            .I(\c0.data_in_frame_28_6 ));
    InMux I__10949 (
            .O(N__59001),
            .I(N__58998));
    LocalMux I__10948 (
            .O(N__58998),
            .I(N__58995));
    Odrv4 I__10947 (
            .O(N__58995),
            .I(\c0.n38_adj_4701 ));
    CascadeMux I__10946 (
            .O(N__58992),
            .I(N__58989));
    InMux I__10945 (
            .O(N__58989),
            .I(N__58986));
    LocalMux I__10944 (
            .O(N__58986),
            .I(\c0.n40_adj_4700 ));
    InMux I__10943 (
            .O(N__58983),
            .I(N__58980));
    LocalMux I__10942 (
            .O(N__58980),
            .I(\c0.n39_adj_4702 ));
    InMux I__10941 (
            .O(N__58977),
            .I(N__58974));
    LocalMux I__10940 (
            .O(N__58974),
            .I(\c0.n10_adj_4669 ));
    InMux I__10939 (
            .O(N__58971),
            .I(N__58968));
    LocalMux I__10938 (
            .O(N__58968),
            .I(N__58965));
    Odrv4 I__10937 (
            .O(N__58965),
            .I(\c0.n35307 ));
    CascadeMux I__10936 (
            .O(N__58962),
            .I(\c0.n16120_cascade_ ));
    InMux I__10935 (
            .O(N__58959),
            .I(N__58950));
    InMux I__10934 (
            .O(N__58958),
            .I(N__58950));
    InMux I__10933 (
            .O(N__58957),
            .I(N__58945));
    InMux I__10932 (
            .O(N__58956),
            .I(N__58945));
    InMux I__10931 (
            .O(N__58955),
            .I(N__58942));
    LocalMux I__10930 (
            .O(N__58950),
            .I(N__58939));
    LocalMux I__10929 (
            .O(N__58945),
            .I(N__58936));
    LocalMux I__10928 (
            .O(N__58942),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__10927 (
            .O(N__58939),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__10926 (
            .O(N__58936),
            .I(\c0.data_in_frame_19_5 ));
    InMux I__10925 (
            .O(N__58929),
            .I(N__58923));
    InMux I__10924 (
            .O(N__58928),
            .I(N__58923));
    LocalMux I__10923 (
            .O(N__58923),
            .I(N__58917));
    InMux I__10922 (
            .O(N__58922),
            .I(N__58914));
    InMux I__10921 (
            .O(N__58921),
            .I(N__58911));
    InMux I__10920 (
            .O(N__58920),
            .I(N__58908));
    Span4Mux_v I__10919 (
            .O(N__58917),
            .I(N__58905));
    LocalMux I__10918 (
            .O(N__58914),
            .I(N__58902));
    LocalMux I__10917 (
            .O(N__58911),
            .I(\c0.data_in_frame_23_3 ));
    LocalMux I__10916 (
            .O(N__58908),
            .I(\c0.data_in_frame_23_3 ));
    Odrv4 I__10915 (
            .O(N__58905),
            .I(\c0.data_in_frame_23_3 ));
    Odrv12 I__10914 (
            .O(N__58902),
            .I(\c0.data_in_frame_23_3 ));
    InMux I__10913 (
            .O(N__58893),
            .I(N__58890));
    LocalMux I__10912 (
            .O(N__58890),
            .I(\c0.n18784 ));
    CascadeMux I__10911 (
            .O(N__58887),
            .I(N__58884));
    InMux I__10910 (
            .O(N__58884),
            .I(N__58875));
    InMux I__10909 (
            .O(N__58883),
            .I(N__58875));
    InMux I__10908 (
            .O(N__58882),
            .I(N__58875));
    LocalMux I__10907 (
            .O(N__58875),
            .I(\c0.data_in_frame_20_4 ));
    InMux I__10906 (
            .O(N__58872),
            .I(N__58868));
    InMux I__10905 (
            .O(N__58871),
            .I(N__58865));
    LocalMux I__10904 (
            .O(N__58868),
            .I(N__58862));
    LocalMux I__10903 (
            .O(N__58865),
            .I(\c0.data_in_frame_22_5 ));
    Odrv4 I__10902 (
            .O(N__58862),
            .I(\c0.data_in_frame_22_5 ));
    InMux I__10901 (
            .O(N__58857),
            .I(N__58854));
    LocalMux I__10900 (
            .O(N__58854),
            .I(N__58851));
    Odrv4 I__10899 (
            .O(N__58851),
            .I(\c0.n6_adj_4675 ));
    InMux I__10898 (
            .O(N__58848),
            .I(N__58842));
    InMux I__10897 (
            .O(N__58847),
            .I(N__58842));
    LocalMux I__10896 (
            .O(N__58842),
            .I(\c0.data_in_frame_29_6 ));
    CascadeMux I__10895 (
            .O(N__58839),
            .I(\c0.n33506_cascade_ ));
    InMux I__10894 (
            .O(N__58836),
            .I(N__58833));
    LocalMux I__10893 (
            .O(N__58833),
            .I(N__58830));
    Span4Mux_h I__10892 (
            .O(N__58830),
            .I(N__58827));
    Odrv4 I__10891 (
            .O(N__58827),
            .I(\c0.n33889 ));
    CascadeMux I__10890 (
            .O(N__58824),
            .I(\c0.n12_adj_4710_cascade_ ));
    InMux I__10889 (
            .O(N__58821),
            .I(N__58817));
    InMux I__10888 (
            .O(N__58820),
            .I(N__58814));
    LocalMux I__10887 (
            .O(N__58817),
            .I(N__58811));
    LocalMux I__10886 (
            .O(N__58814),
            .I(\c0.n32346 ));
    Odrv4 I__10885 (
            .O(N__58811),
            .I(\c0.n32346 ));
    CascadeMux I__10884 (
            .O(N__58806),
            .I(\c0.n18784_cascade_ ));
    InMux I__10883 (
            .O(N__58803),
            .I(N__58800));
    LocalMux I__10882 (
            .O(N__58800),
            .I(\c0.n10_adj_4749 ));
    CascadeMux I__10881 (
            .O(N__58797),
            .I(N__58794));
    InMux I__10880 (
            .O(N__58794),
            .I(N__58790));
    CascadeMux I__10879 (
            .O(N__58793),
            .I(N__58786));
    LocalMux I__10878 (
            .O(N__58790),
            .I(N__58783));
    InMux I__10877 (
            .O(N__58789),
            .I(N__58779));
    InMux I__10876 (
            .O(N__58786),
            .I(N__58776));
    Span4Mux_v I__10875 (
            .O(N__58783),
            .I(N__58773));
    InMux I__10874 (
            .O(N__58782),
            .I(N__58770));
    LocalMux I__10873 (
            .O(N__58779),
            .I(N__58767));
    LocalMux I__10872 (
            .O(N__58776),
            .I(\c0.data_in_frame_23_6 ));
    Odrv4 I__10871 (
            .O(N__58773),
            .I(\c0.data_in_frame_23_6 ));
    LocalMux I__10870 (
            .O(N__58770),
            .I(\c0.data_in_frame_23_6 ));
    Odrv4 I__10869 (
            .O(N__58767),
            .I(\c0.data_in_frame_23_6 ));
    InMux I__10868 (
            .O(N__58758),
            .I(N__58755));
    LocalMux I__10867 (
            .O(N__58755),
            .I(\c0.n33726 ));
    InMux I__10866 (
            .O(N__58752),
            .I(N__58749));
    LocalMux I__10865 (
            .O(N__58749),
            .I(\c0.n33329 ));
    CascadeMux I__10864 (
            .O(N__58746),
            .I(\c0.n33726_cascade_ ));
    CascadeMux I__10863 (
            .O(N__58743),
            .I(N__58740));
    InMux I__10862 (
            .O(N__58740),
            .I(N__58737));
    LocalMux I__10861 (
            .O(N__58737),
            .I(\c0.n15_adj_4747 ));
    InMux I__10860 (
            .O(N__58734),
            .I(N__58730));
    InMux I__10859 (
            .O(N__58733),
            .I(N__58727));
    LocalMux I__10858 (
            .O(N__58730),
            .I(N__58721));
    LocalMux I__10857 (
            .O(N__58727),
            .I(N__58721));
    InMux I__10856 (
            .O(N__58726),
            .I(N__58718));
    Span4Mux_v I__10855 (
            .O(N__58721),
            .I(N__58713));
    LocalMux I__10854 (
            .O(N__58718),
            .I(N__58713));
    Odrv4 I__10853 (
            .O(N__58713),
            .I(\c0.n33532 ));
    CascadeMux I__10852 (
            .O(N__58710),
            .I(N__58706));
    CascadeMux I__10851 (
            .O(N__58709),
            .I(N__58703));
    InMux I__10850 (
            .O(N__58706),
            .I(N__58700));
    InMux I__10849 (
            .O(N__58703),
            .I(N__58697));
    LocalMux I__10848 (
            .O(N__58700),
            .I(N__58694));
    LocalMux I__10847 (
            .O(N__58697),
            .I(\c0.data_in_frame_6_0 ));
    Odrv4 I__10846 (
            .O(N__58694),
            .I(\c0.data_in_frame_6_0 ));
    InMux I__10845 (
            .O(N__58689),
            .I(N__58685));
    InMux I__10844 (
            .O(N__58688),
            .I(N__58682));
    LocalMux I__10843 (
            .O(N__58685),
            .I(N__58675));
    LocalMux I__10842 (
            .O(N__58682),
            .I(N__58672));
    InMux I__10841 (
            .O(N__58681),
            .I(N__58669));
    InMux I__10840 (
            .O(N__58680),
            .I(N__58666));
    CascadeMux I__10839 (
            .O(N__58679),
            .I(N__58663));
    InMux I__10838 (
            .O(N__58678),
            .I(N__58660));
    Span4Mux_v I__10837 (
            .O(N__58675),
            .I(N__58653));
    Span4Mux_v I__10836 (
            .O(N__58672),
            .I(N__58653));
    LocalMux I__10835 (
            .O(N__58669),
            .I(N__58653));
    LocalMux I__10834 (
            .O(N__58666),
            .I(N__58650));
    InMux I__10833 (
            .O(N__58663),
            .I(N__58647));
    LocalMux I__10832 (
            .O(N__58660),
            .I(N__58644));
    Span4Mux_h I__10831 (
            .O(N__58653),
            .I(N__58641));
    Span12Mux_v I__10830 (
            .O(N__58650),
            .I(N__58638));
    LocalMux I__10829 (
            .O(N__58647),
            .I(data_in_frame_1_2));
    Odrv12 I__10828 (
            .O(N__58644),
            .I(data_in_frame_1_2));
    Odrv4 I__10827 (
            .O(N__58641),
            .I(data_in_frame_1_2));
    Odrv12 I__10826 (
            .O(N__58638),
            .I(data_in_frame_1_2));
    InMux I__10825 (
            .O(N__58629),
            .I(N__58626));
    LocalMux I__10824 (
            .O(N__58626),
            .I(N__58623));
    Span4Mux_v I__10823 (
            .O(N__58623),
            .I(N__58620));
    Odrv4 I__10822 (
            .O(N__58620),
            .I(n36096));
    InMux I__10821 (
            .O(N__58617),
            .I(N__58614));
    LocalMux I__10820 (
            .O(N__58614),
            .I(N__58611));
    Sp12to4 I__10819 (
            .O(N__58611),
            .I(N__58608));
    Span12Mux_v I__10818 (
            .O(N__58608),
            .I(N__58605));
    Odrv12 I__10817 (
            .O(N__58605),
            .I(n10_adj_4820));
    CascadeMux I__10816 (
            .O(N__58602),
            .I(N__58598));
    InMux I__10815 (
            .O(N__58601),
            .I(N__58595));
    InMux I__10814 (
            .O(N__58598),
            .I(N__58592));
    LocalMux I__10813 (
            .O(N__58595),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__10812 (
            .O(N__58592),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__10811 (
            .O(N__58587),
            .I(\c0.rx.n30062 ));
    InMux I__10810 (
            .O(N__58584),
            .I(N__58580));
    InMux I__10809 (
            .O(N__58583),
            .I(N__58577));
    LocalMux I__10808 (
            .O(N__58580),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__10807 (
            .O(N__58577),
            .I(\c0.rx.r_Clock_Count_3 ));
    InMux I__10806 (
            .O(N__58572),
            .I(\c0.rx.n30063 ));
    InMux I__10805 (
            .O(N__58569),
            .I(\c0.rx.n30064 ));
    CascadeMux I__10804 (
            .O(N__58566),
            .I(N__58563));
    InMux I__10803 (
            .O(N__58563),
            .I(N__58560));
    LocalMux I__10802 (
            .O(N__58560),
            .I(N__58556));
    InMux I__10801 (
            .O(N__58559),
            .I(N__58551));
    Span4Mux_h I__10800 (
            .O(N__58556),
            .I(N__58548));
    InMux I__10799 (
            .O(N__58555),
            .I(N__58543));
    InMux I__10798 (
            .O(N__58554),
            .I(N__58543));
    LocalMux I__10797 (
            .O(N__58551),
            .I(\c0.rx.r_Clock_Count_5 ));
    Odrv4 I__10796 (
            .O(N__58548),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__10795 (
            .O(N__58543),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__10794 (
            .O(N__58536),
            .I(\c0.rx.n30065 ));
    InMux I__10793 (
            .O(N__58533),
            .I(N__58530));
    LocalMux I__10792 (
            .O(N__58530),
            .I(N__58526));
    InMux I__10791 (
            .O(N__58529),
            .I(N__58521));
    Span12Mux_v I__10790 (
            .O(N__58526),
            .I(N__58518));
    InMux I__10789 (
            .O(N__58525),
            .I(N__58513));
    InMux I__10788 (
            .O(N__58524),
            .I(N__58513));
    LocalMux I__10787 (
            .O(N__58521),
            .I(\c0.rx.r_Clock_Count_6 ));
    Odrv12 I__10786 (
            .O(N__58518),
            .I(\c0.rx.r_Clock_Count_6 ));
    LocalMux I__10785 (
            .O(N__58513),
            .I(\c0.rx.r_Clock_Count_6 ));
    InMux I__10784 (
            .O(N__58506),
            .I(\c0.rx.n30066 ));
    InMux I__10783 (
            .O(N__58503),
            .I(\c0.rx.n30067 ));
    InMux I__10782 (
            .O(N__58500),
            .I(N__58494));
    InMux I__10781 (
            .O(N__58499),
            .I(N__58487));
    InMux I__10780 (
            .O(N__58498),
            .I(N__58487));
    InMux I__10779 (
            .O(N__58497),
            .I(N__58487));
    LocalMux I__10778 (
            .O(N__58494),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__10777 (
            .O(N__58487),
            .I(\c0.rx.r_Clock_Count_7 ));
    CEMux I__10776 (
            .O(N__58482),
            .I(N__58479));
    LocalMux I__10775 (
            .O(N__58479),
            .I(N__58475));
    InMux I__10774 (
            .O(N__58478),
            .I(N__58472));
    Span4Mux_h I__10773 (
            .O(N__58475),
            .I(N__58469));
    LocalMux I__10772 (
            .O(N__58472),
            .I(N__58466));
    Odrv4 I__10771 (
            .O(N__58469),
            .I(n19327));
    Odrv4 I__10770 (
            .O(N__58466),
            .I(n19327));
    SRMux I__10769 (
            .O(N__58461),
            .I(N__58458));
    LocalMux I__10768 (
            .O(N__58458),
            .I(N__58454));
    InMux I__10767 (
            .O(N__58457),
            .I(N__58451));
    Span4Mux_v I__10766 (
            .O(N__58454),
            .I(N__58448));
    LocalMux I__10765 (
            .O(N__58451),
            .I(N__58445));
    Odrv4 I__10764 (
            .O(N__58448),
            .I(n19940));
    Odrv4 I__10763 (
            .O(N__58445),
            .I(n19940));
    CascadeMux I__10762 (
            .O(N__58440),
            .I(N__58433));
    CascadeMux I__10761 (
            .O(N__58439),
            .I(N__58423));
    CascadeMux I__10760 (
            .O(N__58438),
            .I(N__58420));
    InMux I__10759 (
            .O(N__58437),
            .I(N__58417));
    InMux I__10758 (
            .O(N__58436),
            .I(N__58407));
    InMux I__10757 (
            .O(N__58433),
            .I(N__58396));
    InMux I__10756 (
            .O(N__58432),
            .I(N__58396));
    InMux I__10755 (
            .O(N__58431),
            .I(N__58391));
    InMux I__10754 (
            .O(N__58430),
            .I(N__58391));
    InMux I__10753 (
            .O(N__58429),
            .I(N__58384));
    InMux I__10752 (
            .O(N__58428),
            .I(N__58384));
    InMux I__10751 (
            .O(N__58427),
            .I(N__58384));
    InMux I__10750 (
            .O(N__58426),
            .I(N__58374));
    InMux I__10749 (
            .O(N__58423),
            .I(N__58369));
    InMux I__10748 (
            .O(N__58420),
            .I(N__58369));
    LocalMux I__10747 (
            .O(N__58417),
            .I(N__58358));
    InMux I__10746 (
            .O(N__58416),
            .I(N__58349));
    InMux I__10745 (
            .O(N__58415),
            .I(N__58349));
    InMux I__10744 (
            .O(N__58414),
            .I(N__58349));
    InMux I__10743 (
            .O(N__58413),
            .I(N__58349));
    InMux I__10742 (
            .O(N__58412),
            .I(N__58344));
    InMux I__10741 (
            .O(N__58411),
            .I(N__58344));
    InMux I__10740 (
            .O(N__58410),
            .I(N__58341));
    LocalMux I__10739 (
            .O(N__58407),
            .I(N__58338));
    InMux I__10738 (
            .O(N__58406),
            .I(N__58335));
    InMux I__10737 (
            .O(N__58405),
            .I(N__58332));
    InMux I__10736 (
            .O(N__58404),
            .I(N__58323));
    InMux I__10735 (
            .O(N__58403),
            .I(N__58323));
    InMux I__10734 (
            .O(N__58402),
            .I(N__58323));
    InMux I__10733 (
            .O(N__58401),
            .I(N__58323));
    LocalMux I__10732 (
            .O(N__58396),
            .I(N__58313));
    LocalMux I__10731 (
            .O(N__58391),
            .I(N__58308));
    LocalMux I__10730 (
            .O(N__58384),
            .I(N__58308));
    InMux I__10729 (
            .O(N__58383),
            .I(N__58303));
    InMux I__10728 (
            .O(N__58382),
            .I(N__58303));
    InMux I__10727 (
            .O(N__58381),
            .I(N__58295));
    InMux I__10726 (
            .O(N__58380),
            .I(N__58288));
    InMux I__10725 (
            .O(N__58379),
            .I(N__58288));
    InMux I__10724 (
            .O(N__58378),
            .I(N__58288));
    InMux I__10723 (
            .O(N__58377),
            .I(N__58284));
    LocalMux I__10722 (
            .O(N__58374),
            .I(N__58279));
    LocalMux I__10721 (
            .O(N__58369),
            .I(N__58279));
    InMux I__10720 (
            .O(N__58368),
            .I(N__58276));
    InMux I__10719 (
            .O(N__58367),
            .I(N__58273));
    InMux I__10718 (
            .O(N__58366),
            .I(N__58270));
    CascadeMux I__10717 (
            .O(N__58365),
            .I(N__58267));
    InMux I__10716 (
            .O(N__58364),
            .I(N__58258));
    InMux I__10715 (
            .O(N__58363),
            .I(N__58258));
    InMux I__10714 (
            .O(N__58362),
            .I(N__58258));
    InMux I__10713 (
            .O(N__58361),
            .I(N__58258));
    Span4Mux_v I__10712 (
            .O(N__58358),
            .I(N__58249));
    LocalMux I__10711 (
            .O(N__58349),
            .I(N__58249));
    LocalMux I__10710 (
            .O(N__58344),
            .I(N__58249));
    LocalMux I__10709 (
            .O(N__58341),
            .I(N__58249));
    Span4Mux_v I__10708 (
            .O(N__58338),
            .I(N__58240));
    LocalMux I__10707 (
            .O(N__58335),
            .I(N__58240));
    LocalMux I__10706 (
            .O(N__58332),
            .I(N__58240));
    LocalMux I__10705 (
            .O(N__58323),
            .I(N__58240));
    InMux I__10704 (
            .O(N__58322),
            .I(N__58237));
    InMux I__10703 (
            .O(N__58321),
            .I(N__58234));
    InMux I__10702 (
            .O(N__58320),
            .I(N__58227));
    InMux I__10701 (
            .O(N__58319),
            .I(N__58227));
    InMux I__10700 (
            .O(N__58318),
            .I(N__58227));
    InMux I__10699 (
            .O(N__58317),
            .I(N__58222));
    InMux I__10698 (
            .O(N__58316),
            .I(N__58222));
    Span4Mux_v I__10697 (
            .O(N__58313),
            .I(N__58215));
    Span4Mux_v I__10696 (
            .O(N__58308),
            .I(N__58215));
    LocalMux I__10695 (
            .O(N__58303),
            .I(N__58215));
    InMux I__10694 (
            .O(N__58302),
            .I(N__58210));
    InMux I__10693 (
            .O(N__58301),
            .I(N__58210));
    InMux I__10692 (
            .O(N__58300),
            .I(N__58207));
    InMux I__10691 (
            .O(N__58299),
            .I(N__58199));
    InMux I__10690 (
            .O(N__58298),
            .I(N__58199));
    LocalMux I__10689 (
            .O(N__58295),
            .I(N__58196));
    LocalMux I__10688 (
            .O(N__58288),
            .I(N__58193));
    InMux I__10687 (
            .O(N__58287),
            .I(N__58190));
    LocalMux I__10686 (
            .O(N__58284),
            .I(N__58179));
    Span4Mux_h I__10685 (
            .O(N__58279),
            .I(N__58179));
    LocalMux I__10684 (
            .O(N__58276),
            .I(N__58179));
    LocalMux I__10683 (
            .O(N__58273),
            .I(N__58179));
    LocalMux I__10682 (
            .O(N__58270),
            .I(N__58179));
    InMux I__10681 (
            .O(N__58267),
            .I(N__58176));
    LocalMux I__10680 (
            .O(N__58258),
            .I(N__58169));
    Span4Mux_h I__10679 (
            .O(N__58249),
            .I(N__58169));
    Span4Mux_v I__10678 (
            .O(N__58240),
            .I(N__58169));
    LocalMux I__10677 (
            .O(N__58237),
            .I(N__58166));
    LocalMux I__10676 (
            .O(N__58234),
            .I(N__58157));
    LocalMux I__10675 (
            .O(N__58227),
            .I(N__58157));
    LocalMux I__10674 (
            .O(N__58222),
            .I(N__58157));
    Span4Mux_h I__10673 (
            .O(N__58215),
            .I(N__58157));
    LocalMux I__10672 (
            .O(N__58210),
            .I(N__58154));
    LocalMux I__10671 (
            .O(N__58207),
            .I(N__58151));
    InMux I__10670 (
            .O(N__58206),
            .I(N__58148));
    InMux I__10669 (
            .O(N__58205),
            .I(N__58143));
    InMux I__10668 (
            .O(N__58204),
            .I(N__58143));
    LocalMux I__10667 (
            .O(N__58199),
            .I(N__58140));
    Span4Mux_h I__10666 (
            .O(N__58196),
            .I(N__58135));
    Span4Mux_v I__10665 (
            .O(N__58193),
            .I(N__58135));
    LocalMux I__10664 (
            .O(N__58190),
            .I(N__58130));
    Span4Mux_v I__10663 (
            .O(N__58179),
            .I(N__58130));
    LocalMux I__10662 (
            .O(N__58176),
            .I(N__58125));
    Span4Mux_h I__10661 (
            .O(N__58169),
            .I(N__58125));
    Span4Mux_h I__10660 (
            .O(N__58166),
            .I(N__58120));
    Span4Mux_h I__10659 (
            .O(N__58157),
            .I(N__58120));
    Span12Mux_v I__10658 (
            .O(N__58154),
            .I(N__58115));
    Span12Mux_s10_h I__10657 (
            .O(N__58151),
            .I(N__58115));
    LocalMux I__10656 (
            .O(N__58148),
            .I(\c0.n33241 ));
    LocalMux I__10655 (
            .O(N__58143),
            .I(\c0.n33241 ));
    Odrv12 I__10654 (
            .O(N__58140),
            .I(\c0.n33241 ));
    Odrv4 I__10653 (
            .O(N__58135),
            .I(\c0.n33241 ));
    Odrv4 I__10652 (
            .O(N__58130),
            .I(\c0.n33241 ));
    Odrv4 I__10651 (
            .O(N__58125),
            .I(\c0.n33241 ));
    Odrv4 I__10650 (
            .O(N__58120),
            .I(\c0.n33241 ));
    Odrv12 I__10649 (
            .O(N__58115),
            .I(\c0.n33241 ));
    InMux I__10648 (
            .O(N__58098),
            .I(N__58094));
    InMux I__10647 (
            .O(N__58097),
            .I(N__58091));
    LocalMux I__10646 (
            .O(N__58094),
            .I(N__58088));
    LocalMux I__10645 (
            .O(N__58091),
            .I(N__58082));
    Span4Mux_v I__10644 (
            .O(N__58088),
            .I(N__58082));
    CascadeMux I__10643 (
            .O(N__58087),
            .I(N__58079));
    Span4Mux_h I__10642 (
            .O(N__58082),
            .I(N__58076));
    InMux I__10641 (
            .O(N__58079),
            .I(N__58073));
    Span4Mux_h I__10640 (
            .O(N__58076),
            .I(N__58070));
    LocalMux I__10639 (
            .O(N__58073),
            .I(\c0.data_in_frame_9_3 ));
    Odrv4 I__10638 (
            .O(N__58070),
            .I(\c0.data_in_frame_9_3 ));
    CascadeMux I__10637 (
            .O(N__58065),
            .I(\c0.rx.n19345_cascade_ ));
    CascadeMux I__10636 (
            .O(N__58062),
            .I(N__58058));
    CascadeMux I__10635 (
            .O(N__58061),
            .I(N__58055));
    InMux I__10634 (
            .O(N__58058),
            .I(N__58049));
    InMux I__10633 (
            .O(N__58055),
            .I(N__58049));
    InMux I__10632 (
            .O(N__58054),
            .I(N__58046));
    LocalMux I__10631 (
            .O(N__58049),
            .I(N__58043));
    LocalMux I__10630 (
            .O(N__58046),
            .I(\c0.rx.r_SM_Main_2_N_3681_2 ));
    Odrv4 I__10629 (
            .O(N__58043),
            .I(\c0.rx.r_SM_Main_2_N_3681_2 ));
    InMux I__10628 (
            .O(N__58038),
            .I(N__58034));
    InMux I__10627 (
            .O(N__58037),
            .I(N__58031));
    LocalMux I__10626 (
            .O(N__58034),
            .I(N__58028));
    LocalMux I__10625 (
            .O(N__58031),
            .I(N__58023));
    Span12Mux_v I__10624 (
            .O(N__58028),
            .I(N__58023));
    Odrv12 I__10623 (
            .O(N__58023),
            .I(\c0.rx.n17939 ));
    CascadeMux I__10622 (
            .O(N__58020),
            .I(N__58017));
    InMux I__10621 (
            .O(N__58017),
            .I(N__58013));
    InMux I__10620 (
            .O(N__58016),
            .I(N__58010));
    LocalMux I__10619 (
            .O(N__58013),
            .I(N__58006));
    LocalMux I__10618 (
            .O(N__58010),
            .I(N__58002));
    InMux I__10617 (
            .O(N__58009),
            .I(N__57999));
    Span12Mux_h I__10616 (
            .O(N__58006),
            .I(N__57996));
    InMux I__10615 (
            .O(N__58005),
            .I(N__57993));
    Span4Mux_h I__10614 (
            .O(N__58002),
            .I(N__57988));
    LocalMux I__10613 (
            .O(N__57999),
            .I(N__57988));
    Odrv12 I__10612 (
            .O(N__57996),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    LocalMux I__10611 (
            .O(N__57993),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    Odrv4 I__10610 (
            .O(N__57988),
            .I(\c0.FRAME_MATCHER_rx_data_ready_prev ));
    CascadeMux I__10609 (
            .O(N__57981),
            .I(N__57973));
    CascadeMux I__10608 (
            .O(N__57980),
            .I(N__57968));
    CascadeMux I__10607 (
            .O(N__57979),
            .I(N__57959));
    InMux I__10606 (
            .O(N__57978),
            .I(N__57949));
    InMux I__10605 (
            .O(N__57977),
            .I(N__57946));
    InMux I__10604 (
            .O(N__57976),
            .I(N__57942));
    InMux I__10603 (
            .O(N__57973),
            .I(N__57937));
    InMux I__10602 (
            .O(N__57972),
            .I(N__57937));
    InMux I__10601 (
            .O(N__57971),
            .I(N__57930));
    InMux I__10600 (
            .O(N__57968),
            .I(N__57930));
    InMux I__10599 (
            .O(N__57967),
            .I(N__57930));
    InMux I__10598 (
            .O(N__57966),
            .I(N__57923));
    InMux I__10597 (
            .O(N__57965),
            .I(N__57923));
    InMux I__10596 (
            .O(N__57964),
            .I(N__57923));
    InMux I__10595 (
            .O(N__57963),
            .I(N__57914));
    InMux I__10594 (
            .O(N__57962),
            .I(N__57914));
    InMux I__10593 (
            .O(N__57959),
            .I(N__57914));
    InMux I__10592 (
            .O(N__57958),
            .I(N__57914));
    CascadeMux I__10591 (
            .O(N__57957),
            .I(N__57904));
    CascadeMux I__10590 (
            .O(N__57956),
            .I(N__57901));
    InMux I__10589 (
            .O(N__57955),
            .I(N__57891));
    InMux I__10588 (
            .O(N__57954),
            .I(N__57891));
    InMux I__10587 (
            .O(N__57953),
            .I(N__57891));
    InMux I__10586 (
            .O(N__57952),
            .I(N__57891));
    LocalMux I__10585 (
            .O(N__57949),
            .I(N__57886));
    LocalMux I__10584 (
            .O(N__57946),
            .I(N__57886));
    InMux I__10583 (
            .O(N__57945),
            .I(N__57883));
    LocalMux I__10582 (
            .O(N__57942),
            .I(N__57880));
    LocalMux I__10581 (
            .O(N__57937),
            .I(N__57871));
    LocalMux I__10580 (
            .O(N__57930),
            .I(N__57871));
    LocalMux I__10579 (
            .O(N__57923),
            .I(N__57871));
    LocalMux I__10578 (
            .O(N__57914),
            .I(N__57871));
    InMux I__10577 (
            .O(N__57913),
            .I(N__57863));
    InMux I__10576 (
            .O(N__57912),
            .I(N__57863));
    InMux I__10575 (
            .O(N__57911),
            .I(N__57863));
    InMux I__10574 (
            .O(N__57910),
            .I(N__57858));
    InMux I__10573 (
            .O(N__57909),
            .I(N__57858));
    InMux I__10572 (
            .O(N__57908),
            .I(N__57853));
    InMux I__10571 (
            .O(N__57907),
            .I(N__57853));
    InMux I__10570 (
            .O(N__57904),
            .I(N__57848));
    InMux I__10569 (
            .O(N__57901),
            .I(N__57848));
    InMux I__10568 (
            .O(N__57900),
            .I(N__57845));
    LocalMux I__10567 (
            .O(N__57891),
            .I(N__57842));
    Span4Mux_v I__10566 (
            .O(N__57886),
            .I(N__57839));
    LocalMux I__10565 (
            .O(N__57883),
            .I(N__57835));
    Span4Mux_v I__10564 (
            .O(N__57880),
            .I(N__57830));
    Span4Mux_v I__10563 (
            .O(N__57871),
            .I(N__57830));
    InMux I__10562 (
            .O(N__57870),
            .I(N__57826));
    LocalMux I__10561 (
            .O(N__57863),
            .I(N__57823));
    LocalMux I__10560 (
            .O(N__57858),
            .I(N__57816));
    LocalMux I__10559 (
            .O(N__57853),
            .I(N__57816));
    LocalMux I__10558 (
            .O(N__57848),
            .I(N__57816));
    LocalMux I__10557 (
            .O(N__57845),
            .I(N__57809));
    Span4Mux_v I__10556 (
            .O(N__57842),
            .I(N__57809));
    Span4Mux_h I__10555 (
            .O(N__57839),
            .I(N__57809));
    InMux I__10554 (
            .O(N__57838),
            .I(N__57806));
    Span4Mux_v I__10553 (
            .O(N__57835),
            .I(N__57801));
    Span4Mux_h I__10552 (
            .O(N__57830),
            .I(N__57801));
    CascadeMux I__10551 (
            .O(N__57829),
            .I(N__57798));
    LocalMux I__10550 (
            .O(N__57826),
            .I(N__57794));
    Span4Mux_h I__10549 (
            .O(N__57823),
            .I(N__57789));
    Span4Mux_v I__10548 (
            .O(N__57816),
            .I(N__57789));
    Span4Mux_h I__10547 (
            .O(N__57809),
            .I(N__57784));
    LocalMux I__10546 (
            .O(N__57806),
            .I(N__57779));
    Span4Mux_h I__10545 (
            .O(N__57801),
            .I(N__57779));
    InMux I__10544 (
            .O(N__57798),
            .I(N__57776));
    InMux I__10543 (
            .O(N__57797),
            .I(N__57773));
    Span4Mux_v I__10542 (
            .O(N__57794),
            .I(N__57768));
    Span4Mux_h I__10541 (
            .O(N__57789),
            .I(N__57765));
    InMux I__10540 (
            .O(N__57788),
            .I(N__57762));
    InMux I__10539 (
            .O(N__57787),
            .I(N__57759));
    Span4Mux_h I__10538 (
            .O(N__57784),
            .I(N__57756));
    Span4Mux_v I__10537 (
            .O(N__57779),
            .I(N__57751));
    LocalMux I__10536 (
            .O(N__57776),
            .I(N__57751));
    LocalMux I__10535 (
            .O(N__57773),
            .I(N__57748));
    InMux I__10534 (
            .O(N__57772),
            .I(N__57743));
    InMux I__10533 (
            .O(N__57771),
            .I(N__57743));
    Span4Mux_h I__10532 (
            .O(N__57768),
            .I(N__57736));
    Span4Mux_h I__10531 (
            .O(N__57765),
            .I(N__57736));
    LocalMux I__10530 (
            .O(N__57762),
            .I(N__57736));
    LocalMux I__10529 (
            .O(N__57759),
            .I(rx_data_ready));
    Odrv4 I__10528 (
            .O(N__57756),
            .I(rx_data_ready));
    Odrv4 I__10527 (
            .O(N__57751),
            .I(rx_data_ready));
    Odrv4 I__10526 (
            .O(N__57748),
            .I(rx_data_ready));
    LocalMux I__10525 (
            .O(N__57743),
            .I(rx_data_ready));
    Odrv4 I__10524 (
            .O(N__57736),
            .I(rx_data_ready));
    CascadeMux I__10523 (
            .O(N__57723),
            .I(N__57719));
    InMux I__10522 (
            .O(N__57722),
            .I(N__57715));
    InMux I__10521 (
            .O(N__57719),
            .I(N__57710));
    InMux I__10520 (
            .O(N__57718),
            .I(N__57710));
    LocalMux I__10519 (
            .O(N__57715),
            .I(r_Clock_Count_0));
    LocalMux I__10518 (
            .O(N__57710),
            .I(r_Clock_Count_0));
    InMux I__10517 (
            .O(N__57705),
            .I(N__57702));
    LocalMux I__10516 (
            .O(N__57702),
            .I(n226));
    InMux I__10515 (
            .O(N__57699),
            .I(bfn_16_21_0_));
    InMux I__10514 (
            .O(N__57696),
            .I(N__57692));
    InMux I__10513 (
            .O(N__57695),
            .I(N__57689));
    LocalMux I__10512 (
            .O(N__57692),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__10511 (
            .O(N__57689),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__10510 (
            .O(N__57684),
            .I(\c0.rx.n30061 ));
    InMux I__10509 (
            .O(N__57681),
            .I(N__57678));
    LocalMux I__10508 (
            .O(N__57678),
            .I(\c0.n7_adj_4499 ));
    InMux I__10507 (
            .O(N__57675),
            .I(N__57672));
    LocalMux I__10506 (
            .O(N__57672),
            .I(n35818));
    InMux I__10505 (
            .O(N__57669),
            .I(N__57664));
    InMux I__10504 (
            .O(N__57668),
            .I(N__57661));
    InMux I__10503 (
            .O(N__57667),
            .I(N__57658));
    LocalMux I__10502 (
            .O(N__57664),
            .I(N__57653));
    LocalMux I__10501 (
            .O(N__57661),
            .I(N__57653));
    LocalMux I__10500 (
            .O(N__57658),
            .I(\c0.data_in_frame_4_1 ));
    Odrv12 I__10499 (
            .O(N__57653),
            .I(\c0.data_in_frame_4_1 ));
    CascadeMux I__10498 (
            .O(N__57648),
            .I(N__57645));
    InMux I__10497 (
            .O(N__57645),
            .I(N__57642));
    LocalMux I__10496 (
            .O(N__57642),
            .I(N__57636));
    InMux I__10495 (
            .O(N__57641),
            .I(N__57633));
    InMux I__10494 (
            .O(N__57640),
            .I(N__57630));
    CascadeMux I__10493 (
            .O(N__57639),
            .I(N__57627));
    Span4Mux_v I__10492 (
            .O(N__57636),
            .I(N__57624));
    LocalMux I__10491 (
            .O(N__57633),
            .I(N__57621));
    LocalMux I__10490 (
            .O(N__57630),
            .I(N__57618));
    InMux I__10489 (
            .O(N__57627),
            .I(N__57615));
    Span4Mux_h I__10488 (
            .O(N__57624),
            .I(N__57612));
    Span4Mux_v I__10487 (
            .O(N__57621),
            .I(N__57607));
    Span4Mux_v I__10486 (
            .O(N__57618),
            .I(N__57607));
    LocalMux I__10485 (
            .O(N__57615),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__10484 (
            .O(N__57612),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__10483 (
            .O(N__57607),
            .I(\c0.data_in_frame_2_1 ));
    InMux I__10482 (
            .O(N__57600),
            .I(N__57596));
    InMux I__10481 (
            .O(N__57599),
            .I(N__57593));
    LocalMux I__10480 (
            .O(N__57596),
            .I(data_out_frame_13_6));
    LocalMux I__10479 (
            .O(N__57593),
            .I(data_out_frame_13_6));
    InMux I__10478 (
            .O(N__57588),
            .I(N__57584));
    InMux I__10477 (
            .O(N__57587),
            .I(N__57581));
    LocalMux I__10476 (
            .O(N__57584),
            .I(data_out_frame_8_0));
    LocalMux I__10475 (
            .O(N__57581),
            .I(data_out_frame_8_0));
    InMux I__10474 (
            .O(N__57576),
            .I(N__57573));
    LocalMux I__10473 (
            .O(N__57573),
            .I(N__57570));
    Span4Mux_h I__10472 (
            .O(N__57570),
            .I(N__57567));
    Span4Mux_h I__10471 (
            .O(N__57567),
            .I(N__57563));
    InMux I__10470 (
            .O(N__57566),
            .I(N__57560));
    Span4Mux_v I__10469 (
            .O(N__57563),
            .I(N__57557));
    LocalMux I__10468 (
            .O(N__57560),
            .I(data_out_frame_9_7));
    Odrv4 I__10467 (
            .O(N__57557),
            .I(data_out_frame_9_7));
    CascadeMux I__10466 (
            .O(N__57552),
            .I(\c0.n36194_cascade_ ));
    InMux I__10465 (
            .O(N__57549),
            .I(N__57546));
    LocalMux I__10464 (
            .O(N__57546),
            .I(\c0.n11_adj_4655 ));
    InMux I__10463 (
            .O(N__57543),
            .I(N__57540));
    LocalMux I__10462 (
            .O(N__57540),
            .I(n36094));
    InMux I__10461 (
            .O(N__57537),
            .I(N__57534));
    LocalMux I__10460 (
            .O(N__57534),
            .I(N__57531));
    Odrv4 I__10459 (
            .O(N__57531),
            .I(\c0.n5 ));
    InMux I__10458 (
            .O(N__57528),
            .I(N__57524));
    InMux I__10457 (
            .O(N__57527),
            .I(N__57521));
    LocalMux I__10456 (
            .O(N__57524),
            .I(data_out_frame_7_3));
    LocalMux I__10455 (
            .O(N__57521),
            .I(data_out_frame_7_3));
    InMux I__10454 (
            .O(N__57516),
            .I(N__57510));
    InMux I__10453 (
            .O(N__57515),
            .I(N__57510));
    LocalMux I__10452 (
            .O(N__57510),
            .I(data_out_frame_6_3));
    InMux I__10451 (
            .O(N__57507),
            .I(N__57503));
    InMux I__10450 (
            .O(N__57506),
            .I(N__57500));
    LocalMux I__10449 (
            .O(N__57503),
            .I(data_out_frame_12_6));
    LocalMux I__10448 (
            .O(N__57500),
            .I(data_out_frame_12_6));
    CascadeMux I__10447 (
            .O(N__57495),
            .I(\c0.n6_adj_4647_cascade_ ));
    InMux I__10446 (
            .O(N__57492),
            .I(N__57483));
    InMux I__10445 (
            .O(N__57491),
            .I(N__57483));
    InMux I__10444 (
            .O(N__57490),
            .I(N__57483));
    LocalMux I__10443 (
            .O(N__57483),
            .I(N__57480));
    Odrv12 I__10442 (
            .O(N__57480),
            .I(\c0.n28313 ));
    InMux I__10441 (
            .O(N__57477),
            .I(N__57473));
    InMux I__10440 (
            .O(N__57476),
            .I(N__57470));
    LocalMux I__10439 (
            .O(N__57473),
            .I(N__57465));
    LocalMux I__10438 (
            .O(N__57470),
            .I(N__57465));
    Odrv4 I__10437 (
            .O(N__57465),
            .I(data_out_frame_9_2));
    CascadeMux I__10436 (
            .O(N__57462),
            .I(N__57459));
    InMux I__10435 (
            .O(N__57459),
            .I(N__57453));
    InMux I__10434 (
            .O(N__57458),
            .I(N__57453));
    LocalMux I__10433 (
            .O(N__57453),
            .I(data_out_frame_8_2));
    InMux I__10432 (
            .O(N__57450),
            .I(N__57447));
    LocalMux I__10431 (
            .O(N__57447),
            .I(\c0.n36206 ));
    InMux I__10430 (
            .O(N__57444),
            .I(N__57441));
    LocalMux I__10429 (
            .O(N__57441),
            .I(n10));
    InMux I__10428 (
            .O(N__57438),
            .I(N__57435));
    LocalMux I__10427 (
            .O(N__57435),
            .I(N__57432));
    Odrv4 I__10426 (
            .O(N__57432),
            .I(n10_adj_4806));
    InMux I__10425 (
            .O(N__57429),
            .I(N__57426));
    LocalMux I__10424 (
            .O(N__57426),
            .I(N__57423));
    Odrv4 I__10423 (
            .O(N__57423),
            .I(\c0.n35963 ));
    InMux I__10422 (
            .O(N__57420),
            .I(N__57416));
    InMux I__10421 (
            .O(N__57419),
            .I(N__57413));
    LocalMux I__10420 (
            .O(N__57416),
            .I(data_out_frame_11_2));
    LocalMux I__10419 (
            .O(N__57413),
            .I(data_out_frame_11_2));
    InMux I__10418 (
            .O(N__57408),
            .I(N__57402));
    InMux I__10417 (
            .O(N__57407),
            .I(N__57402));
    LocalMux I__10416 (
            .O(N__57402),
            .I(data_out_frame_10_2));
    InMux I__10415 (
            .O(N__57399),
            .I(N__57396));
    LocalMux I__10414 (
            .O(N__57396),
            .I(\c0.n36203 ));
    CascadeMux I__10413 (
            .O(N__57393),
            .I(N__57389));
    CascadeMux I__10412 (
            .O(N__57392),
            .I(N__57385));
    InMux I__10411 (
            .O(N__57389),
            .I(N__57382));
    InMux I__10410 (
            .O(N__57388),
            .I(N__57379));
    InMux I__10409 (
            .O(N__57385),
            .I(N__57376));
    LocalMux I__10408 (
            .O(N__57382),
            .I(N__57373));
    LocalMux I__10407 (
            .O(N__57379),
            .I(\quad_counter0.n3516 ));
    LocalMux I__10406 (
            .O(N__57376),
            .I(\quad_counter0.n3516 ));
    Odrv4 I__10405 (
            .O(N__57373),
            .I(\quad_counter0.n3516 ));
    InMux I__10404 (
            .O(N__57366),
            .I(\quad_counter0.n30456 ));
    InMux I__10403 (
            .O(N__57363),
            .I(N__57360));
    LocalMux I__10402 (
            .O(N__57360),
            .I(\quad_counter0.n12904 ));
    InMux I__10401 (
            .O(N__57357),
            .I(N__57352));
    InMux I__10400 (
            .O(N__57356),
            .I(N__57347));
    InMux I__10399 (
            .O(N__57355),
            .I(N__57347));
    LocalMux I__10398 (
            .O(N__57352),
            .I(N__57344));
    LocalMux I__10397 (
            .O(N__57347),
            .I(\quad_counter0.n3515 ));
    Odrv4 I__10396 (
            .O(N__57344),
            .I(\quad_counter0.n3515 ));
    InMux I__10395 (
            .O(N__57339),
            .I(N__57336));
    LocalMux I__10394 (
            .O(N__57336),
            .I(\quad_counter0.n8_adj_4375 ));
    InMux I__10393 (
            .O(N__57333),
            .I(\quad_counter0.n30457 ));
    InMux I__10392 (
            .O(N__57330),
            .I(N__57327));
    LocalMux I__10391 (
            .O(N__57327),
            .I(\quad_counter0.n12901 ));
    CascadeMux I__10390 (
            .O(N__57324),
            .I(N__57321));
    InMux I__10389 (
            .O(N__57321),
            .I(N__57318));
    LocalMux I__10388 (
            .O(N__57318),
            .I(N__57313));
    InMux I__10387 (
            .O(N__57317),
            .I(N__57310));
    InMux I__10386 (
            .O(N__57316),
            .I(N__57307));
    Odrv4 I__10385 (
            .O(N__57313),
            .I(\quad_counter0.n3514 ));
    LocalMux I__10384 (
            .O(N__57310),
            .I(\quad_counter0.n3514 ));
    LocalMux I__10383 (
            .O(N__57307),
            .I(\quad_counter0.n3514 ));
    InMux I__10382 (
            .O(N__57300),
            .I(\quad_counter0.n30458 ));
    InMux I__10381 (
            .O(N__57297),
            .I(N__57294));
    LocalMux I__10380 (
            .O(N__57294),
            .I(\quad_counter0.n10_adj_4347 ));
    InMux I__10379 (
            .O(N__57291),
            .I(N__57288));
    LocalMux I__10378 (
            .O(N__57288),
            .I(\quad_counter0.n11 ));
    CascadeMux I__10377 (
            .O(N__57285),
            .I(\quad_counter0.n28339_cascade_ ));
    InMux I__10376 (
            .O(N__57282),
            .I(N__57279));
    LocalMux I__10375 (
            .O(N__57279),
            .I(\quad_counter0.n10_adj_4400 ));
    CascadeMux I__10374 (
            .O(N__57276),
            .I(\quad_counter0.n10_adj_4399_cascade_ ));
    CascadeMux I__10373 (
            .O(N__57273),
            .I(N__57270));
    InMux I__10372 (
            .O(N__57270),
            .I(N__57267));
    LocalMux I__10371 (
            .O(N__57267),
            .I(\quad_counter0.n16_adj_4401 ));
    InMux I__10370 (
            .O(N__57264),
            .I(N__57261));
    LocalMux I__10369 (
            .O(N__57261),
            .I(N__57258));
    Span4Mux_h I__10368 (
            .O(N__57258),
            .I(N__57255));
    Odrv4 I__10367 (
            .O(N__57255),
            .I(\quad_counter0.n35976 ));
    CascadeMux I__10366 (
            .O(N__57252),
            .I(\quad_counter0.n35977_cascade_ ));
    InMux I__10365 (
            .O(N__57249),
            .I(N__57246));
    LocalMux I__10364 (
            .O(N__57246),
            .I(N__57243));
    Span4Mux_h I__10363 (
            .O(N__57243),
            .I(N__57240));
    Odrv4 I__10362 (
            .O(N__57240),
            .I(\quad_counter0.n33_adj_4346 ));
    InMux I__10361 (
            .O(N__57237),
            .I(N__57234));
    LocalMux I__10360 (
            .O(N__57234),
            .I(\quad_counter0.n34205 ));
    InMux I__10359 (
            .O(N__57231),
            .I(N__57228));
    LocalMux I__10358 (
            .O(N__57228),
            .I(\quad_counter0.n3508 ));
    InMux I__10357 (
            .O(N__57225),
            .I(N__57222));
    LocalMux I__10356 (
            .O(N__57222),
            .I(\quad_counter0.n3501 ));
    CascadeMux I__10355 (
            .O(N__57219),
            .I(N__57216));
    InMux I__10354 (
            .O(N__57216),
            .I(N__57213));
    LocalMux I__10353 (
            .O(N__57213),
            .I(\quad_counter0.n3504 ));
    InMux I__10352 (
            .O(N__57210),
            .I(N__57207));
    LocalMux I__10351 (
            .O(N__57207),
            .I(\quad_counter0.n3499 ));
    InMux I__10350 (
            .O(N__57204),
            .I(N__57201));
    LocalMux I__10349 (
            .O(N__57201),
            .I(\quad_counter0.n3502 ));
    InMux I__10348 (
            .O(N__57198),
            .I(N__57195));
    LocalMux I__10347 (
            .O(N__57195),
            .I(\quad_counter0.n3498 ));
    CascadeMux I__10346 (
            .O(N__57192),
            .I(\quad_counter0.n31_cascade_ ));
    InMux I__10345 (
            .O(N__57189),
            .I(N__57186));
    LocalMux I__10344 (
            .O(N__57186),
            .I(\quad_counter0.n28_adj_4342 ));
    InMux I__10343 (
            .O(N__57183),
            .I(N__57180));
    LocalMux I__10342 (
            .O(N__57180),
            .I(\quad_counter0.n34 ));
    CascadeMux I__10341 (
            .O(N__57177),
            .I(N__57174));
    InMux I__10340 (
            .O(N__57174),
            .I(N__57171));
    LocalMux I__10339 (
            .O(N__57171),
            .I(\quad_counter0.n35978 ));
    InMux I__10338 (
            .O(N__57168),
            .I(bfn_16_12_0_));
    CascadeMux I__10337 (
            .O(N__57165),
            .I(N__57162));
    InMux I__10336 (
            .O(N__57162),
            .I(N__57158));
    CascadeMux I__10335 (
            .O(N__57161),
            .I(N__57155));
    LocalMux I__10334 (
            .O(N__57158),
            .I(N__57151));
    InMux I__10333 (
            .O(N__57155),
            .I(N__57146));
    InMux I__10332 (
            .O(N__57154),
            .I(N__57146));
    Span4Mux_v I__10331 (
            .O(N__57151),
            .I(N__57143));
    LocalMux I__10330 (
            .O(N__57146),
            .I(\quad_counter0.n3519 ));
    Odrv4 I__10329 (
            .O(N__57143),
            .I(\quad_counter0.n3519 ));
    InMux I__10328 (
            .O(N__57138),
            .I(\quad_counter0.n30453 ));
    CascadeMux I__10327 (
            .O(N__57135),
            .I(N__57132));
    InMux I__10326 (
            .O(N__57132),
            .I(N__57129));
    LocalMux I__10325 (
            .O(N__57129),
            .I(N__57124));
    InMux I__10324 (
            .O(N__57128),
            .I(N__57121));
    InMux I__10323 (
            .O(N__57127),
            .I(N__57118));
    Span4Mux_v I__10322 (
            .O(N__57124),
            .I(N__57115));
    LocalMux I__10321 (
            .O(N__57121),
            .I(\quad_counter0.n3518 ));
    LocalMux I__10320 (
            .O(N__57118),
            .I(\quad_counter0.n3518 ));
    Odrv4 I__10319 (
            .O(N__57115),
            .I(\quad_counter0.n3518 ));
    InMux I__10318 (
            .O(N__57108),
            .I(\quad_counter0.n30454 ));
    InMux I__10317 (
            .O(N__57105),
            .I(N__57102));
    LocalMux I__10316 (
            .O(N__57102),
            .I(\quad_counter0.n12903 ));
    CascadeMux I__10315 (
            .O(N__57099),
            .I(N__57096));
    InMux I__10314 (
            .O(N__57096),
            .I(N__57091));
    InMux I__10313 (
            .O(N__57095),
            .I(N__57088));
    InMux I__10312 (
            .O(N__57094),
            .I(N__57085));
    LocalMux I__10311 (
            .O(N__57091),
            .I(N__57082));
    LocalMux I__10310 (
            .O(N__57088),
            .I(\quad_counter0.n3517 ));
    LocalMux I__10309 (
            .O(N__57085),
            .I(\quad_counter0.n3517 ));
    Odrv4 I__10308 (
            .O(N__57082),
            .I(\quad_counter0.n3517 ));
    InMux I__10307 (
            .O(N__57075),
            .I(N__57072));
    LocalMux I__10306 (
            .O(N__57072),
            .I(\quad_counter0.n9 ));
    InMux I__10305 (
            .O(N__57069),
            .I(\quad_counter0.n30455 ));
    InMux I__10304 (
            .O(N__57066),
            .I(N__57062));
    InMux I__10303 (
            .O(N__57065),
            .I(N__57059));
    LocalMux I__10302 (
            .O(N__57062),
            .I(N__57054));
    LocalMux I__10301 (
            .O(N__57059),
            .I(N__57054));
    Span4Mux_h I__10300 (
            .O(N__57054),
            .I(N__57050));
    InMux I__10299 (
            .O(N__57053),
            .I(N__57047));
    Odrv4 I__10298 (
            .O(N__57050),
            .I(\quad_counter0.n2111 ));
    LocalMux I__10297 (
            .O(N__57047),
            .I(\quad_counter0.n2111 ));
    InMux I__10296 (
            .O(N__57042),
            .I(\quad_counter0.n30238 ));
    CascadeMux I__10295 (
            .O(N__57039),
            .I(N__57033));
    CascadeMux I__10294 (
            .O(N__57038),
            .I(N__57030));
    CascadeMux I__10293 (
            .O(N__57037),
            .I(N__57027));
    CascadeMux I__10292 (
            .O(N__57036),
            .I(N__57024));
    InMux I__10291 (
            .O(N__57033),
            .I(N__57020));
    InMux I__10290 (
            .O(N__57030),
            .I(N__57015));
    InMux I__10289 (
            .O(N__57027),
            .I(N__57015));
    InMux I__10288 (
            .O(N__57024),
            .I(N__57010));
    InMux I__10287 (
            .O(N__57023),
            .I(N__57010));
    LocalMux I__10286 (
            .O(N__57020),
            .I(\quad_counter0.n2144 ));
    LocalMux I__10285 (
            .O(N__57015),
            .I(\quad_counter0.n2144 ));
    LocalMux I__10284 (
            .O(N__57010),
            .I(\quad_counter0.n2144 ));
    CascadeMux I__10283 (
            .O(N__57003),
            .I(N__56995));
    CascadeMux I__10282 (
            .O(N__57002),
            .I(N__56992));
    CascadeMux I__10281 (
            .O(N__57001),
            .I(N__56989));
    CascadeMux I__10280 (
            .O(N__57000),
            .I(N__56986));
    CascadeMux I__10279 (
            .O(N__56999),
            .I(N__56983));
    CascadeMux I__10278 (
            .O(N__56998),
            .I(N__56980));
    InMux I__10277 (
            .O(N__56995),
            .I(N__56975));
    InMux I__10276 (
            .O(N__56992),
            .I(N__56975));
    InMux I__10275 (
            .O(N__56989),
            .I(N__56966));
    InMux I__10274 (
            .O(N__56986),
            .I(N__56966));
    InMux I__10273 (
            .O(N__56983),
            .I(N__56966));
    InMux I__10272 (
            .O(N__56980),
            .I(N__56966));
    LocalMux I__10271 (
            .O(N__56975),
            .I(\quad_counter0.n36157 ));
    LocalMux I__10270 (
            .O(N__56966),
            .I(\quad_counter0.n36157 ));
    CascadeMux I__10269 (
            .O(N__56961),
            .I(\quad_counter0.n10_adj_4389_cascade_ ));
    InMux I__10268 (
            .O(N__56958),
            .I(N__56955));
    LocalMux I__10267 (
            .O(N__56955),
            .I(N__56952));
    Odrv4 I__10266 (
            .O(N__56952),
            .I(\quad_counter0.n14_adj_4418 ));
    CascadeMux I__10265 (
            .O(N__56949),
            .I(\quad_counter0.n15_cascade_ ));
    InMux I__10264 (
            .O(N__56946),
            .I(N__56943));
    LocalMux I__10263 (
            .O(N__56943),
            .I(N__56940));
    Odrv4 I__10262 (
            .O(N__56940),
            .I(\quad_counter0.n3512 ));
    InMux I__10261 (
            .O(N__56937),
            .I(N__56934));
    LocalMux I__10260 (
            .O(N__56934),
            .I(N__56931));
    Odrv4 I__10259 (
            .O(N__56931),
            .I(\quad_counter0.n3513 ));
    CascadeMux I__10258 (
            .O(N__56928),
            .I(N__56925));
    InMux I__10257 (
            .O(N__56925),
            .I(N__56922));
    LocalMux I__10256 (
            .O(N__56922),
            .I(\quad_counter0.n3507 ));
    InMux I__10255 (
            .O(N__56919),
            .I(N__56916));
    LocalMux I__10254 (
            .O(N__56916),
            .I(\quad_counter0.n3500 ));
    InMux I__10253 (
            .O(N__56913),
            .I(N__56909));
    InMux I__10252 (
            .O(N__56912),
            .I(N__56906));
    LocalMux I__10251 (
            .O(N__56909),
            .I(N__56903));
    LocalMux I__10250 (
            .O(N__56906),
            .I(N__56900));
    Odrv12 I__10249 (
            .O(N__56903),
            .I(\quad_counter0.n2119 ));
    Odrv4 I__10248 (
            .O(N__56900),
            .I(\quad_counter0.n2119 ));
    InMux I__10247 (
            .O(N__56895),
            .I(\quad_counter0.n30230 ));
    InMux I__10246 (
            .O(N__56892),
            .I(N__56888));
    InMux I__10245 (
            .O(N__56891),
            .I(N__56885));
    LocalMux I__10244 (
            .O(N__56888),
            .I(N__56880));
    LocalMux I__10243 (
            .O(N__56885),
            .I(N__56880));
    Span4Mux_h I__10242 (
            .O(N__56880),
            .I(N__56876));
    InMux I__10241 (
            .O(N__56879),
            .I(N__56873));
    Odrv4 I__10240 (
            .O(N__56876),
            .I(\quad_counter0.n2118 ));
    LocalMux I__10239 (
            .O(N__56873),
            .I(\quad_counter0.n2118 ));
    InMux I__10238 (
            .O(N__56868),
            .I(\quad_counter0.n30231 ));
    CascadeMux I__10237 (
            .O(N__56865),
            .I(N__56860));
    InMux I__10236 (
            .O(N__56864),
            .I(N__56857));
    InMux I__10235 (
            .O(N__56863),
            .I(N__56854));
    InMux I__10234 (
            .O(N__56860),
            .I(N__56851));
    LocalMux I__10233 (
            .O(N__56857),
            .I(\quad_counter0.n2117 ));
    LocalMux I__10232 (
            .O(N__56854),
            .I(\quad_counter0.n2117 ));
    LocalMux I__10231 (
            .O(N__56851),
            .I(\quad_counter0.n2117 ));
    InMux I__10230 (
            .O(N__56844),
            .I(\quad_counter0.n30232 ));
    InMux I__10229 (
            .O(N__56841),
            .I(N__56836));
    InMux I__10228 (
            .O(N__56840),
            .I(N__56833));
    InMux I__10227 (
            .O(N__56839),
            .I(N__56830));
    LocalMux I__10226 (
            .O(N__56836),
            .I(\quad_counter0.n2116 ));
    LocalMux I__10225 (
            .O(N__56833),
            .I(\quad_counter0.n2116 ));
    LocalMux I__10224 (
            .O(N__56830),
            .I(\quad_counter0.n2116 ));
    InMux I__10223 (
            .O(N__56823),
            .I(\quad_counter0.n30233 ));
    InMux I__10222 (
            .O(N__56820),
            .I(N__56815));
    InMux I__10221 (
            .O(N__56819),
            .I(N__56812));
    InMux I__10220 (
            .O(N__56818),
            .I(N__56809));
    LocalMux I__10219 (
            .O(N__56815),
            .I(\quad_counter0.n2115 ));
    LocalMux I__10218 (
            .O(N__56812),
            .I(\quad_counter0.n2115 ));
    LocalMux I__10217 (
            .O(N__56809),
            .I(\quad_counter0.n2115 ));
    InMux I__10216 (
            .O(N__56802),
            .I(\quad_counter0.n30234 ));
    InMux I__10215 (
            .O(N__56799),
            .I(N__56794));
    InMux I__10214 (
            .O(N__56798),
            .I(N__56791));
    InMux I__10213 (
            .O(N__56797),
            .I(N__56788));
    LocalMux I__10212 (
            .O(N__56794),
            .I(\quad_counter0.n2114 ));
    LocalMux I__10211 (
            .O(N__56791),
            .I(\quad_counter0.n2114 ));
    LocalMux I__10210 (
            .O(N__56788),
            .I(\quad_counter0.n2114 ));
    InMux I__10209 (
            .O(N__56781),
            .I(\quad_counter0.n30235 ));
    InMux I__10208 (
            .O(N__56778),
            .I(N__56774));
    InMux I__10207 (
            .O(N__56777),
            .I(N__56771));
    LocalMux I__10206 (
            .O(N__56774),
            .I(N__56765));
    LocalMux I__10205 (
            .O(N__56771),
            .I(N__56765));
    InMux I__10204 (
            .O(N__56770),
            .I(N__56762));
    Odrv4 I__10203 (
            .O(N__56765),
            .I(\quad_counter0.n2113 ));
    LocalMux I__10202 (
            .O(N__56762),
            .I(\quad_counter0.n2113 ));
    InMux I__10201 (
            .O(N__56757),
            .I(\quad_counter0.n30236 ));
    InMux I__10200 (
            .O(N__56754),
            .I(N__56750));
    InMux I__10199 (
            .O(N__56753),
            .I(N__56747));
    LocalMux I__10198 (
            .O(N__56750),
            .I(N__56741));
    LocalMux I__10197 (
            .O(N__56747),
            .I(N__56741));
    InMux I__10196 (
            .O(N__56746),
            .I(N__56738));
    Odrv4 I__10195 (
            .O(N__56741),
            .I(\quad_counter0.n2112 ));
    LocalMux I__10194 (
            .O(N__56738),
            .I(\quad_counter0.n2112 ));
    InMux I__10193 (
            .O(N__56733),
            .I(bfn_16_7_0_));
    InMux I__10192 (
            .O(N__56730),
            .I(N__56725));
    InMux I__10191 (
            .O(N__56729),
            .I(N__56722));
    CascadeMux I__10190 (
            .O(N__56728),
            .I(N__56718));
    LocalMux I__10189 (
            .O(N__56725),
            .I(N__56714));
    LocalMux I__10188 (
            .O(N__56722),
            .I(N__56711));
    InMux I__10187 (
            .O(N__56721),
            .I(N__56708));
    InMux I__10186 (
            .O(N__56718),
            .I(N__56705));
    InMux I__10185 (
            .O(N__56717),
            .I(N__56702));
    Span4Mux_h I__10184 (
            .O(N__56714),
            .I(N__56695));
    Span4Mux_h I__10183 (
            .O(N__56711),
            .I(N__56695));
    LocalMux I__10182 (
            .O(N__56708),
            .I(N__56695));
    LocalMux I__10181 (
            .O(N__56705),
            .I(\c0.data_in_frame_16_2 ));
    LocalMux I__10180 (
            .O(N__56702),
            .I(\c0.data_in_frame_16_2 ));
    Odrv4 I__10179 (
            .O(N__56695),
            .I(\c0.data_in_frame_16_2 ));
    InMux I__10178 (
            .O(N__56688),
            .I(N__56684));
    InMux I__10177 (
            .O(N__56687),
            .I(N__56681));
    LocalMux I__10176 (
            .O(N__56684),
            .I(N__56678));
    LocalMux I__10175 (
            .O(N__56681),
            .I(N__56673));
    Span4Mux_v I__10174 (
            .O(N__56678),
            .I(N__56673));
    Odrv4 I__10173 (
            .O(N__56673),
            .I(\c0.n32241 ));
    InMux I__10172 (
            .O(N__56670),
            .I(N__56667));
    LocalMux I__10171 (
            .O(N__56667),
            .I(N__56664));
    Span4Mux_v I__10170 (
            .O(N__56664),
            .I(N__56661));
    Odrv4 I__10169 (
            .O(N__56661),
            .I(\c0.n33618 ));
    CascadeMux I__10168 (
            .O(N__56658),
            .I(\c0.n33618_cascade_ ));
    CascadeMux I__10167 (
            .O(N__56655),
            .I(N__56652));
    InMux I__10166 (
            .O(N__56652),
            .I(N__56649));
    LocalMux I__10165 (
            .O(N__56649),
            .I(\c0.n6462 ));
    CascadeMux I__10164 (
            .O(N__56646),
            .I(N__56643));
    InMux I__10163 (
            .O(N__56643),
            .I(N__56640));
    LocalMux I__10162 (
            .O(N__56640),
            .I(\c0.n22_adj_4670 ));
    InMux I__10161 (
            .O(N__56637),
            .I(N__56634));
    LocalMux I__10160 (
            .O(N__56634),
            .I(N__56631));
    Span4Mux_h I__10159 (
            .O(N__56631),
            .I(N__56628));
    Odrv4 I__10158 (
            .O(N__56628),
            .I(\c0.n33514 ));
    InMux I__10157 (
            .O(N__56625),
            .I(N__56619));
    InMux I__10156 (
            .O(N__56624),
            .I(N__56619));
    LocalMux I__10155 (
            .O(N__56619),
            .I(N__56616));
    Span4Mux_h I__10154 (
            .O(N__56616),
            .I(N__56613));
    Odrv4 I__10153 (
            .O(N__56613),
            .I(\c0.n18166 ));
    InMux I__10152 (
            .O(N__56610),
            .I(N__56605));
    InMux I__10151 (
            .O(N__56609),
            .I(N__56600));
    InMux I__10150 (
            .O(N__56608),
            .I(N__56600));
    LocalMux I__10149 (
            .O(N__56605),
            .I(N__56597));
    LocalMux I__10148 (
            .O(N__56600),
            .I(N__56594));
    Span4Mux_h I__10147 (
            .O(N__56597),
            .I(N__56591));
    Odrv4 I__10146 (
            .O(N__56594),
            .I(\c0.n31417 ));
    Odrv4 I__10145 (
            .O(N__56591),
            .I(\c0.n31417 ));
    InMux I__10144 (
            .O(N__56586),
            .I(N__56580));
    InMux I__10143 (
            .O(N__56585),
            .I(N__56580));
    LocalMux I__10142 (
            .O(N__56580),
            .I(N__56577));
    Span4Mux_h I__10141 (
            .O(N__56577),
            .I(N__56574));
    Span4Mux_h I__10140 (
            .O(N__56574),
            .I(N__56571));
    Odrv4 I__10139 (
            .O(N__56571),
            .I(\c0.n33833 ));
    InMux I__10138 (
            .O(N__56568),
            .I(N__56564));
    InMux I__10137 (
            .O(N__56567),
            .I(N__56561));
    LocalMux I__10136 (
            .O(N__56564),
            .I(N__56555));
    LocalMux I__10135 (
            .O(N__56561),
            .I(N__56555));
    InMux I__10134 (
            .O(N__56560),
            .I(N__56552));
    Span4Mux_h I__10133 (
            .O(N__56555),
            .I(N__56549));
    LocalMux I__10132 (
            .O(N__56552),
            .I(N__56546));
    Odrv4 I__10131 (
            .O(N__56549),
            .I(\c0.n18487 ));
    Odrv12 I__10130 (
            .O(N__56546),
            .I(\c0.n18487 ));
    InMux I__10129 (
            .O(N__56541),
            .I(N__56538));
    LocalMux I__10128 (
            .O(N__56538),
            .I(N__56535));
    Odrv4 I__10127 (
            .O(N__56535),
            .I(\c0.n33621 ));
    InMux I__10126 (
            .O(N__56532),
            .I(N__56529));
    LocalMux I__10125 (
            .O(N__56529),
            .I(\c0.n17702 ));
    CascadeMux I__10124 (
            .O(N__56526),
            .I(\c0.n17702_cascade_ ));
    InMux I__10123 (
            .O(N__56523),
            .I(bfn_16_6_0_));
    CascadeMux I__10122 (
            .O(N__56520),
            .I(N__56517));
    InMux I__10121 (
            .O(N__56517),
            .I(N__56513));
    InMux I__10120 (
            .O(N__56516),
            .I(N__56510));
    LocalMux I__10119 (
            .O(N__56513),
            .I(\c0.data_in_frame_14_4 ));
    LocalMux I__10118 (
            .O(N__56510),
            .I(\c0.data_in_frame_14_4 ));
    InMux I__10117 (
            .O(N__56505),
            .I(N__56502));
    LocalMux I__10116 (
            .O(N__56502),
            .I(N__56499));
    Odrv12 I__10115 (
            .O(N__56499),
            .I(\c0.n20_adj_4627 ));
    CascadeMux I__10114 (
            .O(N__56496),
            .I(N__56493));
    InMux I__10113 (
            .O(N__56493),
            .I(N__56489));
    CascadeMux I__10112 (
            .O(N__56492),
            .I(N__56485));
    LocalMux I__10111 (
            .O(N__56489),
            .I(N__56482));
    CascadeMux I__10110 (
            .O(N__56488),
            .I(N__56478));
    InMux I__10109 (
            .O(N__56485),
            .I(N__56475));
    Span4Mux_h I__10108 (
            .O(N__56482),
            .I(N__56472));
    InMux I__10107 (
            .O(N__56481),
            .I(N__56467));
    InMux I__10106 (
            .O(N__56478),
            .I(N__56467));
    LocalMux I__10105 (
            .O(N__56475),
            .I(\c0.data_in_frame_20_5 ));
    Odrv4 I__10104 (
            .O(N__56472),
            .I(\c0.data_in_frame_20_5 ));
    LocalMux I__10103 (
            .O(N__56467),
            .I(\c0.data_in_frame_20_5 ));
    InMux I__10102 (
            .O(N__56460),
            .I(N__56457));
    LocalMux I__10101 (
            .O(N__56457),
            .I(N__56451));
    InMux I__10100 (
            .O(N__56456),
            .I(N__56448));
    InMux I__10099 (
            .O(N__56455),
            .I(N__56443));
    InMux I__10098 (
            .O(N__56454),
            .I(N__56443));
    Span4Mux_h I__10097 (
            .O(N__56451),
            .I(N__56438));
    LocalMux I__10096 (
            .O(N__56448),
            .I(N__56438));
    LocalMux I__10095 (
            .O(N__56443),
            .I(N__56435));
    Span4Mux_v I__10094 (
            .O(N__56438),
            .I(N__56432));
    Odrv4 I__10093 (
            .O(N__56435),
            .I(\c0.n32357 ));
    Odrv4 I__10092 (
            .O(N__56432),
            .I(\c0.n32357 ));
    CascadeMux I__10091 (
            .O(N__56427),
            .I(\c0.n32026_cascade_ ));
    InMux I__10090 (
            .O(N__56424),
            .I(N__56421));
    LocalMux I__10089 (
            .O(N__56421),
            .I(\c0.n16_adj_4667 ));
    InMux I__10088 (
            .O(N__56418),
            .I(N__56415));
    LocalMux I__10087 (
            .O(N__56415),
            .I(N__56411));
    InMux I__10086 (
            .O(N__56414),
            .I(N__56408));
    Span4Mux_h I__10085 (
            .O(N__56411),
            .I(N__56405));
    LocalMux I__10084 (
            .O(N__56408),
            .I(N__56402));
    Odrv4 I__10083 (
            .O(N__56405),
            .I(\c0.n31940 ));
    Odrv4 I__10082 (
            .O(N__56402),
            .I(\c0.n31940 ));
    InMux I__10081 (
            .O(N__56397),
            .I(N__56394));
    LocalMux I__10080 (
            .O(N__56394),
            .I(\c0.n24_adj_4671 ));
    InMux I__10079 (
            .O(N__56391),
            .I(N__56385));
    InMux I__10078 (
            .O(N__56390),
            .I(N__56385));
    LocalMux I__10077 (
            .O(N__56385),
            .I(\c0.n32026 ));
    InMux I__10076 (
            .O(N__56382),
            .I(N__56376));
    InMux I__10075 (
            .O(N__56381),
            .I(N__56376));
    LocalMux I__10074 (
            .O(N__56376),
            .I(N__56373));
    Sp12to4 I__10073 (
            .O(N__56373),
            .I(N__56369));
    InMux I__10072 (
            .O(N__56372),
            .I(N__56365));
    Span12Mux_s8_v I__10071 (
            .O(N__56369),
            .I(N__56362));
    InMux I__10070 (
            .O(N__56368),
            .I(N__56359));
    LocalMux I__10069 (
            .O(N__56365),
            .I(\c0.data_in_frame_16_0 ));
    Odrv12 I__10068 (
            .O(N__56362),
            .I(\c0.data_in_frame_16_0 ));
    LocalMux I__10067 (
            .O(N__56359),
            .I(\c0.data_in_frame_16_0 ));
    InMux I__10066 (
            .O(N__56352),
            .I(N__56345));
    InMux I__10065 (
            .O(N__56351),
            .I(N__56345));
    InMux I__10064 (
            .O(N__56350),
            .I(N__56342));
    LocalMux I__10063 (
            .O(N__56345),
            .I(N__56339));
    LocalMux I__10062 (
            .O(N__56342),
            .I(N__56334));
    Span4Mux_h I__10061 (
            .O(N__56339),
            .I(N__56334));
    Odrv4 I__10060 (
            .O(N__56334),
            .I(\c0.n33601 ));
    InMux I__10059 (
            .O(N__56331),
            .I(N__56324));
    InMux I__10058 (
            .O(N__56330),
            .I(N__56324));
    InMux I__10057 (
            .O(N__56329),
            .I(N__56321));
    LocalMux I__10056 (
            .O(N__56324),
            .I(N__56318));
    LocalMux I__10055 (
            .O(N__56321),
            .I(N__56315));
    Odrv4 I__10054 (
            .O(N__56318),
            .I(\c0.n33827 ));
    Odrv4 I__10053 (
            .O(N__56315),
            .I(\c0.n33827 ));
    InMux I__10052 (
            .O(N__56310),
            .I(N__56307));
    LocalMux I__10051 (
            .O(N__56307),
            .I(\c0.n18974 ));
    CascadeMux I__10050 (
            .O(N__56304),
            .I(\c0.n18974_cascade_ ));
    CascadeMux I__10049 (
            .O(N__56301),
            .I(N__56297));
    InMux I__10048 (
            .O(N__56300),
            .I(N__56292));
    InMux I__10047 (
            .O(N__56297),
            .I(N__56292));
    LocalMux I__10046 (
            .O(N__56292),
            .I(N__56287));
    InMux I__10045 (
            .O(N__56291),
            .I(N__56282));
    InMux I__10044 (
            .O(N__56290),
            .I(N__56282));
    Odrv12 I__10043 (
            .O(N__56287),
            .I(\c0.data_in_frame_18_1 ));
    LocalMux I__10042 (
            .O(N__56282),
            .I(\c0.data_in_frame_18_1 ));
    CascadeMux I__10041 (
            .O(N__56277),
            .I(N__56274));
    InMux I__10040 (
            .O(N__56274),
            .I(N__56269));
    InMux I__10039 (
            .O(N__56273),
            .I(N__56264));
    InMux I__10038 (
            .O(N__56272),
            .I(N__56264));
    LocalMux I__10037 (
            .O(N__56269),
            .I(\c0.data_in_frame_20_3 ));
    LocalMux I__10036 (
            .O(N__56264),
            .I(\c0.data_in_frame_20_3 ));
    InMux I__10035 (
            .O(N__56259),
            .I(N__56256));
    LocalMux I__10034 (
            .O(N__56256),
            .I(\c0.n6_adj_4661 ));
    InMux I__10033 (
            .O(N__56253),
            .I(N__56250));
    LocalMux I__10032 (
            .O(N__56250),
            .I(N__56245));
    InMux I__10031 (
            .O(N__56249),
            .I(N__56242));
    InMux I__10030 (
            .O(N__56248),
            .I(N__56239));
    Span4Mux_h I__10029 (
            .O(N__56245),
            .I(N__56236));
    LocalMux I__10028 (
            .O(N__56242),
            .I(\c0.data_in_frame_12_2 ));
    LocalMux I__10027 (
            .O(N__56239),
            .I(\c0.data_in_frame_12_2 ));
    Odrv4 I__10026 (
            .O(N__56236),
            .I(\c0.data_in_frame_12_2 ));
    CascadeMux I__10025 (
            .O(N__56229),
            .I(N__56224));
    CascadeMux I__10024 (
            .O(N__56228),
            .I(N__56221));
    InMux I__10023 (
            .O(N__56227),
            .I(N__56217));
    InMux I__10022 (
            .O(N__56224),
            .I(N__56214));
    InMux I__10021 (
            .O(N__56221),
            .I(N__56209));
    InMux I__10020 (
            .O(N__56220),
            .I(N__56209));
    LocalMux I__10019 (
            .O(N__56217),
            .I(N__56206));
    LocalMux I__10018 (
            .O(N__56214),
            .I(\c0.data_in_frame_15_1 ));
    LocalMux I__10017 (
            .O(N__56209),
            .I(\c0.data_in_frame_15_1 ));
    Odrv4 I__10016 (
            .O(N__56206),
            .I(\c0.data_in_frame_15_1 ));
    CascadeMux I__10015 (
            .O(N__56199),
            .I(N__56196));
    InMux I__10014 (
            .O(N__56196),
            .I(N__56193));
    LocalMux I__10013 (
            .O(N__56193),
            .I(N__56189));
    InMux I__10012 (
            .O(N__56192),
            .I(N__56186));
    Odrv4 I__10011 (
            .O(N__56189),
            .I(\c0.n32087 ));
    LocalMux I__10010 (
            .O(N__56186),
            .I(\c0.n32087 ));
    CascadeMux I__10009 (
            .O(N__56181),
            .I(\c0.n33864_cascade_ ));
    InMux I__10008 (
            .O(N__56178),
            .I(N__56174));
    InMux I__10007 (
            .O(N__56177),
            .I(N__56171));
    LocalMux I__10006 (
            .O(N__56174),
            .I(\c0.n33979 ));
    LocalMux I__10005 (
            .O(N__56171),
            .I(\c0.n33979 ));
    InMux I__10004 (
            .O(N__56166),
            .I(N__56162));
    InMux I__10003 (
            .O(N__56165),
            .I(N__56159));
    LocalMux I__10002 (
            .O(N__56162),
            .I(N__56156));
    LocalMux I__10001 (
            .O(N__56159),
            .I(\c0.data_in_frame_28_3 ));
    Odrv4 I__10000 (
            .O(N__56156),
            .I(\c0.data_in_frame_28_3 ));
    InMux I__9999 (
            .O(N__56151),
            .I(N__56148));
    LocalMux I__9998 (
            .O(N__56148),
            .I(\c0.n34566 ));
    InMux I__9997 (
            .O(N__56145),
            .I(N__56142));
    LocalMux I__9996 (
            .O(N__56142),
            .I(\c0.n24_adj_4760 ));
    CascadeMux I__9995 (
            .O(N__56139),
            .I(N__56136));
    InMux I__9994 (
            .O(N__56136),
            .I(N__56130));
    InMux I__9993 (
            .O(N__56135),
            .I(N__56130));
    LocalMux I__9992 (
            .O(N__56130),
            .I(\c0.data_in_frame_28_1 ));
    CascadeMux I__9991 (
            .O(N__56127),
            .I(\c0.n17531_cascade_ ));
    CascadeMux I__9990 (
            .O(N__56124),
            .I(N__56121));
    InMux I__9989 (
            .O(N__56121),
            .I(N__56118));
    LocalMux I__9988 (
            .O(N__56118),
            .I(N__56115));
    Span4Mux_h I__9987 (
            .O(N__56115),
            .I(N__56110));
    InMux I__9986 (
            .O(N__56114),
            .I(N__56105));
    InMux I__9985 (
            .O(N__56113),
            .I(N__56105));
    Odrv4 I__9984 (
            .O(N__56110),
            .I(\c0.n17545 ));
    LocalMux I__9983 (
            .O(N__56105),
            .I(\c0.n17545 ));
    InMux I__9982 (
            .O(N__56100),
            .I(N__56097));
    LocalMux I__9981 (
            .O(N__56097),
            .I(N__56094));
    Odrv12 I__9980 (
            .O(N__56094),
            .I(\c0.n18588 ));
    CascadeMux I__9979 (
            .O(N__56091),
            .I(N__56088));
    InMux I__9978 (
            .O(N__56088),
            .I(N__56084));
    InMux I__9977 (
            .O(N__56087),
            .I(N__56081));
    LocalMux I__9976 (
            .O(N__56084),
            .I(\c0.data_in_frame_20_2 ));
    LocalMux I__9975 (
            .O(N__56081),
            .I(\c0.data_in_frame_20_2 ));
    CascadeMux I__9974 (
            .O(N__56076),
            .I(N__56072));
    CascadeMux I__9973 (
            .O(N__56075),
            .I(N__56069));
    InMux I__9972 (
            .O(N__56072),
            .I(N__56063));
    InMux I__9971 (
            .O(N__56069),
            .I(N__56063));
    CascadeMux I__9970 (
            .O(N__56068),
            .I(N__56060));
    LocalMux I__9969 (
            .O(N__56063),
            .I(N__56056));
    InMux I__9968 (
            .O(N__56060),
            .I(N__56053));
    InMux I__9967 (
            .O(N__56059),
            .I(N__56050));
    Span4Mux_h I__9966 (
            .O(N__56056),
            .I(N__56047));
    LocalMux I__9965 (
            .O(N__56053),
            .I(\c0.data_in_frame_15_3 ));
    LocalMux I__9964 (
            .O(N__56050),
            .I(\c0.data_in_frame_15_3 ));
    Odrv4 I__9963 (
            .O(N__56047),
            .I(\c0.data_in_frame_15_3 ));
    CascadeMux I__9962 (
            .O(N__56040),
            .I(N__56037));
    InMux I__9961 (
            .O(N__56037),
            .I(N__56034));
    LocalMux I__9960 (
            .O(N__56034),
            .I(N__56031));
    Odrv4 I__9959 (
            .O(N__56031),
            .I(\c0.n18373 ));
    InMux I__9958 (
            .O(N__56028),
            .I(N__56022));
    InMux I__9957 (
            .O(N__56027),
            .I(N__56022));
    LocalMux I__9956 (
            .O(N__56022),
            .I(N__56018));
    InMux I__9955 (
            .O(N__56021),
            .I(N__56015));
    Span4Mux_v I__9954 (
            .O(N__56018),
            .I(N__56012));
    LocalMux I__9953 (
            .O(N__56015),
            .I(\c0.data_in_frame_23_7 ));
    Odrv4 I__9952 (
            .O(N__56012),
            .I(\c0.data_in_frame_23_7 ));
    InMux I__9951 (
            .O(N__56007),
            .I(N__56004));
    LocalMux I__9950 (
            .O(N__56004),
            .I(N__56001));
    Span4Mux_h I__9949 (
            .O(N__56001),
            .I(N__55998));
    Odrv4 I__9948 (
            .O(N__55998),
            .I(\c0.n33813 ));
    InMux I__9947 (
            .O(N__55995),
            .I(N__55992));
    LocalMux I__9946 (
            .O(N__55992),
            .I(N__55988));
    CascadeMux I__9945 (
            .O(N__55991),
            .I(N__55983));
    Span4Mux_h I__9944 (
            .O(N__55988),
            .I(N__55980));
    InMux I__9943 (
            .O(N__55987),
            .I(N__55977));
    InMux I__9942 (
            .O(N__55986),
            .I(N__55974));
    InMux I__9941 (
            .O(N__55983),
            .I(N__55971));
    Span4Mux_h I__9940 (
            .O(N__55980),
            .I(N__55968));
    LocalMux I__9939 (
            .O(N__55977),
            .I(N__55963));
    LocalMux I__9938 (
            .O(N__55974),
            .I(N__55963));
    LocalMux I__9937 (
            .O(N__55971),
            .I(\c0.data_in_frame_13_7 ));
    Odrv4 I__9936 (
            .O(N__55968),
            .I(\c0.data_in_frame_13_7 ));
    Odrv12 I__9935 (
            .O(N__55963),
            .I(\c0.data_in_frame_13_7 ));
    InMux I__9934 (
            .O(N__55956),
            .I(N__55953));
    LocalMux I__9933 (
            .O(N__55953),
            .I(N__55950));
    Odrv4 I__9932 (
            .O(N__55950),
            .I(\c0.n14_adj_4538 ));
    CascadeMux I__9931 (
            .O(N__55947),
            .I(\c0.n34727_cascade_ ));
    InMux I__9930 (
            .O(N__55944),
            .I(N__55941));
    LocalMux I__9929 (
            .O(N__55941),
            .I(N__55938));
    Odrv4 I__9928 (
            .O(N__55938),
            .I(\c0.n29_adj_4761 ));
    CascadeMux I__9927 (
            .O(N__55935),
            .I(N__55923));
    CascadeMux I__9926 (
            .O(N__55934),
            .I(N__55920));
    CascadeMux I__9925 (
            .O(N__55933),
            .I(N__55917));
    CascadeMux I__9924 (
            .O(N__55932),
            .I(N__55913));
    InMux I__9923 (
            .O(N__55931),
            .I(N__55908));
    InMux I__9922 (
            .O(N__55930),
            .I(N__55908));
    CascadeMux I__9921 (
            .O(N__55929),
            .I(N__55905));
    CascadeMux I__9920 (
            .O(N__55928),
            .I(N__55902));
    CascadeMux I__9919 (
            .O(N__55927),
            .I(N__55899));
    InMux I__9918 (
            .O(N__55926),
            .I(N__55895));
    InMux I__9917 (
            .O(N__55923),
            .I(N__55892));
    InMux I__9916 (
            .O(N__55920),
            .I(N__55887));
    InMux I__9915 (
            .O(N__55917),
            .I(N__55887));
    InMux I__9914 (
            .O(N__55916),
            .I(N__55882));
    InMux I__9913 (
            .O(N__55913),
            .I(N__55882));
    LocalMux I__9912 (
            .O(N__55908),
            .I(N__55879));
    InMux I__9911 (
            .O(N__55905),
            .I(N__55876));
    InMux I__9910 (
            .O(N__55902),
            .I(N__55869));
    InMux I__9909 (
            .O(N__55899),
            .I(N__55869));
    InMux I__9908 (
            .O(N__55898),
            .I(N__55869));
    LocalMux I__9907 (
            .O(N__55895),
            .I(N__55866));
    LocalMux I__9906 (
            .O(N__55892),
            .I(N__55863));
    LocalMux I__9905 (
            .O(N__55887),
            .I(N__55860));
    LocalMux I__9904 (
            .O(N__55882),
            .I(N__55855));
    Span4Mux_v I__9903 (
            .O(N__55879),
            .I(N__55855));
    LocalMux I__9902 (
            .O(N__55876),
            .I(N__55852));
    LocalMux I__9901 (
            .O(N__55869),
            .I(N__55849));
    Span4Mux_h I__9900 (
            .O(N__55866),
            .I(N__55846));
    Span4Mux_h I__9899 (
            .O(N__55863),
            .I(N__55841));
    Span4Mux_v I__9898 (
            .O(N__55860),
            .I(N__55841));
    Span4Mux_v I__9897 (
            .O(N__55855),
            .I(N__55838));
    Span4Mux_v I__9896 (
            .O(N__55852),
            .I(N__55835));
    Span4Mux_h I__9895 (
            .O(N__55849),
            .I(N__55830));
    Span4Mux_h I__9894 (
            .O(N__55846),
            .I(N__55830));
    Span4Mux_v I__9893 (
            .O(N__55841),
            .I(N__55827));
    Span4Mux_v I__9892 (
            .O(N__55838),
            .I(N__55824));
    Span4Mux_h I__9891 (
            .O(N__55835),
            .I(N__55819));
    Span4Mux_v I__9890 (
            .O(N__55830),
            .I(N__55819));
    Span4Mux_v I__9889 (
            .O(N__55827),
            .I(N__55814));
    Span4Mux_h I__9888 (
            .O(N__55824),
            .I(N__55814));
    Span4Mux_v I__9887 (
            .O(N__55819),
            .I(N__55811));
    Odrv4 I__9886 (
            .O(N__55814),
            .I(r_Rx_Data));
    Odrv4 I__9885 (
            .O(N__55811),
            .I(r_Rx_Data));
    CascadeMux I__9884 (
            .O(N__55806),
            .I(\c0.rx.n35769_cascade_ ));
    InMux I__9883 (
            .O(N__55803),
            .I(N__55795));
    InMux I__9882 (
            .O(N__55802),
            .I(N__55795));
    InMux I__9881 (
            .O(N__55801),
            .I(N__55792));
    InMux I__9880 (
            .O(N__55800),
            .I(N__55789));
    LocalMux I__9879 (
            .O(N__55795),
            .I(\c0.rx.r_SM_Main_2_N_3687_0 ));
    LocalMux I__9878 (
            .O(N__55792),
            .I(\c0.rx.r_SM_Main_2_N_3687_0 ));
    LocalMux I__9877 (
            .O(N__55789),
            .I(\c0.rx.r_SM_Main_2_N_3687_0 ));
    InMux I__9876 (
            .O(N__55782),
            .I(N__55779));
    LocalMux I__9875 (
            .O(N__55779),
            .I(\c0.rx.n35738 ));
    InMux I__9874 (
            .O(N__55776),
            .I(N__55771));
    InMux I__9873 (
            .O(N__55775),
            .I(N__55768));
    CascadeMux I__9872 (
            .O(N__55774),
            .I(N__55765));
    LocalMux I__9871 (
            .O(N__55771),
            .I(N__55762));
    LocalMux I__9870 (
            .O(N__55768),
            .I(N__55759));
    InMux I__9869 (
            .O(N__55765),
            .I(N__55756));
    Span4Mux_h I__9868 (
            .O(N__55762),
            .I(N__55753));
    Span4Mux_h I__9867 (
            .O(N__55759),
            .I(N__55750));
    LocalMux I__9866 (
            .O(N__55756),
            .I(\c0.data_in_frame_3_4 ));
    Odrv4 I__9865 (
            .O(N__55753),
            .I(\c0.data_in_frame_3_4 ));
    Odrv4 I__9864 (
            .O(N__55750),
            .I(\c0.data_in_frame_3_4 ));
    CascadeMux I__9863 (
            .O(N__55743),
            .I(\c0.rx.n33223_cascade_ ));
    InMux I__9862 (
            .O(N__55740),
            .I(N__55737));
    LocalMux I__9861 (
            .O(N__55737),
            .I(\c0.rx.n35950 ));
    InMux I__9860 (
            .O(N__55734),
            .I(N__55730));
    InMux I__9859 (
            .O(N__55733),
            .I(N__55725));
    LocalMux I__9858 (
            .O(N__55730),
            .I(N__55722));
    InMux I__9857 (
            .O(N__55729),
            .I(N__55719));
    CascadeMux I__9856 (
            .O(N__55728),
            .I(N__55716));
    LocalMux I__9855 (
            .O(N__55725),
            .I(N__55709));
    Span4Mux_v I__9854 (
            .O(N__55722),
            .I(N__55709));
    LocalMux I__9853 (
            .O(N__55719),
            .I(N__55709));
    InMux I__9852 (
            .O(N__55716),
            .I(N__55706));
    Span4Mux_h I__9851 (
            .O(N__55709),
            .I(N__55703));
    LocalMux I__9850 (
            .O(N__55706),
            .I(\c0.data_in_frame_13_1 ));
    Odrv4 I__9849 (
            .O(N__55703),
            .I(\c0.data_in_frame_13_1 ));
    CascadeMux I__9848 (
            .O(N__55698),
            .I(\c0.n33233_cascade_ ));
    InMux I__9847 (
            .O(N__55695),
            .I(N__55692));
    LocalMux I__9846 (
            .O(N__55692),
            .I(N__55688));
    CascadeMux I__9845 (
            .O(N__55691),
            .I(N__55684));
    Span4Mux_v I__9844 (
            .O(N__55688),
            .I(N__55681));
    InMux I__9843 (
            .O(N__55687),
            .I(N__55676));
    InMux I__9842 (
            .O(N__55684),
            .I(N__55676));
    Span4Mux_v I__9841 (
            .O(N__55681),
            .I(N__55673));
    LocalMux I__9840 (
            .O(N__55676),
            .I(N__55670));
    Odrv4 I__9839 (
            .O(N__55673),
            .I(\c0.n63_adj_4633 ));
    Odrv4 I__9838 (
            .O(N__55670),
            .I(\c0.n63_adj_4633 ));
    InMux I__9837 (
            .O(N__55665),
            .I(N__55662));
    LocalMux I__9836 (
            .O(N__55662),
            .I(N__55659));
    Odrv4 I__9835 (
            .O(N__55659),
            .I(\c0.n35633 ));
    CascadeMux I__9834 (
            .O(N__55656),
            .I(N__55653));
    InMux I__9833 (
            .O(N__55653),
            .I(N__55650));
    LocalMux I__9832 (
            .O(N__55650),
            .I(N__55647));
    Span4Mux_v I__9831 (
            .O(N__55647),
            .I(N__55643));
    InMux I__9830 (
            .O(N__55646),
            .I(N__55640));
    Odrv4 I__9829 (
            .O(N__55643),
            .I(\c0.n27708 ));
    LocalMux I__9828 (
            .O(N__55640),
            .I(\c0.n27708 ));
    InMux I__9827 (
            .O(N__55635),
            .I(N__55632));
    LocalMux I__9826 (
            .O(N__55632),
            .I(n35992));
    CascadeMux I__9825 (
            .O(N__55629),
            .I(\c0.rx.r_SM_Main_2_N_3681_2_cascade_ ));
    InMux I__9824 (
            .O(N__55626),
            .I(N__55620));
    InMux I__9823 (
            .O(N__55625),
            .I(N__55617));
    InMux I__9822 (
            .O(N__55624),
            .I(N__55614));
    InMux I__9821 (
            .O(N__55623),
            .I(N__55610));
    LocalMux I__9820 (
            .O(N__55620),
            .I(N__55607));
    LocalMux I__9819 (
            .O(N__55617),
            .I(N__55603));
    LocalMux I__9818 (
            .O(N__55614),
            .I(N__55600));
    InMux I__9817 (
            .O(N__55613),
            .I(N__55597));
    LocalMux I__9816 (
            .O(N__55610),
            .I(N__55592));
    Span4Mux_v I__9815 (
            .O(N__55607),
            .I(N__55592));
    InMux I__9814 (
            .O(N__55606),
            .I(N__55589));
    Span4Mux_v I__9813 (
            .O(N__55603),
            .I(N__55584));
    Span4Mux_h I__9812 (
            .O(N__55600),
            .I(N__55584));
    LocalMux I__9811 (
            .O(N__55597),
            .I(N__55581));
    Span4Mux_h I__9810 (
            .O(N__55592),
            .I(N__55578));
    LocalMux I__9809 (
            .O(N__55589),
            .I(N__55571));
    Span4Mux_h I__9808 (
            .O(N__55584),
            .I(N__55571));
    Span4Mux_v I__9807 (
            .O(N__55581),
            .I(N__55571));
    Odrv4 I__9806 (
            .O(N__55578),
            .I(\c0.rx.r_Bit_Index_0 ));
    Odrv4 I__9805 (
            .O(N__55571),
            .I(\c0.rx.r_Bit_Index_0 ));
    CascadeMux I__9804 (
            .O(N__55566),
            .I(\c0.rx.n34091_cascade_ ));
    InMux I__9803 (
            .O(N__55563),
            .I(N__55559));
    InMux I__9802 (
            .O(N__55562),
            .I(N__55554));
    LocalMux I__9801 (
            .O(N__55559),
            .I(N__55551));
    InMux I__9800 (
            .O(N__55558),
            .I(N__55545));
    InMux I__9799 (
            .O(N__55557),
            .I(N__55542));
    LocalMux I__9798 (
            .O(N__55554),
            .I(N__55539));
    Span4Mux_v I__9797 (
            .O(N__55551),
            .I(N__55536));
    InMux I__9796 (
            .O(N__55550),
            .I(N__55533));
    InMux I__9795 (
            .O(N__55549),
            .I(N__55530));
    InMux I__9794 (
            .O(N__55548),
            .I(N__55527));
    LocalMux I__9793 (
            .O(N__55545),
            .I(N__55520));
    LocalMux I__9792 (
            .O(N__55542),
            .I(N__55520));
    Span12Mux_v I__9791 (
            .O(N__55539),
            .I(N__55520));
    Span4Mux_h I__9790 (
            .O(N__55536),
            .I(N__55517));
    LocalMux I__9789 (
            .O(N__55533),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__9788 (
            .O(N__55530),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__9787 (
            .O(N__55527),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv12 I__9786 (
            .O(N__55520),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv4 I__9785 (
            .O(N__55517),
            .I(\c0.rx.r_Bit_Index_1 ));
    InMux I__9784 (
            .O(N__55506),
            .I(N__55503));
    LocalMux I__9783 (
            .O(N__55503),
            .I(\c0.rx.n28401 ));
    InMux I__9782 (
            .O(N__55500),
            .I(N__55497));
    LocalMux I__9781 (
            .O(N__55497),
            .I(\c0.rx.n29888 ));
    InMux I__9780 (
            .O(N__55494),
            .I(N__55491));
    LocalMux I__9779 (
            .O(N__55491),
            .I(N__55486));
    InMux I__9778 (
            .O(N__55490),
            .I(N__55481));
    InMux I__9777 (
            .O(N__55489),
            .I(N__55481));
    Odrv4 I__9776 (
            .O(N__55486),
            .I(\c0.rx.n34091 ));
    LocalMux I__9775 (
            .O(N__55481),
            .I(\c0.rx.n34091 ));
    InMux I__9774 (
            .O(N__55476),
            .I(N__55473));
    LocalMux I__9773 (
            .O(N__55473),
            .I(N__55470));
    Span4Mux_h I__9772 (
            .O(N__55470),
            .I(N__55467));
    Span4Mux_h I__9771 (
            .O(N__55467),
            .I(N__55464));
    Odrv4 I__9770 (
            .O(N__55464),
            .I(\c0.rx.n3821 ));
    CascadeMux I__9769 (
            .O(N__55461),
            .I(\c0.rx.n29888_cascade_ ));
    InMux I__9768 (
            .O(N__55458),
            .I(N__55455));
    LocalMux I__9767 (
            .O(N__55455),
            .I(N__55452));
    Span4Mux_h I__9766 (
            .O(N__55452),
            .I(N__55449));
    Span4Mux_h I__9765 (
            .O(N__55449),
            .I(N__55443));
    InMux I__9764 (
            .O(N__55448),
            .I(N__55440));
    InMux I__9763 (
            .O(N__55447),
            .I(N__55437));
    InMux I__9762 (
            .O(N__55446),
            .I(N__55432));
    Span4Mux_h I__9761 (
            .O(N__55443),
            .I(N__55429));
    LocalMux I__9760 (
            .O(N__55440),
            .I(N__55424));
    LocalMux I__9759 (
            .O(N__55437),
            .I(N__55424));
    InMux I__9758 (
            .O(N__55436),
            .I(N__55421));
    InMux I__9757 (
            .O(N__55435),
            .I(N__55418));
    LocalMux I__9756 (
            .O(N__55432),
            .I(\c0.rx.r_Bit_Index_2 ));
    Odrv4 I__9755 (
            .O(N__55429),
            .I(\c0.rx.r_Bit_Index_2 ));
    Odrv12 I__9754 (
            .O(N__55424),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__9753 (
            .O(N__55421),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__9752 (
            .O(N__55418),
            .I(\c0.rx.r_Bit_Index_2 ));
    CascadeMux I__9751 (
            .O(N__55407),
            .I(N__55404));
    InMux I__9750 (
            .O(N__55404),
            .I(N__55401));
    LocalMux I__9749 (
            .O(N__55401),
            .I(N__55395));
    InMux I__9748 (
            .O(N__55400),
            .I(N__55390));
    InMux I__9747 (
            .O(N__55399),
            .I(N__55390));
    CascadeMux I__9746 (
            .O(N__55398),
            .I(N__55387));
    Span4Mux_v I__9745 (
            .O(N__55395),
            .I(N__55382));
    LocalMux I__9744 (
            .O(N__55390),
            .I(N__55382));
    InMux I__9743 (
            .O(N__55387),
            .I(N__55379));
    Span4Mux_h I__9742 (
            .O(N__55382),
            .I(N__55376));
    LocalMux I__9741 (
            .O(N__55379),
            .I(\c0.data_in_frame_5_7 ));
    Odrv4 I__9740 (
            .O(N__55376),
            .I(\c0.data_in_frame_5_7 ));
    CascadeMux I__9739 (
            .O(N__55371),
            .I(N__55367));
    InMux I__9738 (
            .O(N__55370),
            .I(N__55364));
    InMux I__9737 (
            .O(N__55367),
            .I(N__55361));
    LocalMux I__9736 (
            .O(N__55364),
            .I(N__55358));
    LocalMux I__9735 (
            .O(N__55361),
            .I(N__55353));
    Span4Mux_h I__9734 (
            .O(N__55358),
            .I(N__55353));
    Span4Mux_h I__9733 (
            .O(N__55353),
            .I(N__55350));
    Odrv4 I__9732 (
            .O(N__55350),
            .I(\c0.n5024 ));
    CascadeMux I__9731 (
            .O(N__55347),
            .I(n35991_cascade_));
    InMux I__9730 (
            .O(N__55344),
            .I(N__55341));
    LocalMux I__9729 (
            .O(N__55341),
            .I(\c0.n11_adj_4626 ));
    CascadeMux I__9728 (
            .O(N__55338),
            .I(\c0.rx.n28401_cascade_ ));
    CascadeMux I__9727 (
            .O(N__55335),
            .I(n28381_cascade_));
    InMux I__9726 (
            .O(N__55332),
            .I(N__55329));
    LocalMux I__9725 (
            .O(N__55329),
            .I(n1));
    InMux I__9724 (
            .O(N__55326),
            .I(N__55322));
    InMux I__9723 (
            .O(N__55325),
            .I(N__55319));
    LocalMux I__9722 (
            .O(N__55322),
            .I(data_out_frame_7_6));
    LocalMux I__9721 (
            .O(N__55319),
            .I(data_out_frame_7_6));
    InMux I__9720 (
            .O(N__55314),
            .I(N__55308));
    InMux I__9719 (
            .O(N__55313),
            .I(N__55308));
    LocalMux I__9718 (
            .O(N__55308),
            .I(data_out_frame_6_2));
    InMux I__9717 (
            .O(N__55305),
            .I(N__55302));
    LocalMux I__9716 (
            .O(N__55302),
            .I(\c0.n5_adj_4511 ));
    InMux I__9715 (
            .O(N__55299),
            .I(N__55296));
    LocalMux I__9714 (
            .O(N__55296),
            .I(N__55293));
    Odrv4 I__9713 (
            .O(N__55293),
            .I(\c0.n36209 ));
    InMux I__9712 (
            .O(N__55290),
            .I(N__55284));
    InMux I__9711 (
            .O(N__55289),
            .I(N__55284));
    LocalMux I__9710 (
            .O(N__55284),
            .I(data_out_frame_8_1));
    CascadeMux I__9709 (
            .O(N__55281),
            .I(\c0.n36212_cascade_ ));
    InMux I__9708 (
            .O(N__55278),
            .I(N__55275));
    LocalMux I__9707 (
            .O(N__55275),
            .I(N__55272));
    Span4Mux_v I__9706 (
            .O(N__55272),
            .I(N__55269));
    Odrv4 I__9705 (
            .O(N__55269),
            .I(n36092));
    InMux I__9704 (
            .O(N__55266),
            .I(N__55263));
    LocalMux I__9703 (
            .O(N__55263),
            .I(N__55260));
    Odrv4 I__9702 (
            .O(N__55260),
            .I(n36088));
    InMux I__9701 (
            .O(N__55257),
            .I(N__55254));
    LocalMux I__9700 (
            .O(N__55254),
            .I(N__55251));
    Odrv4 I__9699 (
            .O(N__55251),
            .I(n35820));
    InMux I__9698 (
            .O(N__55248),
            .I(N__55245));
    LocalMux I__9697 (
            .O(N__55245),
            .I(N__55242));
    Odrv4 I__9696 (
            .O(N__55242),
            .I(\c0.n17959 ));
    CascadeMux I__9695 (
            .O(N__55239),
            .I(N__55236));
    InMux I__9694 (
            .O(N__55236),
            .I(N__55232));
    InMux I__9693 (
            .O(N__55235),
            .I(N__55228));
    LocalMux I__9692 (
            .O(N__55232),
            .I(N__55225));
    InMux I__9691 (
            .O(N__55231),
            .I(N__55222));
    LocalMux I__9690 (
            .O(N__55228),
            .I(N__55219));
    Span4Mux_h I__9689 (
            .O(N__55225),
            .I(N__55216));
    LocalMux I__9688 (
            .O(N__55222),
            .I(N__55213));
    Span4Mux_h I__9687 (
            .O(N__55219),
            .I(N__55210));
    Span4Mux_h I__9686 (
            .O(N__55216),
            .I(N__55207));
    Span12Mux_v I__9685 (
            .O(N__55213),
            .I(N__55204));
    Odrv4 I__9684 (
            .O(N__55210),
            .I(\c0.n30906 ));
    Odrv4 I__9683 (
            .O(N__55207),
            .I(\c0.n30906 ));
    Odrv12 I__9682 (
            .O(N__55204),
            .I(\c0.n30906 ));
    InMux I__9681 (
            .O(N__55197),
            .I(N__55191));
    InMux I__9680 (
            .O(N__55196),
            .I(N__55191));
    LocalMux I__9679 (
            .O(N__55191),
            .I(data_out_frame_10_1));
    InMux I__9678 (
            .O(N__55188),
            .I(N__55182));
    InMux I__9677 (
            .O(N__55187),
            .I(N__55182));
    LocalMux I__9676 (
            .O(N__55182),
            .I(data_out_frame_11_1));
    InMux I__9675 (
            .O(N__55179),
            .I(N__55176));
    LocalMux I__9674 (
            .O(N__55176),
            .I(N__55173));
    Odrv4 I__9673 (
            .O(N__55173),
            .I(\c0.n35833 ));
    InMux I__9672 (
            .O(N__55170),
            .I(N__55167));
    LocalMux I__9671 (
            .O(N__55167),
            .I(n35835));
    InMux I__9670 (
            .O(N__55164),
            .I(N__55158));
    InMux I__9669 (
            .O(N__55163),
            .I(N__55158));
    LocalMux I__9668 (
            .O(N__55158),
            .I(data_out_frame_9_0));
    InMux I__9667 (
            .O(N__55155),
            .I(N__55152));
    LocalMux I__9666 (
            .O(N__55152),
            .I(N__55149));
    Odrv12 I__9665 (
            .O(N__55149),
            .I(\c0.n11 ));
    CascadeMux I__9664 (
            .O(N__55146),
            .I(\c0.n36200_cascade_ ));
    InMux I__9663 (
            .O(N__55143),
            .I(N__55140));
    LocalMux I__9662 (
            .O(N__55140),
            .I(N__55136));
    CascadeMux I__9661 (
            .O(N__55139),
            .I(N__55133));
    Span4Mux_h I__9660 (
            .O(N__55136),
            .I(N__55130));
    InMux I__9659 (
            .O(N__55133),
            .I(N__55127));
    Span4Mux_h I__9658 (
            .O(N__55130),
            .I(N__55124));
    LocalMux I__9657 (
            .O(N__55127),
            .I(r_Tx_Data_3));
    Odrv4 I__9656 (
            .O(N__55124),
            .I(r_Tx_Data_3));
    InMux I__9655 (
            .O(N__55119),
            .I(N__55115));
    InMux I__9654 (
            .O(N__55118),
            .I(N__55112));
    LocalMux I__9653 (
            .O(N__55115),
            .I(N__55109));
    LocalMux I__9652 (
            .O(N__55112),
            .I(data_out_frame_12_0));
    Odrv4 I__9651 (
            .O(N__55109),
            .I(data_out_frame_12_0));
    InMux I__9650 (
            .O(N__55104),
            .I(N__55100));
    InMux I__9649 (
            .O(N__55103),
            .I(N__55097));
    LocalMux I__9648 (
            .O(N__55100),
            .I(data_out_frame_13_0));
    LocalMux I__9647 (
            .O(N__55097),
            .I(data_out_frame_13_0));
    InMux I__9646 (
            .O(N__55092),
            .I(N__55088));
    InMux I__9645 (
            .O(N__55091),
            .I(N__55085));
    LocalMux I__9644 (
            .O(N__55088),
            .I(\c0.byte_transmit_counter_7 ));
    LocalMux I__9643 (
            .O(N__55085),
            .I(\c0.byte_transmit_counter_7 ));
    InMux I__9642 (
            .O(N__55080),
            .I(N__55076));
    InMux I__9641 (
            .O(N__55079),
            .I(N__55073));
    LocalMux I__9640 (
            .O(N__55076),
            .I(\c0.byte_transmit_counter_6 ));
    LocalMux I__9639 (
            .O(N__55073),
            .I(\c0.byte_transmit_counter_6 ));
    CascadeMux I__9638 (
            .O(N__55068),
            .I(N__55065));
    InMux I__9637 (
            .O(N__55065),
            .I(N__55056));
    InMux I__9636 (
            .O(N__55064),
            .I(N__55056));
    InMux I__9635 (
            .O(N__55063),
            .I(N__55056));
    LocalMux I__9634 (
            .O(N__55056),
            .I(N__55053));
    Odrv4 I__9633 (
            .O(N__55053),
            .I(\c0.n4_adj_4646 ));
    CascadeMux I__9632 (
            .O(N__55050),
            .I(N__55046));
    CascadeMux I__9631 (
            .O(N__55049),
            .I(N__55043));
    InMux I__9630 (
            .O(N__55046),
            .I(N__55040));
    InMux I__9629 (
            .O(N__55043),
            .I(N__55037));
    LocalMux I__9628 (
            .O(N__55040),
            .I(N__55034));
    LocalMux I__9627 (
            .O(N__55037),
            .I(N__55029));
    Span4Mux_h I__9626 (
            .O(N__55034),
            .I(N__55029));
    Odrv4 I__9625 (
            .O(N__55029),
            .I(r_Tx_Data_7));
    CascadeMux I__9624 (
            .O(N__55026),
            .I(n36084_cascade_));
    InMux I__9623 (
            .O(N__55023),
            .I(N__55020));
    LocalMux I__9622 (
            .O(N__55020),
            .I(N__55017));
    Span4Mux_h I__9621 (
            .O(N__55017),
            .I(N__55014));
    Odrv4 I__9620 (
            .O(N__55014),
            .I(n10_adj_4804));
    InMux I__9619 (
            .O(N__55011),
            .I(N__55008));
    LocalMux I__9618 (
            .O(N__55008),
            .I(N__55004));
    InMux I__9617 (
            .O(N__55007),
            .I(N__55001));
    Span12Mux_h I__9616 (
            .O(N__55004),
            .I(N__54998));
    LocalMux I__9615 (
            .O(N__55001),
            .I(r_Tx_Data_0));
    Odrv12 I__9614 (
            .O(N__54998),
            .I(r_Tx_Data_0));
    InMux I__9613 (
            .O(N__54993),
            .I(N__54990));
    LocalMux I__9612 (
            .O(N__54990),
            .I(N__54987));
    Odrv4 I__9611 (
            .O(N__54987),
            .I(\quad_counter0.n3503 ));
    InMux I__9610 (
            .O(N__54984),
            .I(bfn_15_11_0_));
    InMux I__9609 (
            .O(N__54981),
            .I(N__54977));
    InMux I__9608 (
            .O(N__54980),
            .I(N__54974));
    LocalMux I__9607 (
            .O(N__54977),
            .I(N__54968));
    LocalMux I__9606 (
            .O(N__54974),
            .I(N__54968));
    InMux I__9605 (
            .O(N__54973),
            .I(N__54965));
    Odrv4 I__9604 (
            .O(N__54968),
            .I(\quad_counter0.n3403 ));
    LocalMux I__9603 (
            .O(N__54965),
            .I(\quad_counter0.n3403 ));
    InMux I__9602 (
            .O(N__54960),
            .I(\quad_counter0.n30441 ));
    InMux I__9601 (
            .O(N__54957),
            .I(N__54953));
    InMux I__9600 (
            .O(N__54956),
            .I(N__54950));
    LocalMux I__9599 (
            .O(N__54953),
            .I(N__54944));
    LocalMux I__9598 (
            .O(N__54950),
            .I(N__54944));
    InMux I__9597 (
            .O(N__54949),
            .I(N__54941));
    Odrv12 I__9596 (
            .O(N__54944),
            .I(\quad_counter0.n3402 ));
    LocalMux I__9595 (
            .O(N__54941),
            .I(\quad_counter0.n3402 ));
    InMux I__9594 (
            .O(N__54936),
            .I(\quad_counter0.n30442 ));
    InMux I__9593 (
            .O(N__54933),
            .I(N__54928));
    InMux I__9592 (
            .O(N__54932),
            .I(N__54925));
    CascadeMux I__9591 (
            .O(N__54931),
            .I(N__54922));
    LocalMux I__9590 (
            .O(N__54928),
            .I(N__54917));
    LocalMux I__9589 (
            .O(N__54925),
            .I(N__54917));
    InMux I__9588 (
            .O(N__54922),
            .I(N__54914));
    Odrv4 I__9587 (
            .O(N__54917),
            .I(\quad_counter0.n3401 ));
    LocalMux I__9586 (
            .O(N__54914),
            .I(\quad_counter0.n3401 ));
    InMux I__9585 (
            .O(N__54909),
            .I(\quad_counter0.n30443 ));
    InMux I__9584 (
            .O(N__54906),
            .I(N__54902));
    InMux I__9583 (
            .O(N__54905),
            .I(N__54899));
    LocalMux I__9582 (
            .O(N__54902),
            .I(N__54893));
    LocalMux I__9581 (
            .O(N__54899),
            .I(N__54893));
    InMux I__9580 (
            .O(N__54898),
            .I(N__54890));
    Odrv4 I__9579 (
            .O(N__54893),
            .I(\quad_counter0.n3400 ));
    LocalMux I__9578 (
            .O(N__54890),
            .I(\quad_counter0.n3400 ));
    InMux I__9577 (
            .O(N__54885),
            .I(\quad_counter0.n30444 ));
    InMux I__9576 (
            .O(N__54882),
            .I(N__54878));
    InMux I__9575 (
            .O(N__54881),
            .I(N__54875));
    LocalMux I__9574 (
            .O(N__54878),
            .I(N__54869));
    LocalMux I__9573 (
            .O(N__54875),
            .I(N__54869));
    InMux I__9572 (
            .O(N__54874),
            .I(N__54866));
    Odrv12 I__9571 (
            .O(N__54869),
            .I(\quad_counter0.n3399 ));
    LocalMux I__9570 (
            .O(N__54866),
            .I(\quad_counter0.n3399 ));
    InMux I__9569 (
            .O(N__54861),
            .I(\quad_counter0.n30445 ));
    InMux I__9568 (
            .O(N__54858),
            .I(N__54854));
    InMux I__9567 (
            .O(N__54857),
            .I(N__54851));
    LocalMux I__9566 (
            .O(N__54854),
            .I(N__54845));
    LocalMux I__9565 (
            .O(N__54851),
            .I(N__54845));
    InMux I__9564 (
            .O(N__54850),
            .I(N__54842));
    Odrv4 I__9563 (
            .O(N__54845),
            .I(\quad_counter0.n3398 ));
    LocalMux I__9562 (
            .O(N__54842),
            .I(\quad_counter0.n3398 ));
    CascadeMux I__9561 (
            .O(N__54837),
            .I(N__54818));
    CascadeMux I__9560 (
            .O(N__54836),
            .I(N__54815));
    CascadeMux I__9559 (
            .O(N__54835),
            .I(N__54812));
    CascadeMux I__9558 (
            .O(N__54834),
            .I(N__54809));
    CascadeMux I__9557 (
            .O(N__54833),
            .I(N__54806));
    CascadeMux I__9556 (
            .O(N__54832),
            .I(N__54803));
    CascadeMux I__9555 (
            .O(N__54831),
            .I(N__54800));
    CascadeMux I__9554 (
            .O(N__54830),
            .I(N__54797));
    CascadeMux I__9553 (
            .O(N__54829),
            .I(N__54794));
    CascadeMux I__9552 (
            .O(N__54828),
            .I(N__54791));
    CascadeMux I__9551 (
            .O(N__54827),
            .I(N__54788));
    CascadeMux I__9550 (
            .O(N__54826),
            .I(N__54785));
    CascadeMux I__9549 (
            .O(N__54825),
            .I(N__54782));
    CascadeMux I__9548 (
            .O(N__54824),
            .I(N__54779));
    CascadeMux I__9547 (
            .O(N__54823),
            .I(N__54776));
    CascadeMux I__9546 (
            .O(N__54822),
            .I(N__54773));
    CascadeMux I__9545 (
            .O(N__54821),
            .I(N__54770));
    InMux I__9544 (
            .O(N__54818),
            .I(N__54762));
    InMux I__9543 (
            .O(N__54815),
            .I(N__54762));
    InMux I__9542 (
            .O(N__54812),
            .I(N__54762));
    InMux I__9541 (
            .O(N__54809),
            .I(N__54753));
    InMux I__9540 (
            .O(N__54806),
            .I(N__54753));
    InMux I__9539 (
            .O(N__54803),
            .I(N__54753));
    InMux I__9538 (
            .O(N__54800),
            .I(N__54753));
    InMux I__9537 (
            .O(N__54797),
            .I(N__54744));
    InMux I__9536 (
            .O(N__54794),
            .I(N__54744));
    InMux I__9535 (
            .O(N__54791),
            .I(N__54744));
    InMux I__9534 (
            .O(N__54788),
            .I(N__54744));
    InMux I__9533 (
            .O(N__54785),
            .I(N__54735));
    InMux I__9532 (
            .O(N__54782),
            .I(N__54735));
    InMux I__9531 (
            .O(N__54779),
            .I(N__54735));
    InMux I__9530 (
            .O(N__54776),
            .I(N__54735));
    InMux I__9529 (
            .O(N__54773),
            .I(N__54730));
    InMux I__9528 (
            .O(N__54770),
            .I(N__54730));
    InMux I__9527 (
            .O(N__54769),
            .I(N__54727));
    LocalMux I__9526 (
            .O(N__54762),
            .I(\quad_counter0.n3431 ));
    LocalMux I__9525 (
            .O(N__54753),
            .I(\quad_counter0.n3431 ));
    LocalMux I__9524 (
            .O(N__54744),
            .I(\quad_counter0.n3431 ));
    LocalMux I__9523 (
            .O(N__54735),
            .I(\quad_counter0.n3431 ));
    LocalMux I__9522 (
            .O(N__54730),
            .I(\quad_counter0.n3431 ));
    LocalMux I__9521 (
            .O(N__54727),
            .I(\quad_counter0.n3431 ));
    InMux I__9520 (
            .O(N__54714),
            .I(\quad_counter0.n30446 ));
    CascadeMux I__9519 (
            .O(N__54711),
            .I(N__54708));
    InMux I__9518 (
            .O(N__54708),
            .I(N__54705));
    LocalMux I__9517 (
            .O(N__54705),
            .I(N__54702));
    Odrv4 I__9516 (
            .O(N__54702),
            .I(\quad_counter0.n3497 ));
    CascadeMux I__9515 (
            .O(N__54699),
            .I(N__54691));
    CascadeMux I__9514 (
            .O(N__54698),
            .I(N__54688));
    CascadeMux I__9513 (
            .O(N__54697),
            .I(N__54685));
    CascadeMux I__9512 (
            .O(N__54696),
            .I(N__54682));
    CascadeMux I__9511 (
            .O(N__54695),
            .I(N__54679));
    CascadeMux I__9510 (
            .O(N__54694),
            .I(N__54676));
    InMux I__9509 (
            .O(N__54691),
            .I(N__54671));
    InMux I__9508 (
            .O(N__54688),
            .I(N__54671));
    InMux I__9507 (
            .O(N__54685),
            .I(N__54662));
    InMux I__9506 (
            .O(N__54682),
            .I(N__54662));
    InMux I__9505 (
            .O(N__54679),
            .I(N__54662));
    InMux I__9504 (
            .O(N__54676),
            .I(N__54662));
    LocalMux I__9503 (
            .O(N__54671),
            .I(\quad_counter0.n36150 ));
    LocalMux I__9502 (
            .O(N__54662),
            .I(\quad_counter0.n36150 ));
    CascadeMux I__9501 (
            .O(N__54657),
            .I(N__54645));
    CascadeMux I__9500 (
            .O(N__54656),
            .I(N__54642));
    CascadeMux I__9499 (
            .O(N__54655),
            .I(N__54639));
    CascadeMux I__9498 (
            .O(N__54654),
            .I(N__54636));
    CascadeMux I__9497 (
            .O(N__54653),
            .I(N__54633));
    CascadeMux I__9496 (
            .O(N__54652),
            .I(N__54630));
    CascadeMux I__9495 (
            .O(N__54651),
            .I(N__54627));
    CascadeMux I__9494 (
            .O(N__54650),
            .I(N__54624));
    CascadeMux I__9493 (
            .O(N__54649),
            .I(N__54621));
    CascadeMux I__9492 (
            .O(N__54648),
            .I(N__54618));
    InMux I__9491 (
            .O(N__54645),
            .I(N__54611));
    InMux I__9490 (
            .O(N__54642),
            .I(N__54611));
    InMux I__9489 (
            .O(N__54639),
            .I(N__54611));
    InMux I__9488 (
            .O(N__54636),
            .I(N__54602));
    InMux I__9487 (
            .O(N__54633),
            .I(N__54602));
    InMux I__9486 (
            .O(N__54630),
            .I(N__54602));
    InMux I__9485 (
            .O(N__54627),
            .I(N__54602));
    InMux I__9484 (
            .O(N__54624),
            .I(N__54597));
    InMux I__9483 (
            .O(N__54621),
            .I(N__54597));
    InMux I__9482 (
            .O(N__54618),
            .I(N__54594));
    LocalMux I__9481 (
            .O(N__54611),
            .I(\quad_counter0.n2639 ));
    LocalMux I__9480 (
            .O(N__54602),
            .I(\quad_counter0.n2639 ));
    LocalMux I__9479 (
            .O(N__54597),
            .I(\quad_counter0.n2639 ));
    LocalMux I__9478 (
            .O(N__54594),
            .I(\quad_counter0.n2639 ));
    InMux I__9477 (
            .O(N__54585),
            .I(N__54582));
    LocalMux I__9476 (
            .O(N__54582),
            .I(\quad_counter0.n3511 ));
    InMux I__9475 (
            .O(N__54579),
            .I(bfn_15_10_0_));
    InMux I__9474 (
            .O(N__54576),
            .I(N__54571));
    InMux I__9473 (
            .O(N__54575),
            .I(N__54568));
    CascadeMux I__9472 (
            .O(N__54574),
            .I(N__54565));
    LocalMux I__9471 (
            .O(N__54571),
            .I(N__54560));
    LocalMux I__9470 (
            .O(N__54568),
            .I(N__54560));
    InMux I__9469 (
            .O(N__54565),
            .I(N__54557));
    Odrv12 I__9468 (
            .O(N__54560),
            .I(\quad_counter0.n3411 ));
    LocalMux I__9467 (
            .O(N__54557),
            .I(\quad_counter0.n3411 ));
    InMux I__9466 (
            .O(N__54552),
            .I(N__54549));
    LocalMux I__9465 (
            .O(N__54549),
            .I(\quad_counter0.n3510 ));
    InMux I__9464 (
            .O(N__54546),
            .I(\quad_counter0.n30433 ));
    InMux I__9463 (
            .O(N__54543),
            .I(N__54538));
    InMux I__9462 (
            .O(N__54542),
            .I(N__54535));
    CascadeMux I__9461 (
            .O(N__54541),
            .I(N__54532));
    LocalMux I__9460 (
            .O(N__54538),
            .I(N__54527));
    LocalMux I__9459 (
            .O(N__54535),
            .I(N__54527));
    InMux I__9458 (
            .O(N__54532),
            .I(N__54524));
    Odrv12 I__9457 (
            .O(N__54527),
            .I(\quad_counter0.n3410 ));
    LocalMux I__9456 (
            .O(N__54524),
            .I(\quad_counter0.n3410 ));
    InMux I__9455 (
            .O(N__54519),
            .I(N__54516));
    LocalMux I__9454 (
            .O(N__54516),
            .I(\quad_counter0.n3509 ));
    InMux I__9453 (
            .O(N__54513),
            .I(\quad_counter0.n30434 ));
    InMux I__9452 (
            .O(N__54510),
            .I(N__54505));
    InMux I__9451 (
            .O(N__54509),
            .I(N__54502));
    CascadeMux I__9450 (
            .O(N__54508),
            .I(N__54499));
    LocalMux I__9449 (
            .O(N__54505),
            .I(N__54494));
    LocalMux I__9448 (
            .O(N__54502),
            .I(N__54494));
    InMux I__9447 (
            .O(N__54499),
            .I(N__54491));
    Odrv4 I__9446 (
            .O(N__54494),
            .I(\quad_counter0.n3409 ));
    LocalMux I__9445 (
            .O(N__54491),
            .I(\quad_counter0.n3409 ));
    InMux I__9444 (
            .O(N__54486),
            .I(\quad_counter0.n30435 ));
    InMux I__9443 (
            .O(N__54483),
            .I(N__54479));
    InMux I__9442 (
            .O(N__54482),
            .I(N__54476));
    LocalMux I__9441 (
            .O(N__54479),
            .I(N__54470));
    LocalMux I__9440 (
            .O(N__54476),
            .I(N__54470));
    InMux I__9439 (
            .O(N__54475),
            .I(N__54467));
    Odrv4 I__9438 (
            .O(N__54470),
            .I(\quad_counter0.n3408 ));
    LocalMux I__9437 (
            .O(N__54467),
            .I(\quad_counter0.n3408 ));
    InMux I__9436 (
            .O(N__54462),
            .I(\quad_counter0.n30436 ));
    InMux I__9435 (
            .O(N__54459),
            .I(N__54455));
    InMux I__9434 (
            .O(N__54458),
            .I(N__54452));
    LocalMux I__9433 (
            .O(N__54455),
            .I(N__54446));
    LocalMux I__9432 (
            .O(N__54452),
            .I(N__54446));
    InMux I__9431 (
            .O(N__54451),
            .I(N__54443));
    Odrv4 I__9430 (
            .O(N__54446),
            .I(\quad_counter0.n3407 ));
    LocalMux I__9429 (
            .O(N__54443),
            .I(\quad_counter0.n3407 ));
    InMux I__9428 (
            .O(N__54438),
            .I(N__54435));
    LocalMux I__9427 (
            .O(N__54435),
            .I(\quad_counter0.n3506 ));
    InMux I__9426 (
            .O(N__54432),
            .I(\quad_counter0.n30437 ));
    InMux I__9425 (
            .O(N__54429),
            .I(N__54425));
    InMux I__9424 (
            .O(N__54428),
            .I(N__54422));
    LocalMux I__9423 (
            .O(N__54425),
            .I(N__54416));
    LocalMux I__9422 (
            .O(N__54422),
            .I(N__54416));
    InMux I__9421 (
            .O(N__54421),
            .I(N__54413));
    Odrv4 I__9420 (
            .O(N__54416),
            .I(\quad_counter0.n3406 ));
    LocalMux I__9419 (
            .O(N__54413),
            .I(\quad_counter0.n3406 ));
    InMux I__9418 (
            .O(N__54408),
            .I(N__54405));
    LocalMux I__9417 (
            .O(N__54405),
            .I(\quad_counter0.n3505 ));
    InMux I__9416 (
            .O(N__54402),
            .I(\quad_counter0.n30438 ));
    InMux I__9415 (
            .O(N__54399),
            .I(N__54395));
    InMux I__9414 (
            .O(N__54398),
            .I(N__54392));
    LocalMux I__9413 (
            .O(N__54395),
            .I(N__54386));
    LocalMux I__9412 (
            .O(N__54392),
            .I(N__54386));
    InMux I__9411 (
            .O(N__54391),
            .I(N__54383));
    Odrv12 I__9410 (
            .O(N__54386),
            .I(\quad_counter0.n3405 ));
    LocalMux I__9409 (
            .O(N__54383),
            .I(\quad_counter0.n3405 ));
    InMux I__9408 (
            .O(N__54378),
            .I(\quad_counter0.n30439 ));
    InMux I__9407 (
            .O(N__54375),
            .I(N__54371));
    InMux I__9406 (
            .O(N__54374),
            .I(N__54368));
    LocalMux I__9405 (
            .O(N__54371),
            .I(N__54363));
    LocalMux I__9404 (
            .O(N__54368),
            .I(N__54363));
    Span4Mux_h I__9403 (
            .O(N__54363),
            .I(N__54359));
    InMux I__9402 (
            .O(N__54362),
            .I(N__54356));
    Odrv4 I__9401 (
            .O(N__54359),
            .I(\quad_counter0.n3404 ));
    LocalMux I__9400 (
            .O(N__54356),
            .I(\quad_counter0.n3404 ));
    InMux I__9399 (
            .O(N__54351),
            .I(bfn_15_9_0_));
    InMux I__9398 (
            .O(N__54348),
            .I(N__54343));
    InMux I__9397 (
            .O(N__54347),
            .I(N__54340));
    CascadeMux I__9396 (
            .O(N__54346),
            .I(N__54337));
    LocalMux I__9395 (
            .O(N__54343),
            .I(N__54332));
    LocalMux I__9394 (
            .O(N__54340),
            .I(N__54332));
    InMux I__9393 (
            .O(N__54337),
            .I(N__54329));
    Odrv12 I__9392 (
            .O(N__54332),
            .I(\quad_counter0.n3419 ));
    LocalMux I__9391 (
            .O(N__54329),
            .I(\quad_counter0.n3419 ));
    InMux I__9390 (
            .O(N__54324),
            .I(\quad_counter0.n30425 ));
    InMux I__9389 (
            .O(N__54321),
            .I(N__54317));
    InMux I__9388 (
            .O(N__54320),
            .I(N__54314));
    LocalMux I__9387 (
            .O(N__54317),
            .I(N__54308));
    LocalMux I__9386 (
            .O(N__54314),
            .I(N__54308));
    InMux I__9385 (
            .O(N__54313),
            .I(N__54305));
    Odrv12 I__9384 (
            .O(N__54308),
            .I(\quad_counter0.n3418 ));
    LocalMux I__9383 (
            .O(N__54305),
            .I(\quad_counter0.n3418 ));
    InMux I__9382 (
            .O(N__54300),
            .I(\quad_counter0.n30426 ));
    InMux I__9381 (
            .O(N__54297),
            .I(N__54292));
    InMux I__9380 (
            .O(N__54296),
            .I(N__54289));
    CascadeMux I__9379 (
            .O(N__54295),
            .I(N__54286));
    LocalMux I__9378 (
            .O(N__54292),
            .I(N__54281));
    LocalMux I__9377 (
            .O(N__54289),
            .I(N__54281));
    InMux I__9376 (
            .O(N__54286),
            .I(N__54278));
    Odrv4 I__9375 (
            .O(N__54281),
            .I(\quad_counter0.n3417 ));
    LocalMux I__9374 (
            .O(N__54278),
            .I(\quad_counter0.n3417 ));
    InMux I__9373 (
            .O(N__54273),
            .I(\quad_counter0.n30427 ));
    InMux I__9372 (
            .O(N__54270),
            .I(N__54266));
    InMux I__9371 (
            .O(N__54269),
            .I(N__54263));
    LocalMux I__9370 (
            .O(N__54266),
            .I(N__54257));
    LocalMux I__9369 (
            .O(N__54263),
            .I(N__54257));
    InMux I__9368 (
            .O(N__54262),
            .I(N__54254));
    Odrv4 I__9367 (
            .O(N__54257),
            .I(\quad_counter0.n3416 ));
    LocalMux I__9366 (
            .O(N__54254),
            .I(\quad_counter0.n3416 ));
    InMux I__9365 (
            .O(N__54249),
            .I(\quad_counter0.n30428 ));
    InMux I__9364 (
            .O(N__54246),
            .I(N__54242));
    InMux I__9363 (
            .O(N__54245),
            .I(N__54239));
    LocalMux I__9362 (
            .O(N__54242),
            .I(N__54233));
    LocalMux I__9361 (
            .O(N__54239),
            .I(N__54233));
    InMux I__9360 (
            .O(N__54238),
            .I(N__54230));
    Odrv4 I__9359 (
            .O(N__54233),
            .I(\quad_counter0.n3415 ));
    LocalMux I__9358 (
            .O(N__54230),
            .I(\quad_counter0.n3415 ));
    InMux I__9357 (
            .O(N__54225),
            .I(\quad_counter0.n30429 ));
    InMux I__9356 (
            .O(N__54222),
            .I(N__54218));
    InMux I__9355 (
            .O(N__54221),
            .I(N__54215));
    LocalMux I__9354 (
            .O(N__54218),
            .I(N__54209));
    LocalMux I__9353 (
            .O(N__54215),
            .I(N__54209));
    InMux I__9352 (
            .O(N__54214),
            .I(N__54206));
    Odrv4 I__9351 (
            .O(N__54209),
            .I(\quad_counter0.n3414 ));
    LocalMux I__9350 (
            .O(N__54206),
            .I(\quad_counter0.n3414 ));
    CascadeMux I__9349 (
            .O(N__54201),
            .I(N__54193));
    CascadeMux I__9348 (
            .O(N__54200),
            .I(N__54190));
    CascadeMux I__9347 (
            .O(N__54199),
            .I(N__54187));
    CascadeMux I__9346 (
            .O(N__54198),
            .I(N__54184));
    CascadeMux I__9345 (
            .O(N__54197),
            .I(N__54181));
    CascadeMux I__9344 (
            .O(N__54196),
            .I(N__54178));
    InMux I__9343 (
            .O(N__54193),
            .I(N__54173));
    InMux I__9342 (
            .O(N__54190),
            .I(N__54173));
    InMux I__9341 (
            .O(N__54187),
            .I(N__54164));
    InMux I__9340 (
            .O(N__54184),
            .I(N__54164));
    InMux I__9339 (
            .O(N__54181),
            .I(N__54164));
    InMux I__9338 (
            .O(N__54178),
            .I(N__54164));
    LocalMux I__9337 (
            .O(N__54173),
            .I(\quad_counter0.n36139 ));
    LocalMux I__9336 (
            .O(N__54164),
            .I(\quad_counter0.n36139 ));
    InMux I__9335 (
            .O(N__54159),
            .I(\quad_counter0.n30430 ));
    InMux I__9334 (
            .O(N__54156),
            .I(N__54152));
    InMux I__9333 (
            .O(N__54155),
            .I(N__54149));
    LocalMux I__9332 (
            .O(N__54152),
            .I(N__54143));
    LocalMux I__9331 (
            .O(N__54149),
            .I(N__54143));
    InMux I__9330 (
            .O(N__54148),
            .I(N__54140));
    Odrv12 I__9329 (
            .O(N__54143),
            .I(\quad_counter0.n3413 ));
    LocalMux I__9328 (
            .O(N__54140),
            .I(\quad_counter0.n3413 ));
    InMux I__9327 (
            .O(N__54135),
            .I(\quad_counter0.n30431 ));
    InMux I__9326 (
            .O(N__54132),
            .I(N__54128));
    InMux I__9325 (
            .O(N__54131),
            .I(N__54125));
    LocalMux I__9324 (
            .O(N__54128),
            .I(N__54120));
    LocalMux I__9323 (
            .O(N__54125),
            .I(N__54120));
    Span4Mux_h I__9322 (
            .O(N__54120),
            .I(N__54116));
    InMux I__9321 (
            .O(N__54119),
            .I(N__54113));
    Odrv4 I__9320 (
            .O(N__54116),
            .I(\quad_counter0.n3412 ));
    LocalMux I__9319 (
            .O(N__54113),
            .I(\quad_counter0.n3412 ));
    InMux I__9318 (
            .O(N__54108),
            .I(N__54105));
    LocalMux I__9317 (
            .O(N__54105),
            .I(\quad_counter0.n2081 ));
    CascadeMux I__9316 (
            .O(N__54102),
            .I(N__54099));
    InMux I__9315 (
            .O(N__54099),
            .I(N__54095));
    InMux I__9314 (
            .O(N__54098),
            .I(N__54092));
    LocalMux I__9313 (
            .O(N__54095),
            .I(N__54089));
    LocalMux I__9312 (
            .O(N__54092),
            .I(\quad_counter0.n2014 ));
    Odrv4 I__9311 (
            .O(N__54089),
            .I(\quad_counter0.n2014 ));
    CascadeMux I__9310 (
            .O(N__54084),
            .I(N__54081));
    InMux I__9309 (
            .O(N__54081),
            .I(N__54077));
    CascadeMux I__9308 (
            .O(N__54080),
            .I(N__54074));
    LocalMux I__9307 (
            .O(N__54077),
            .I(N__54070));
    InMux I__9306 (
            .O(N__54074),
            .I(N__54067));
    InMux I__9305 (
            .O(N__54073),
            .I(N__54064));
    Odrv4 I__9304 (
            .O(N__54070),
            .I(\quad_counter0.n2015 ));
    LocalMux I__9303 (
            .O(N__54067),
            .I(\quad_counter0.n2015 ));
    LocalMux I__9302 (
            .O(N__54064),
            .I(\quad_counter0.n2015 ));
    InMux I__9301 (
            .O(N__54057),
            .I(N__54054));
    LocalMux I__9300 (
            .O(N__54054),
            .I(\quad_counter0.n2082 ));
    InMux I__9299 (
            .O(N__54051),
            .I(N__54048));
    LocalMux I__9298 (
            .O(N__54048),
            .I(N__54045));
    Span4Mux_v I__9297 (
            .O(N__54045),
            .I(N__54040));
    InMux I__9296 (
            .O(N__54044),
            .I(N__54037));
    InMux I__9295 (
            .O(N__54043),
            .I(N__54034));
    Odrv4 I__9294 (
            .O(N__54040),
            .I(\quad_counter0.n1919 ));
    LocalMux I__9293 (
            .O(N__54037),
            .I(\quad_counter0.n1919 ));
    LocalMux I__9292 (
            .O(N__54034),
            .I(\quad_counter0.n1919 ));
    CascadeMux I__9291 (
            .O(N__54027),
            .I(N__54024));
    InMux I__9290 (
            .O(N__54024),
            .I(N__54021));
    LocalMux I__9289 (
            .O(N__54021),
            .I(N__54018));
    Span4Mux_v I__9288 (
            .O(N__54018),
            .I(N__54015));
    Odrv4 I__9287 (
            .O(N__54015),
            .I(\quad_counter0.n1986 ));
    CascadeMux I__9286 (
            .O(N__54012),
            .I(N__54006));
    InMux I__9285 (
            .O(N__54011),
            .I(N__54002));
    InMux I__9284 (
            .O(N__54010),
            .I(N__53999));
    CascadeMux I__9283 (
            .O(N__54009),
            .I(N__53995));
    InMux I__9282 (
            .O(N__54006),
            .I(N__53991));
    InMux I__9281 (
            .O(N__54005),
            .I(N__53988));
    LocalMux I__9280 (
            .O(N__54002),
            .I(N__53983));
    LocalMux I__9279 (
            .O(N__53999),
            .I(N__53983));
    InMux I__9278 (
            .O(N__53998),
            .I(N__53976));
    InMux I__9277 (
            .O(N__53995),
            .I(N__53976));
    InMux I__9276 (
            .O(N__53994),
            .I(N__53976));
    LocalMux I__9275 (
            .O(N__53991),
            .I(\quad_counter0.n1946 ));
    LocalMux I__9274 (
            .O(N__53988),
            .I(\quad_counter0.n1946 ));
    Odrv4 I__9273 (
            .O(N__53983),
            .I(\quad_counter0.n1946 ));
    LocalMux I__9272 (
            .O(N__53976),
            .I(\quad_counter0.n1946 ));
    CascadeMux I__9271 (
            .O(N__53967),
            .I(N__53963));
    InMux I__9270 (
            .O(N__53966),
            .I(N__53960));
    InMux I__9269 (
            .O(N__53963),
            .I(N__53957));
    LocalMux I__9268 (
            .O(N__53960),
            .I(\quad_counter0.n2018 ));
    LocalMux I__9267 (
            .O(N__53957),
            .I(\quad_counter0.n2018 ));
    InMux I__9266 (
            .O(N__53952),
            .I(N__53949));
    LocalMux I__9265 (
            .O(N__53949),
            .I(\quad_counter0.n2085 ));
    CascadeMux I__9264 (
            .O(N__53946),
            .I(\quad_counter0.n2018_cascade_ ));
    InMux I__9263 (
            .O(N__53943),
            .I(N__53938));
    CascadeMux I__9262 (
            .O(N__53942),
            .I(N__53935));
    CascadeMux I__9261 (
            .O(N__53941),
            .I(N__53932));
    LocalMux I__9260 (
            .O(N__53938),
            .I(N__53929));
    InMux I__9259 (
            .O(N__53935),
            .I(N__53926));
    InMux I__9258 (
            .O(N__53932),
            .I(N__53923));
    Odrv12 I__9257 (
            .O(N__53929),
            .I(\quad_counter0.n2016 ));
    LocalMux I__9256 (
            .O(N__53926),
            .I(\quad_counter0.n2016 ));
    LocalMux I__9255 (
            .O(N__53923),
            .I(\quad_counter0.n2016 ));
    CascadeMux I__9254 (
            .O(N__53916),
            .I(N__53913));
    InMux I__9253 (
            .O(N__53913),
            .I(N__53910));
    LocalMux I__9252 (
            .O(N__53910),
            .I(\quad_counter0.n2083 ));
    CascadeMux I__9251 (
            .O(N__53907),
            .I(N__53901));
    CascadeMux I__9250 (
            .O(N__53906),
            .I(N__53897));
    CascadeMux I__9249 (
            .O(N__53905),
            .I(N__53893));
    InMux I__9248 (
            .O(N__53904),
            .I(N__53888));
    InMux I__9247 (
            .O(N__53901),
            .I(N__53883));
    InMux I__9246 (
            .O(N__53900),
            .I(N__53883));
    InMux I__9245 (
            .O(N__53897),
            .I(N__53872));
    InMux I__9244 (
            .O(N__53896),
            .I(N__53872));
    InMux I__9243 (
            .O(N__53893),
            .I(N__53872));
    InMux I__9242 (
            .O(N__53892),
            .I(N__53872));
    InMux I__9241 (
            .O(N__53891),
            .I(N__53872));
    LocalMux I__9240 (
            .O(N__53888),
            .I(\quad_counter0.n2045 ));
    LocalMux I__9239 (
            .O(N__53883),
            .I(\quad_counter0.n2045 ));
    LocalMux I__9238 (
            .O(N__53872),
            .I(\quad_counter0.n2045 ));
    CascadeMux I__9237 (
            .O(N__53865),
            .I(\quad_counter0.n8_adj_4380_cascade_ ));
    InMux I__9236 (
            .O(N__53862),
            .I(N__53859));
    LocalMux I__9235 (
            .O(N__53859),
            .I(\quad_counter0.n7_adj_4381 ));
    CascadeMux I__9234 (
            .O(N__53856),
            .I(\quad_counter0.n35542_cascade_ ));
    InMux I__9233 (
            .O(N__53853),
            .I(N__53850));
    LocalMux I__9232 (
            .O(N__53850),
            .I(N__53847));
    Span4Mux_h I__9231 (
            .O(N__53847),
            .I(N__53843));
    InMux I__9230 (
            .O(N__53846),
            .I(N__53840));
    Odrv4 I__9229 (
            .O(N__53843),
            .I(\c0.n33653 ));
    LocalMux I__9228 (
            .O(N__53840),
            .I(\c0.n33653 ));
    CascadeMux I__9227 (
            .O(N__53835),
            .I(\c0.n15_adj_4664_cascade_ ));
    InMux I__9226 (
            .O(N__53832),
            .I(N__53829));
    LocalMux I__9225 (
            .O(N__53829),
            .I(\c0.n14_adj_4663 ));
    InMux I__9224 (
            .O(N__53826),
            .I(N__53820));
    InMux I__9223 (
            .O(N__53825),
            .I(N__53820));
    LocalMux I__9222 (
            .O(N__53820),
            .I(\c0.n33939 ));
    InMux I__9221 (
            .O(N__53817),
            .I(N__53814));
    LocalMux I__9220 (
            .O(N__53814),
            .I(N__53809));
    InMux I__9219 (
            .O(N__53813),
            .I(N__53804));
    InMux I__9218 (
            .O(N__53812),
            .I(N__53804));
    Span4Mux_v I__9217 (
            .O(N__53809),
            .I(N__53798));
    LocalMux I__9216 (
            .O(N__53804),
            .I(N__53798));
    InMux I__9215 (
            .O(N__53803),
            .I(N__53795));
    Span4Mux_v I__9214 (
            .O(N__53798),
            .I(N__53792));
    LocalMux I__9213 (
            .O(N__53795),
            .I(\c0.data_in_frame_20_7 ));
    Odrv4 I__9212 (
            .O(N__53792),
            .I(\c0.data_in_frame_20_7 ));
    CascadeMux I__9211 (
            .O(N__53787),
            .I(N__53784));
    InMux I__9210 (
            .O(N__53784),
            .I(N__53779));
    InMux I__9209 (
            .O(N__53783),
            .I(N__53774));
    InMux I__9208 (
            .O(N__53782),
            .I(N__53774));
    LocalMux I__9207 (
            .O(N__53779),
            .I(\c0.data_in_frame_20_6 ));
    LocalMux I__9206 (
            .O(N__53774),
            .I(\c0.data_in_frame_20_6 ));
    CascadeMux I__9205 (
            .O(N__53769),
            .I(N__53766));
    InMux I__9204 (
            .O(N__53766),
            .I(N__53758));
    InMux I__9203 (
            .O(N__53765),
            .I(N__53758));
    CascadeMux I__9202 (
            .O(N__53764),
            .I(N__53755));
    CascadeMux I__9201 (
            .O(N__53763),
            .I(N__53752));
    LocalMux I__9200 (
            .O(N__53758),
            .I(N__53749));
    InMux I__9199 (
            .O(N__53755),
            .I(N__53744));
    InMux I__9198 (
            .O(N__53752),
            .I(N__53744));
    Odrv4 I__9197 (
            .O(N__53749),
            .I(\c0.data_in_frame_23_2 ));
    LocalMux I__9196 (
            .O(N__53744),
            .I(\c0.data_in_frame_23_2 ));
    InMux I__9195 (
            .O(N__53739),
            .I(N__53733));
    InMux I__9194 (
            .O(N__53738),
            .I(N__53733));
    LocalMux I__9193 (
            .O(N__53733),
            .I(\c0.n18559 ));
    CascadeMux I__9192 (
            .O(N__53730),
            .I(\c0.n6404_cascade_ ));
    InMux I__9191 (
            .O(N__53727),
            .I(N__53723));
    InMux I__9190 (
            .O(N__53726),
            .I(N__53720));
    LocalMux I__9189 (
            .O(N__53723),
            .I(\c0.n32390 ));
    LocalMux I__9188 (
            .O(N__53720),
            .I(\c0.n32390 ));
    InMux I__9187 (
            .O(N__53715),
            .I(N__53711));
    CascadeMux I__9186 (
            .O(N__53714),
            .I(N__53707));
    LocalMux I__9185 (
            .O(N__53711),
            .I(N__53703));
    InMux I__9184 (
            .O(N__53710),
            .I(N__53700));
    InMux I__9183 (
            .O(N__53707),
            .I(N__53697));
    InMux I__9182 (
            .O(N__53706),
            .I(N__53694));
    Span4Mux_h I__9181 (
            .O(N__53703),
            .I(N__53691));
    LocalMux I__9180 (
            .O(N__53700),
            .I(N__53688));
    LocalMux I__9179 (
            .O(N__53697),
            .I(\c0.data_in_frame_16_6 ));
    LocalMux I__9178 (
            .O(N__53694),
            .I(\c0.data_in_frame_16_6 ));
    Odrv4 I__9177 (
            .O(N__53691),
            .I(\c0.data_in_frame_16_6 ));
    Odrv12 I__9176 (
            .O(N__53688),
            .I(\c0.data_in_frame_16_6 ));
    CascadeMux I__9175 (
            .O(N__53679),
            .I(N__53674));
    InMux I__9174 (
            .O(N__53678),
            .I(N__53671));
    InMux I__9173 (
            .O(N__53677),
            .I(N__53668));
    InMux I__9172 (
            .O(N__53674),
            .I(N__53665));
    LocalMux I__9171 (
            .O(N__53671),
            .I(\quad_counter0.n2017 ));
    LocalMux I__9170 (
            .O(N__53668),
            .I(\quad_counter0.n2017 ));
    LocalMux I__9169 (
            .O(N__53665),
            .I(\quad_counter0.n2017 ));
    InMux I__9168 (
            .O(N__53658),
            .I(N__53655));
    LocalMux I__9167 (
            .O(N__53655),
            .I(\quad_counter0.n2084 ));
    CascadeMux I__9166 (
            .O(N__53652),
            .I(\c0.n18578_cascade_ ));
    CascadeMux I__9165 (
            .O(N__53649),
            .I(\c0.n15_adj_4746_cascade_ ));
    InMux I__9164 (
            .O(N__53646),
            .I(N__53643));
    LocalMux I__9163 (
            .O(N__53643),
            .I(\c0.n14_adj_4578 ));
    CascadeMux I__9162 (
            .O(N__53640),
            .I(\c0.n32087_cascade_ ));
    InMux I__9161 (
            .O(N__53637),
            .I(N__53633));
    InMux I__9160 (
            .O(N__53636),
            .I(N__53630));
    LocalMux I__9159 (
            .O(N__53633),
            .I(\c0.data_in_frame_26_5 ));
    LocalMux I__9158 (
            .O(N__53630),
            .I(\c0.data_in_frame_26_5 ));
    InMux I__9157 (
            .O(N__53625),
            .I(N__53622));
    LocalMux I__9156 (
            .O(N__53622),
            .I(N__53618));
    InMux I__9155 (
            .O(N__53621),
            .I(N__53615));
    Span4Mux_h I__9154 (
            .O(N__53618),
            .I(N__53612));
    LocalMux I__9153 (
            .O(N__53615),
            .I(\c0.n33966 ));
    Odrv4 I__9152 (
            .O(N__53612),
            .I(\c0.n33966 ));
    InMux I__9151 (
            .O(N__53607),
            .I(N__53602));
    CascadeMux I__9150 (
            .O(N__53606),
            .I(N__53599));
    InMux I__9149 (
            .O(N__53605),
            .I(N__53596));
    LocalMux I__9148 (
            .O(N__53602),
            .I(N__53591));
    InMux I__9147 (
            .O(N__53599),
            .I(N__53588));
    LocalMux I__9146 (
            .O(N__53596),
            .I(N__53585));
    InMux I__9145 (
            .O(N__53595),
            .I(N__53580));
    InMux I__9144 (
            .O(N__53594),
            .I(N__53580));
    Span4Mux_v I__9143 (
            .O(N__53591),
            .I(N__53577));
    LocalMux I__9142 (
            .O(N__53588),
            .I(\c0.data_in_frame_16_3 ));
    Odrv4 I__9141 (
            .O(N__53585),
            .I(\c0.data_in_frame_16_3 ));
    LocalMux I__9140 (
            .O(N__53580),
            .I(\c0.data_in_frame_16_3 ));
    Odrv4 I__9139 (
            .O(N__53577),
            .I(\c0.data_in_frame_16_3 ));
    InMux I__9138 (
            .O(N__53568),
            .I(N__53565));
    LocalMux I__9137 (
            .O(N__53565),
            .I(N__53562));
    Span4Mux_v I__9136 (
            .O(N__53562),
            .I(N__53558));
    InMux I__9135 (
            .O(N__53561),
            .I(N__53555));
    Odrv4 I__9134 (
            .O(N__53558),
            .I(\c0.n33526 ));
    LocalMux I__9133 (
            .O(N__53555),
            .I(\c0.n33526 ));
    InMux I__9132 (
            .O(N__53550),
            .I(N__53545));
    CascadeMux I__9131 (
            .O(N__53549),
            .I(N__53542));
    InMux I__9130 (
            .O(N__53548),
            .I(N__53539));
    LocalMux I__9129 (
            .O(N__53545),
            .I(N__53536));
    InMux I__9128 (
            .O(N__53542),
            .I(N__53532));
    LocalMux I__9127 (
            .O(N__53539),
            .I(N__53527));
    Span4Mux_v I__9126 (
            .O(N__53536),
            .I(N__53527));
    InMux I__9125 (
            .O(N__53535),
            .I(N__53524));
    LocalMux I__9124 (
            .O(N__53532),
            .I(N__53519));
    Span4Mux_v I__9123 (
            .O(N__53527),
            .I(N__53519));
    LocalMux I__9122 (
            .O(N__53524),
            .I(\c0.data_in_frame_18_5 ));
    Odrv4 I__9121 (
            .O(N__53519),
            .I(\c0.data_in_frame_18_5 ));
    InMux I__9120 (
            .O(N__53514),
            .I(N__53511));
    LocalMux I__9119 (
            .O(N__53511),
            .I(N__53507));
    InMux I__9118 (
            .O(N__53510),
            .I(N__53504));
    Span4Mux_h I__9117 (
            .O(N__53507),
            .I(N__53498));
    LocalMux I__9116 (
            .O(N__53504),
            .I(N__53498));
    InMux I__9115 (
            .O(N__53503),
            .I(N__53495));
    Span4Mux_v I__9114 (
            .O(N__53498),
            .I(N__53489));
    LocalMux I__9113 (
            .O(N__53495),
            .I(N__53489));
    InMux I__9112 (
            .O(N__53494),
            .I(N__53486));
    Span4Mux_h I__9111 (
            .O(N__53489),
            .I(N__53483));
    LocalMux I__9110 (
            .O(N__53486),
            .I(N__53480));
    Odrv4 I__9109 (
            .O(N__53483),
            .I(\c0.n31651 ));
    Odrv12 I__9108 (
            .O(N__53480),
            .I(\c0.n31651 ));
    CascadeMux I__9107 (
            .O(N__53475),
            .I(\c0.n18559_cascade_ ));
    InMux I__9106 (
            .O(N__53472),
            .I(N__53467));
    InMux I__9105 (
            .O(N__53471),
            .I(N__53462));
    InMux I__9104 (
            .O(N__53470),
            .I(N__53462));
    LocalMux I__9103 (
            .O(N__53467),
            .I(N__53459));
    LocalMux I__9102 (
            .O(N__53462),
            .I(N__53456));
    Span4Mux_v I__9101 (
            .O(N__53459),
            .I(N__53452));
    Span4Mux_h I__9100 (
            .O(N__53456),
            .I(N__53449));
    InMux I__9099 (
            .O(N__53455),
            .I(N__53446));
    Odrv4 I__9098 (
            .O(N__53452),
            .I(\c0.n33972 ));
    Odrv4 I__9097 (
            .O(N__53449),
            .I(\c0.n33972 ));
    LocalMux I__9096 (
            .O(N__53446),
            .I(\c0.n33972 ));
    CascadeMux I__9095 (
            .O(N__53439),
            .I(\c0.n6023_cascade_ ));
    InMux I__9094 (
            .O(N__53436),
            .I(N__53433));
    LocalMux I__9093 (
            .O(N__53433),
            .I(N__53427));
    InMux I__9092 (
            .O(N__53432),
            .I(N__53424));
    InMux I__9091 (
            .O(N__53431),
            .I(N__53419));
    InMux I__9090 (
            .O(N__53430),
            .I(N__53419));
    Span4Mux_v I__9089 (
            .O(N__53427),
            .I(N__53416));
    LocalMux I__9088 (
            .O(N__53424),
            .I(N__53413));
    LocalMux I__9087 (
            .O(N__53419),
            .I(\c0.data_in_frame_17_0 ));
    Odrv4 I__9086 (
            .O(N__53416),
            .I(\c0.data_in_frame_17_0 ));
    Odrv4 I__9085 (
            .O(N__53413),
            .I(\c0.data_in_frame_17_0 ));
    InMux I__9084 (
            .O(N__53406),
            .I(N__53401));
    InMux I__9083 (
            .O(N__53405),
            .I(N__53396));
    InMux I__9082 (
            .O(N__53404),
            .I(N__53396));
    LocalMux I__9081 (
            .O(N__53401),
            .I(N__53393));
    LocalMux I__9080 (
            .O(N__53396),
            .I(\c0.n33458 ));
    Odrv4 I__9079 (
            .O(N__53393),
            .I(\c0.n33458 ));
    InMux I__9078 (
            .O(N__53388),
            .I(N__53385));
    LocalMux I__9077 (
            .O(N__53385),
            .I(N__53382));
    Odrv4 I__9076 (
            .O(N__53382),
            .I(\c0.n19108 ));
    InMux I__9075 (
            .O(N__53379),
            .I(N__53376));
    LocalMux I__9074 (
            .O(N__53376),
            .I(N__53373));
    Span4Mux_h I__9073 (
            .O(N__53373),
            .I(N__53370));
    Odrv4 I__9072 (
            .O(N__53370),
            .I(\c0.n10_adj_4709 ));
    CascadeMux I__9071 (
            .O(N__53367),
            .I(\c0.n33621_cascade_ ));
    InMux I__9070 (
            .O(N__53364),
            .I(N__53355));
    InMux I__9069 (
            .O(N__53363),
            .I(N__53355));
    CascadeMux I__9068 (
            .O(N__53362),
            .I(N__53352));
    CascadeMux I__9067 (
            .O(N__53361),
            .I(N__53349));
    InMux I__9066 (
            .O(N__53360),
            .I(N__53346));
    LocalMux I__9065 (
            .O(N__53355),
            .I(N__53343));
    InMux I__9064 (
            .O(N__53352),
            .I(N__53340));
    InMux I__9063 (
            .O(N__53349),
            .I(N__53337));
    LocalMux I__9062 (
            .O(N__53346),
            .I(N__53334));
    Span4Mux_h I__9061 (
            .O(N__53343),
            .I(N__53331));
    LocalMux I__9060 (
            .O(N__53340),
            .I(N__53328));
    LocalMux I__9059 (
            .O(N__53337),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__9058 (
            .O(N__53334),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__9057 (
            .O(N__53331),
            .I(\c0.data_in_frame_16_7 ));
    Odrv4 I__9056 (
            .O(N__53328),
            .I(\c0.data_in_frame_16_7 ));
    InMux I__9055 (
            .O(N__53319),
            .I(N__53315));
    CascadeMux I__9054 (
            .O(N__53318),
            .I(N__53312));
    LocalMux I__9053 (
            .O(N__53315),
            .I(N__53308));
    InMux I__9052 (
            .O(N__53312),
            .I(N__53303));
    InMux I__9051 (
            .O(N__53311),
            .I(N__53303));
    Span4Mux_h I__9050 (
            .O(N__53308),
            .I(N__53300));
    LocalMux I__9049 (
            .O(N__53303),
            .I(\c0.data_in_frame_19_3 ));
    Odrv4 I__9048 (
            .O(N__53300),
            .I(\c0.data_in_frame_19_3 ));
    InMux I__9047 (
            .O(N__53295),
            .I(N__53292));
    LocalMux I__9046 (
            .O(N__53292),
            .I(N__53289));
    Odrv4 I__9045 (
            .O(N__53289),
            .I(\c0.n12_adj_4712 ));
    CascadeMux I__9044 (
            .O(N__53286),
            .I(\c0.n8_adj_4711_cascade_ ));
    InMux I__9043 (
            .O(N__53283),
            .I(N__53280));
    LocalMux I__9042 (
            .O(N__53280),
            .I(N__53277));
    Odrv12 I__9041 (
            .O(N__53277),
            .I(\c0.n19060 ));
    InMux I__9040 (
            .O(N__53274),
            .I(N__53268));
    InMux I__9039 (
            .O(N__53273),
            .I(N__53268));
    LocalMux I__9038 (
            .O(N__53268),
            .I(\c0.data_in_frame_28_4 ));
    CascadeMux I__9037 (
            .O(N__53265),
            .I(\c0.n12_adj_4748_cascade_ ));
    InMux I__9036 (
            .O(N__53262),
            .I(N__53259));
    LocalMux I__9035 (
            .O(N__53259),
            .I(\c0.n33517 ));
    CascadeMux I__9034 (
            .O(N__53256),
            .I(\c0.n33517_cascade_ ));
    InMux I__9033 (
            .O(N__53253),
            .I(N__53250));
    LocalMux I__9032 (
            .O(N__53250),
            .I(N__53247));
    Span4Mux_v I__9031 (
            .O(N__53247),
            .I(N__53244));
    Odrv4 I__9030 (
            .O(N__53244),
            .I(\c0.n33441 ));
    InMux I__9029 (
            .O(N__53241),
            .I(N__53238));
    LocalMux I__9028 (
            .O(N__53238),
            .I(N__53234));
    InMux I__9027 (
            .O(N__53237),
            .I(N__53231));
    Odrv12 I__9026 (
            .O(N__53234),
            .I(\c0.n33768 ));
    LocalMux I__9025 (
            .O(N__53231),
            .I(\c0.n33768 ));
    InMux I__9024 (
            .O(N__53226),
            .I(N__53222));
    InMux I__9023 (
            .O(N__53225),
            .I(N__53218));
    LocalMux I__9022 (
            .O(N__53222),
            .I(N__53215));
    CascadeMux I__9021 (
            .O(N__53221),
            .I(N__53212));
    LocalMux I__9020 (
            .O(N__53218),
            .I(N__53208));
    Span4Mux_v I__9019 (
            .O(N__53215),
            .I(N__53204));
    InMux I__9018 (
            .O(N__53212),
            .I(N__53201));
    InMux I__9017 (
            .O(N__53211),
            .I(N__53198));
    Span12Mux_s8_v I__9016 (
            .O(N__53208),
            .I(N__53195));
    InMux I__9015 (
            .O(N__53207),
            .I(N__53192));
    Span4Mux_h I__9014 (
            .O(N__53204),
            .I(N__53189));
    LocalMux I__9013 (
            .O(N__53201),
            .I(\c0.data_in_frame_12_4 ));
    LocalMux I__9012 (
            .O(N__53198),
            .I(\c0.data_in_frame_12_4 ));
    Odrv12 I__9011 (
            .O(N__53195),
            .I(\c0.data_in_frame_12_4 ));
    LocalMux I__9010 (
            .O(N__53192),
            .I(\c0.data_in_frame_12_4 ));
    Odrv4 I__9009 (
            .O(N__53189),
            .I(\c0.data_in_frame_12_4 ));
    CascadeMux I__9008 (
            .O(N__53178),
            .I(\c0.n33768_cascade_ ));
    InMux I__9007 (
            .O(N__53175),
            .I(N__53171));
    InMux I__9006 (
            .O(N__53174),
            .I(N__53168));
    LocalMux I__9005 (
            .O(N__53171),
            .I(N__53165));
    LocalMux I__9004 (
            .O(N__53168),
            .I(N__53162));
    Span4Mux_v I__9003 (
            .O(N__53165),
            .I(N__53159));
    Odrv4 I__9002 (
            .O(N__53162),
            .I(\c0.n33417 ));
    Odrv4 I__9001 (
            .O(N__53159),
            .I(\c0.n33417 ));
    InMux I__9000 (
            .O(N__53154),
            .I(N__53150));
    InMux I__8999 (
            .O(N__53153),
            .I(N__53147));
    LocalMux I__8998 (
            .O(N__53150),
            .I(N__53142));
    LocalMux I__8997 (
            .O(N__53147),
            .I(N__53142));
    Span4Mux_v I__8996 (
            .O(N__53142),
            .I(N__53139));
    Odrv4 I__8995 (
            .O(N__53139),
            .I(\c0.n6023 ));
    InMux I__8994 (
            .O(N__53136),
            .I(N__53133));
    LocalMux I__8993 (
            .O(N__53133),
            .I(N__53130));
    Span4Mux_v I__8992 (
            .O(N__53130),
            .I(N__53126));
    CascadeMux I__8991 (
            .O(N__53129),
            .I(N__53122));
    Sp12to4 I__8990 (
            .O(N__53126),
            .I(N__53118));
    InMux I__8989 (
            .O(N__53125),
            .I(N__53115));
    InMux I__8988 (
            .O(N__53122),
            .I(N__53110));
    InMux I__8987 (
            .O(N__53121),
            .I(N__53110));
    Odrv12 I__8986 (
            .O(N__53118),
            .I(\c0.data_in_frame_15_7 ));
    LocalMux I__8985 (
            .O(N__53115),
            .I(\c0.data_in_frame_15_7 ));
    LocalMux I__8984 (
            .O(N__53110),
            .I(\c0.data_in_frame_15_7 ));
    CascadeMux I__8983 (
            .O(N__53103),
            .I(N__53100));
    InMux I__8982 (
            .O(N__53100),
            .I(N__53093));
    InMux I__8981 (
            .O(N__53099),
            .I(N__53088));
    InMux I__8980 (
            .O(N__53098),
            .I(N__53088));
    InMux I__8979 (
            .O(N__53097),
            .I(N__53085));
    InMux I__8978 (
            .O(N__53096),
            .I(N__53082));
    LocalMux I__8977 (
            .O(N__53093),
            .I(N__53077));
    LocalMux I__8976 (
            .O(N__53088),
            .I(N__53077));
    LocalMux I__8975 (
            .O(N__53085),
            .I(\c0.data_in_frame_13_6 ));
    LocalMux I__8974 (
            .O(N__53082),
            .I(\c0.data_in_frame_13_6 ));
    Odrv4 I__8973 (
            .O(N__53077),
            .I(\c0.data_in_frame_13_6 ));
    InMux I__8972 (
            .O(N__53070),
            .I(N__53067));
    LocalMux I__8971 (
            .O(N__53067),
            .I(N__53064));
    Span4Mux_v I__8970 (
            .O(N__53064),
            .I(N__53061));
    Odrv4 I__8969 (
            .O(N__53061),
            .I(\c0.n6_adj_4715 ));
    CascadeMux I__8968 (
            .O(N__53058),
            .I(\c0.n31480_cascade_ ));
    InMux I__8967 (
            .O(N__53055),
            .I(N__53051));
    InMux I__8966 (
            .O(N__53054),
            .I(N__53048));
    LocalMux I__8965 (
            .O(N__53051),
            .I(N__53045));
    LocalMux I__8964 (
            .O(N__53048),
            .I(N__53039));
    Span4Mux_h I__8963 (
            .O(N__53045),
            .I(N__53039));
    InMux I__8962 (
            .O(N__53044),
            .I(N__53036));
    Odrv4 I__8961 (
            .O(N__53039),
            .I(\c0.n33422 ));
    LocalMux I__8960 (
            .O(N__53036),
            .I(\c0.n33422 ));
    InMux I__8959 (
            .O(N__53031),
            .I(N__53028));
    LocalMux I__8958 (
            .O(N__53028),
            .I(N__53024));
    CascadeMux I__8957 (
            .O(N__53027),
            .I(N__53018));
    Span4Mux_h I__8956 (
            .O(N__53024),
            .I(N__53014));
    InMux I__8955 (
            .O(N__53023),
            .I(N__53011));
    InMux I__8954 (
            .O(N__53022),
            .I(N__53006));
    InMux I__8953 (
            .O(N__53021),
            .I(N__53006));
    InMux I__8952 (
            .O(N__53018),
            .I(N__53001));
    InMux I__8951 (
            .O(N__53017),
            .I(N__53001));
    Odrv4 I__8950 (
            .O(N__53014),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__8949 (
            .O(N__53011),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__8948 (
            .O(N__53006),
            .I(\c0.data_in_frame_13_5 ));
    LocalMux I__8947 (
            .O(N__53001),
            .I(\c0.data_in_frame_13_5 ));
    CascadeMux I__8946 (
            .O(N__52992),
            .I(N__52989));
    InMux I__8945 (
            .O(N__52989),
            .I(N__52985));
    InMux I__8944 (
            .O(N__52988),
            .I(N__52982));
    LocalMux I__8943 (
            .O(N__52985),
            .I(\c0.n33610 ));
    LocalMux I__8942 (
            .O(N__52982),
            .I(\c0.n33610 ));
    InMux I__8941 (
            .O(N__52977),
            .I(N__52973));
    InMux I__8940 (
            .O(N__52976),
            .I(N__52970));
    LocalMux I__8939 (
            .O(N__52973),
            .I(N__52967));
    LocalMux I__8938 (
            .O(N__52970),
            .I(N__52964));
    Span4Mux_v I__8937 (
            .O(N__52967),
            .I(N__52961));
    Odrv4 I__8936 (
            .O(N__52964),
            .I(\c0.n35077 ));
    Odrv4 I__8935 (
            .O(N__52961),
            .I(\c0.n35077 ));
    InMux I__8934 (
            .O(N__52956),
            .I(N__52952));
    CascadeMux I__8933 (
            .O(N__52955),
            .I(N__52949));
    LocalMux I__8932 (
            .O(N__52952),
            .I(N__52944));
    InMux I__8931 (
            .O(N__52949),
            .I(N__52937));
    InMux I__8930 (
            .O(N__52948),
            .I(N__52937));
    InMux I__8929 (
            .O(N__52947),
            .I(N__52937));
    Odrv12 I__8928 (
            .O(N__52944),
            .I(\c0.data_in_frame_13_0 ));
    LocalMux I__8927 (
            .O(N__52937),
            .I(\c0.data_in_frame_13_0 ));
    InMux I__8926 (
            .O(N__52932),
            .I(N__52929));
    LocalMux I__8925 (
            .O(N__52929),
            .I(N__52926));
    Span4Mux_h I__8924 (
            .O(N__52926),
            .I(N__52923));
    Odrv4 I__8923 (
            .O(N__52923),
            .I(\c0.n12_adj_4714 ));
    CascadeMux I__8922 (
            .O(N__52920),
            .I(\c0.n33913_cascade_ ));
    InMux I__8921 (
            .O(N__52917),
            .I(N__52914));
    LocalMux I__8920 (
            .O(N__52914),
            .I(\c0.n18881 ));
    InMux I__8919 (
            .O(N__52911),
            .I(N__52907));
    InMux I__8918 (
            .O(N__52910),
            .I(N__52904));
    LocalMux I__8917 (
            .O(N__52907),
            .I(N__52901));
    LocalMux I__8916 (
            .O(N__52904),
            .I(N__52898));
    Span4Mux_h I__8915 (
            .O(N__52901),
            .I(N__52895));
    Odrv4 I__8914 (
            .O(N__52898),
            .I(\c0.n18847 ));
    Odrv4 I__8913 (
            .O(N__52895),
            .I(\c0.n18847 ));
    CascadeMux I__8912 (
            .O(N__52890),
            .I(\c0.n16010_cascade_ ));
    InMux I__8911 (
            .O(N__52887),
            .I(N__52884));
    LocalMux I__8910 (
            .O(N__52884),
            .I(N__52881));
    Span4Mux_v I__8909 (
            .O(N__52881),
            .I(N__52876));
    InMux I__8908 (
            .O(N__52880),
            .I(N__52873));
    InMux I__8907 (
            .O(N__52879),
            .I(N__52870));
    Odrv4 I__8906 (
            .O(N__52876),
            .I(\c0.n31526 ));
    LocalMux I__8905 (
            .O(N__52873),
            .I(\c0.n31526 ));
    LocalMux I__8904 (
            .O(N__52870),
            .I(\c0.n31526 ));
    InMux I__8903 (
            .O(N__52863),
            .I(N__52860));
    LocalMux I__8902 (
            .O(N__52860),
            .I(N__52856));
    InMux I__8901 (
            .O(N__52859),
            .I(N__52853));
    Span4Mux_v I__8900 (
            .O(N__52856),
            .I(N__52850));
    LocalMux I__8899 (
            .O(N__52853),
            .I(\c0.n33591 ));
    Odrv4 I__8898 (
            .O(N__52850),
            .I(\c0.n33591 ));
    CascadeMux I__8897 (
            .O(N__52845),
            .I(\c0.n32241_cascade_ ));
    InMux I__8896 (
            .O(N__52842),
            .I(N__52836));
    InMux I__8895 (
            .O(N__52841),
            .I(N__52836));
    LocalMux I__8894 (
            .O(N__52836),
            .I(\c0.n16010 ));
    InMux I__8893 (
            .O(N__52833),
            .I(N__52827));
    InMux I__8892 (
            .O(N__52832),
            .I(N__52824));
    InMux I__8891 (
            .O(N__52831),
            .I(N__52818));
    InMux I__8890 (
            .O(N__52830),
            .I(N__52818));
    LocalMux I__8889 (
            .O(N__52827),
            .I(N__52815));
    LocalMux I__8888 (
            .O(N__52824),
            .I(N__52812));
    InMux I__8887 (
            .O(N__52823),
            .I(N__52809));
    LocalMux I__8886 (
            .O(N__52818),
            .I(N__52806));
    Span4Mux_v I__8885 (
            .O(N__52815),
            .I(N__52802));
    Span4Mux_v I__8884 (
            .O(N__52812),
            .I(N__52799));
    LocalMux I__8883 (
            .O(N__52809),
            .I(N__52796));
    Span4Mux_h I__8882 (
            .O(N__52806),
            .I(N__52793));
    InMux I__8881 (
            .O(N__52805),
            .I(N__52790));
    Odrv4 I__8880 (
            .O(N__52802),
            .I(\c0.n18805 ));
    Odrv4 I__8879 (
            .O(N__52799),
            .I(\c0.n18805 ));
    Odrv4 I__8878 (
            .O(N__52796),
            .I(\c0.n18805 ));
    Odrv4 I__8877 (
            .O(N__52793),
            .I(\c0.n18805 ));
    LocalMux I__8876 (
            .O(N__52790),
            .I(\c0.n18805 ));
    CascadeMux I__8875 (
            .O(N__52779),
            .I(N__52776));
    InMux I__8874 (
            .O(N__52776),
            .I(N__52773));
    LocalMux I__8873 (
            .O(N__52773),
            .I(N__52769));
    InMux I__8872 (
            .O(N__52772),
            .I(N__52766));
    Odrv12 I__8871 (
            .O(N__52769),
            .I(\c0.n34012 ));
    LocalMux I__8870 (
            .O(N__52766),
            .I(\c0.n34012 ));
    InMux I__8869 (
            .O(N__52761),
            .I(N__52758));
    LocalMux I__8868 (
            .O(N__52758),
            .I(N__52753));
    InMux I__8867 (
            .O(N__52757),
            .I(N__52750));
    InMux I__8866 (
            .O(N__52756),
            .I(N__52747));
    Span4Mux_v I__8865 (
            .O(N__52753),
            .I(N__52744));
    LocalMux I__8864 (
            .O(N__52750),
            .I(N__52740));
    LocalMux I__8863 (
            .O(N__52747),
            .I(N__52737));
    Span4Mux_h I__8862 (
            .O(N__52744),
            .I(N__52734));
    InMux I__8861 (
            .O(N__52743),
            .I(N__52731));
    Odrv12 I__8860 (
            .O(N__52740),
            .I(\c0.n18438 ));
    Odrv4 I__8859 (
            .O(N__52737),
            .I(\c0.n18438 ));
    Odrv4 I__8858 (
            .O(N__52734),
            .I(\c0.n18438 ));
    LocalMux I__8857 (
            .O(N__52731),
            .I(\c0.n18438 ));
    InMux I__8856 (
            .O(N__52722),
            .I(N__52718));
    InMux I__8855 (
            .O(N__52721),
            .I(N__52715));
    LocalMux I__8854 (
            .O(N__52718),
            .I(N__52712));
    LocalMux I__8853 (
            .O(N__52715),
            .I(\c0.n33629 ));
    Odrv4 I__8852 (
            .O(N__52712),
            .I(\c0.n33629 ));
    InMux I__8851 (
            .O(N__52707),
            .I(N__52698));
    InMux I__8850 (
            .O(N__52706),
            .I(N__52698));
    InMux I__8849 (
            .O(N__52705),
            .I(N__52698));
    LocalMux I__8848 (
            .O(N__52698),
            .I(\c0.data_in_frame_15_2 ));
    CascadeMux I__8847 (
            .O(N__52695),
            .I(N__52692));
    InMux I__8846 (
            .O(N__52692),
            .I(N__52689));
    LocalMux I__8845 (
            .O(N__52689),
            .I(N__52686));
    Odrv4 I__8844 (
            .O(N__52686),
            .I(\c0.n33321 ));
    InMux I__8843 (
            .O(N__52683),
            .I(N__52678));
    CascadeMux I__8842 (
            .O(N__52682),
            .I(N__52675));
    InMux I__8841 (
            .O(N__52681),
            .I(N__52672));
    LocalMux I__8840 (
            .O(N__52678),
            .I(N__52669));
    InMux I__8839 (
            .O(N__52675),
            .I(N__52666));
    LocalMux I__8838 (
            .O(N__52672),
            .I(N__52663));
    Span4Mux_h I__8837 (
            .O(N__52669),
            .I(N__52660));
    LocalMux I__8836 (
            .O(N__52666),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__8835 (
            .O(N__52663),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__8834 (
            .O(N__52660),
            .I(\c0.data_in_frame_3_7 ));
    InMux I__8833 (
            .O(N__52653),
            .I(N__52648));
    InMux I__8832 (
            .O(N__52652),
            .I(N__52645));
    CascadeMux I__8831 (
            .O(N__52651),
            .I(N__52642));
    LocalMux I__8830 (
            .O(N__52648),
            .I(N__52637));
    LocalMux I__8829 (
            .O(N__52645),
            .I(N__52637));
    InMux I__8828 (
            .O(N__52642),
            .I(N__52634));
    Span4Mux_h I__8827 (
            .O(N__52637),
            .I(N__52631));
    LocalMux I__8826 (
            .O(N__52634),
            .I(\c0.data_in_frame_15_6 ));
    Odrv4 I__8825 (
            .O(N__52631),
            .I(\c0.data_in_frame_15_6 ));
    CascadeMux I__8824 (
            .O(N__52626),
            .I(N__52623));
    InMux I__8823 (
            .O(N__52623),
            .I(N__52618));
    InMux I__8822 (
            .O(N__52622),
            .I(N__52615));
    InMux I__8821 (
            .O(N__52621),
            .I(N__52612));
    LocalMux I__8820 (
            .O(N__52618),
            .I(\c0.data_in_frame_12_1 ));
    LocalMux I__8819 (
            .O(N__52615),
            .I(\c0.data_in_frame_12_1 ));
    LocalMux I__8818 (
            .O(N__52612),
            .I(\c0.data_in_frame_12_1 ));
    InMux I__8817 (
            .O(N__52605),
            .I(N__52601));
    InMux I__8816 (
            .O(N__52604),
            .I(N__52598));
    LocalMux I__8815 (
            .O(N__52601),
            .I(N__52595));
    LocalMux I__8814 (
            .O(N__52598),
            .I(N__52592));
    Span4Mux_v I__8813 (
            .O(N__52595),
            .I(N__52589));
    Span4Mux_h I__8812 (
            .O(N__52592),
            .I(N__52586));
    Odrv4 I__8811 (
            .O(N__52589),
            .I(\c0.n33843 ));
    Odrv4 I__8810 (
            .O(N__52586),
            .I(\c0.n33843 ));
    InMux I__8809 (
            .O(N__52581),
            .I(N__52578));
    LocalMux I__8808 (
            .O(N__52578),
            .I(N__52575));
    Span4Mux_v I__8807 (
            .O(N__52575),
            .I(N__52572));
    Odrv4 I__8806 (
            .O(N__52572),
            .I(\c0.n31_adj_4740 ));
    InMux I__8805 (
            .O(N__52569),
            .I(N__52566));
    LocalMux I__8804 (
            .O(N__52566),
            .I(N__52563));
    Span4Mux_h I__8803 (
            .O(N__52563),
            .I(N__52560));
    Odrv4 I__8802 (
            .O(N__52560),
            .I(n4_adj_4807));
    CascadeMux I__8801 (
            .O(N__52557),
            .I(n4_adj_4807_cascade_));
    InMux I__8800 (
            .O(N__52554),
            .I(N__52551));
    LocalMux I__8799 (
            .O(N__52551),
            .I(N__52548));
    Span4Mux_h I__8798 (
            .O(N__52548),
            .I(N__52545));
    Span4Mux_h I__8797 (
            .O(N__52545),
            .I(N__52539));
    InMux I__8796 (
            .O(N__52544),
            .I(N__52532));
    InMux I__8795 (
            .O(N__52543),
            .I(N__52532));
    InMux I__8794 (
            .O(N__52542),
            .I(N__52532));
    Span4Mux_h I__8793 (
            .O(N__52539),
            .I(N__52529));
    LocalMux I__8792 (
            .O(N__52532),
            .I(n18031));
    Odrv4 I__8791 (
            .O(N__52529),
            .I(n18031));
    InMux I__8790 (
            .O(N__52524),
            .I(N__52520));
    InMux I__8789 (
            .O(N__52523),
            .I(N__52516));
    LocalMux I__8788 (
            .O(N__52520),
            .I(N__52513));
    InMux I__8787 (
            .O(N__52519),
            .I(N__52510));
    LocalMux I__8786 (
            .O(N__52516),
            .I(N__52506));
    Span4Mux_h I__8785 (
            .O(N__52513),
            .I(N__52503));
    LocalMux I__8784 (
            .O(N__52510),
            .I(N__52500));
    InMux I__8783 (
            .O(N__52509),
            .I(N__52497));
    Span4Mux_h I__8782 (
            .O(N__52506),
            .I(N__52494));
    Sp12to4 I__8781 (
            .O(N__52503),
            .I(N__52489));
    Span12Mux_h I__8780 (
            .O(N__52500),
            .I(N__52489));
    LocalMux I__8779 (
            .O(N__52497),
            .I(\c0.data_in_frame_5_2 ));
    Odrv4 I__8778 (
            .O(N__52494),
            .I(\c0.data_in_frame_5_2 ));
    Odrv12 I__8777 (
            .O(N__52489),
            .I(\c0.data_in_frame_5_2 ));
    InMux I__8776 (
            .O(N__52482),
            .I(N__52478));
    InMux I__8775 (
            .O(N__52481),
            .I(N__52474));
    LocalMux I__8774 (
            .O(N__52478),
            .I(N__52471));
    CascadeMux I__8773 (
            .O(N__52477),
            .I(N__52468));
    LocalMux I__8772 (
            .O(N__52474),
            .I(N__52465));
    Span4Mux_v I__8771 (
            .O(N__52471),
            .I(N__52462));
    InMux I__8770 (
            .O(N__52468),
            .I(N__52459));
    Span4Mux_v I__8769 (
            .O(N__52465),
            .I(N__52456));
    Span4Mux_h I__8768 (
            .O(N__52462),
            .I(N__52453));
    LocalMux I__8767 (
            .O(N__52459),
            .I(N__52448));
    Span4Mux_h I__8766 (
            .O(N__52456),
            .I(N__52448));
    Odrv4 I__8765 (
            .O(N__52453),
            .I(\c0.data_in_frame_14_3 ));
    Odrv4 I__8764 (
            .O(N__52448),
            .I(\c0.data_in_frame_14_3 ));
    InMux I__8763 (
            .O(N__52443),
            .I(N__52440));
    LocalMux I__8762 (
            .O(N__52440),
            .I(N__52437));
    Odrv12 I__8761 (
            .O(N__52437),
            .I(\c0.n6_adj_4546 ));
    InMux I__8760 (
            .O(N__52434),
            .I(N__52430));
    InMux I__8759 (
            .O(N__52433),
            .I(N__52427));
    LocalMux I__8758 (
            .O(N__52430),
            .I(N__52421));
    LocalMux I__8757 (
            .O(N__52427),
            .I(N__52421));
    InMux I__8756 (
            .O(N__52426),
            .I(N__52418));
    Span4Mux_v I__8755 (
            .O(N__52421),
            .I(N__52415));
    LocalMux I__8754 (
            .O(N__52418),
            .I(\c0.data_in_frame_4_0 ));
    Odrv4 I__8753 (
            .O(N__52415),
            .I(\c0.data_in_frame_4_0 ));
    InMux I__8752 (
            .O(N__52410),
            .I(N__52407));
    LocalMux I__8751 (
            .O(N__52407),
            .I(\c0.n18663 ));
    CascadeMux I__8750 (
            .O(N__52404),
            .I(\c0.n33344_cascade_ ));
    InMux I__8749 (
            .O(N__52401),
            .I(N__52398));
    LocalMux I__8748 (
            .O(N__52398),
            .I(N__52393));
    InMux I__8747 (
            .O(N__52397),
            .I(N__52390));
    CascadeMux I__8746 (
            .O(N__52396),
            .I(N__52386));
    Span4Mux_h I__8745 (
            .O(N__52393),
            .I(N__52381));
    LocalMux I__8744 (
            .O(N__52390),
            .I(N__52381));
    InMux I__8743 (
            .O(N__52389),
            .I(N__52378));
    InMux I__8742 (
            .O(N__52386),
            .I(N__52375));
    Span4Mux_v I__8741 (
            .O(N__52381),
            .I(N__52372));
    LocalMux I__8740 (
            .O(N__52378),
            .I(N__52369));
    LocalMux I__8739 (
            .O(N__52375),
            .I(\c0.data_in_frame_3_6 ));
    Odrv4 I__8738 (
            .O(N__52372),
            .I(\c0.data_in_frame_3_6 ));
    Odrv4 I__8737 (
            .O(N__52369),
            .I(\c0.data_in_frame_3_6 ));
    CascadeMux I__8736 (
            .O(N__52362),
            .I(\c0.n10_adj_4770_cascade_ ));
    InMux I__8735 (
            .O(N__52359),
            .I(N__52356));
    LocalMux I__8734 (
            .O(N__52356),
            .I(N__52351));
    InMux I__8733 (
            .O(N__52355),
            .I(N__52346));
    InMux I__8732 (
            .O(N__52354),
            .I(N__52343));
    Span4Mux_v I__8731 (
            .O(N__52351),
            .I(N__52340));
    InMux I__8730 (
            .O(N__52350),
            .I(N__52335));
    InMux I__8729 (
            .O(N__52349),
            .I(N__52335));
    LocalMux I__8728 (
            .O(N__52346),
            .I(N__52332));
    LocalMux I__8727 (
            .O(N__52343),
            .I(N__52329));
    Span4Mux_h I__8726 (
            .O(N__52340),
            .I(N__52324));
    LocalMux I__8725 (
            .O(N__52335),
            .I(N__52324));
    Span12Mux_h I__8724 (
            .O(N__52332),
            .I(N__52321));
    Odrv4 I__8723 (
            .O(N__52329),
            .I(\c0.n18314 ));
    Odrv4 I__8722 (
            .O(N__52324),
            .I(\c0.n18314 ));
    Odrv12 I__8721 (
            .O(N__52321),
            .I(\c0.n18314 ));
    CascadeMux I__8720 (
            .O(N__52314),
            .I(N__52311));
    InMux I__8719 (
            .O(N__52311),
            .I(N__52305));
    InMux I__8718 (
            .O(N__52310),
            .I(N__52305));
    LocalMux I__8717 (
            .O(N__52305),
            .I(\c0.data_in_frame_6_2 ));
    InMux I__8716 (
            .O(N__52302),
            .I(N__52299));
    LocalMux I__8715 (
            .O(N__52299),
            .I(N__52296));
    Span4Mux_h I__8714 (
            .O(N__52296),
            .I(N__52292));
    CascadeMux I__8713 (
            .O(N__52295),
            .I(N__52288));
    Span4Mux_h I__8712 (
            .O(N__52292),
            .I(N__52284));
    InMux I__8711 (
            .O(N__52291),
            .I(N__52281));
    InMux I__8710 (
            .O(N__52288),
            .I(N__52276));
    InMux I__8709 (
            .O(N__52287),
            .I(N__52276));
    Odrv4 I__8708 (
            .O(N__52284),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__8707 (
            .O(N__52281),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__8706 (
            .O(N__52276),
            .I(\c0.data_in_frame_4_3 ));
    CascadeMux I__8705 (
            .O(N__52269),
            .I(N__52265));
    InMux I__8704 (
            .O(N__52268),
            .I(N__52262));
    InMux I__8703 (
            .O(N__52265),
            .I(N__52256));
    LocalMux I__8702 (
            .O(N__52262),
            .I(N__52253));
    InMux I__8701 (
            .O(N__52261),
            .I(N__52250));
    InMux I__8700 (
            .O(N__52260),
            .I(N__52245));
    InMux I__8699 (
            .O(N__52259),
            .I(N__52245));
    LocalMux I__8698 (
            .O(N__52256),
            .I(\c0.data_in_frame_2_0 ));
    Odrv4 I__8697 (
            .O(N__52253),
            .I(\c0.data_in_frame_2_0 ));
    LocalMux I__8696 (
            .O(N__52250),
            .I(\c0.data_in_frame_2_0 ));
    LocalMux I__8695 (
            .O(N__52245),
            .I(\c0.data_in_frame_2_0 ));
    InMux I__8694 (
            .O(N__52236),
            .I(N__52233));
    LocalMux I__8693 (
            .O(N__52233),
            .I(\c0.n33692 ));
    CascadeMux I__8692 (
            .O(N__52230),
            .I(\c0.rx.n6_cascade_ ));
    CascadeMux I__8691 (
            .O(N__52227),
            .I(\c0.rx.n35949_cascade_ ));
    CascadeMux I__8690 (
            .O(N__52224),
            .I(\c0.n18663_cascade_ ));
    CascadeMux I__8689 (
            .O(N__52221),
            .I(\c0.n33397_cascade_ ));
    InMux I__8688 (
            .O(N__52218),
            .I(N__52215));
    LocalMux I__8687 (
            .O(N__52215),
            .I(N__52211));
    InMux I__8686 (
            .O(N__52214),
            .I(N__52208));
    Span4Mux_v I__8685 (
            .O(N__52211),
            .I(N__52203));
    LocalMux I__8684 (
            .O(N__52208),
            .I(N__52203));
    Odrv4 I__8683 (
            .O(N__52203),
            .I(\c0.n33604 ));
    InMux I__8682 (
            .O(N__52200),
            .I(N__52196));
    InMux I__8681 (
            .O(N__52199),
            .I(N__52193));
    LocalMux I__8680 (
            .O(N__52196),
            .I(N__52187));
    LocalMux I__8679 (
            .O(N__52193),
            .I(N__52187));
    CascadeMux I__8678 (
            .O(N__52192),
            .I(N__52184));
    Span4Mux_v I__8677 (
            .O(N__52187),
            .I(N__52181));
    InMux I__8676 (
            .O(N__52184),
            .I(N__52178));
    Span4Mux_h I__8675 (
            .O(N__52181),
            .I(N__52175));
    LocalMux I__8674 (
            .O(N__52178),
            .I(\c0.data_in_frame_9_0 ));
    Odrv4 I__8673 (
            .O(N__52175),
            .I(\c0.data_in_frame_9_0 ));
    InMux I__8672 (
            .O(N__52170),
            .I(N__52167));
    LocalMux I__8671 (
            .O(N__52167),
            .I(N__52163));
    CascadeMux I__8670 (
            .O(N__52166),
            .I(N__52159));
    Span4Mux_h I__8669 (
            .O(N__52163),
            .I(N__52155));
    CascadeMux I__8668 (
            .O(N__52162),
            .I(N__52150));
    InMux I__8667 (
            .O(N__52159),
            .I(N__52144));
    InMux I__8666 (
            .O(N__52158),
            .I(N__52144));
    Span4Mux_h I__8665 (
            .O(N__52155),
            .I(N__52141));
    InMux I__8664 (
            .O(N__52154),
            .I(N__52136));
    InMux I__8663 (
            .O(N__52153),
            .I(N__52136));
    InMux I__8662 (
            .O(N__52150),
            .I(N__52131));
    InMux I__8661 (
            .O(N__52149),
            .I(N__52131));
    LocalMux I__8660 (
            .O(N__52144),
            .I(\c0.data_in_frame_0_2 ));
    Odrv4 I__8659 (
            .O(N__52141),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__8658 (
            .O(N__52136),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__8657 (
            .O(N__52131),
            .I(\c0.data_in_frame_0_2 ));
    CascadeMux I__8656 (
            .O(N__52122),
            .I(N__52116));
    InMux I__8655 (
            .O(N__52121),
            .I(N__52113));
    InMux I__8654 (
            .O(N__52120),
            .I(N__52110));
    CascadeMux I__8653 (
            .O(N__52119),
            .I(N__52107));
    InMux I__8652 (
            .O(N__52116),
            .I(N__52099));
    LocalMux I__8651 (
            .O(N__52113),
            .I(N__52096));
    LocalMux I__8650 (
            .O(N__52110),
            .I(N__52093));
    InMux I__8649 (
            .O(N__52107),
            .I(N__52088));
    InMux I__8648 (
            .O(N__52106),
            .I(N__52088));
    InMux I__8647 (
            .O(N__52105),
            .I(N__52079));
    InMux I__8646 (
            .O(N__52104),
            .I(N__52079));
    InMux I__8645 (
            .O(N__52103),
            .I(N__52079));
    InMux I__8644 (
            .O(N__52102),
            .I(N__52079));
    LocalMux I__8643 (
            .O(N__52099),
            .I(N__52072));
    Span4Mux_h I__8642 (
            .O(N__52096),
            .I(N__52072));
    Span4Mux_h I__8641 (
            .O(N__52093),
            .I(N__52072));
    LocalMux I__8640 (
            .O(N__52088),
            .I(\c0.data_in_frame_0_3 ));
    LocalMux I__8639 (
            .O(N__52079),
            .I(\c0.data_in_frame_0_3 ));
    Odrv4 I__8638 (
            .O(N__52072),
            .I(\c0.data_in_frame_0_3 ));
    CascadeMux I__8637 (
            .O(N__52065),
            .I(N__52056));
    InMux I__8636 (
            .O(N__52064),
            .I(N__52053));
    CascadeMux I__8635 (
            .O(N__52063),
            .I(N__52049));
    InMux I__8634 (
            .O(N__52062),
            .I(N__52044));
    InMux I__8633 (
            .O(N__52061),
            .I(N__52044));
    InMux I__8632 (
            .O(N__52060),
            .I(N__52039));
    InMux I__8631 (
            .O(N__52059),
            .I(N__52039));
    InMux I__8630 (
            .O(N__52056),
            .I(N__52036));
    LocalMux I__8629 (
            .O(N__52053),
            .I(N__52033));
    InMux I__8628 (
            .O(N__52052),
            .I(N__52030));
    InMux I__8627 (
            .O(N__52049),
            .I(N__52027));
    LocalMux I__8626 (
            .O(N__52044),
            .I(N__52022));
    LocalMux I__8625 (
            .O(N__52039),
            .I(N__52022));
    LocalMux I__8624 (
            .O(N__52036),
            .I(\c0.data_in_frame_0_1 ));
    Odrv4 I__8623 (
            .O(N__52033),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8622 (
            .O(N__52030),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8621 (
            .O(N__52027),
            .I(\c0.data_in_frame_0_1 ));
    Odrv12 I__8620 (
            .O(N__52022),
            .I(\c0.data_in_frame_0_1 ));
    InMux I__8619 (
            .O(N__52011),
            .I(N__52008));
    LocalMux I__8618 (
            .O(N__52008),
            .I(\c0.n28 ));
    InMux I__8617 (
            .O(N__52005),
            .I(N__52002));
    LocalMux I__8616 (
            .O(N__52002),
            .I(\c0.n32 ));
    CascadeMux I__8615 (
            .O(N__51999),
            .I(N__51996));
    InMux I__8614 (
            .O(N__51996),
            .I(N__51992));
    InMux I__8613 (
            .O(N__51995),
            .I(N__51989));
    LocalMux I__8612 (
            .O(N__51992),
            .I(\c0.data_in_frame_6_3 ));
    LocalMux I__8611 (
            .O(N__51989),
            .I(\c0.data_in_frame_6_3 ));
    InMux I__8610 (
            .O(N__51984),
            .I(N__51978));
    InMux I__8609 (
            .O(N__51983),
            .I(N__51978));
    LocalMux I__8608 (
            .O(N__51978),
            .I(data_out_frame_5_2));
    InMux I__8607 (
            .O(N__51975),
            .I(N__51969));
    InMux I__8606 (
            .O(N__51974),
            .I(N__51969));
    LocalMux I__8605 (
            .O(N__51969),
            .I(data_out_frame_6_0));
    InMux I__8604 (
            .O(N__51966),
            .I(N__51960));
    InMux I__8603 (
            .O(N__51965),
            .I(N__51960));
    LocalMux I__8602 (
            .O(N__51960),
            .I(data_out_frame_7_0));
    InMux I__8601 (
            .O(N__51957),
            .I(N__51954));
    LocalMux I__8600 (
            .O(N__51954),
            .I(N__51950));
    InMux I__8599 (
            .O(N__51953),
            .I(N__51947));
    Odrv4 I__8598 (
            .O(N__51950),
            .I(\c0.n27710 ));
    LocalMux I__8597 (
            .O(N__51947),
            .I(\c0.n27710 ));
    SRMux I__8596 (
            .O(N__51942),
            .I(N__51939));
    LocalMux I__8595 (
            .O(N__51939),
            .I(N__51935));
    InMux I__8594 (
            .O(N__51938),
            .I(N__51932));
    Span4Mux_v I__8593 (
            .O(N__51935),
            .I(N__51926));
    LocalMux I__8592 (
            .O(N__51932),
            .I(N__51926));
    InMux I__8591 (
            .O(N__51931),
            .I(N__51923));
    Span4Mux_h I__8590 (
            .O(N__51926),
            .I(N__51920));
    LocalMux I__8589 (
            .O(N__51923),
            .I(N__51917));
    Span4Mux_h I__8588 (
            .O(N__51920),
            .I(N__51914));
    Span4Mux_h I__8587 (
            .O(N__51917),
            .I(N__51911));
    Odrv4 I__8586 (
            .O(N__51914),
            .I(\c0.n34190 ));
    Odrv4 I__8585 (
            .O(N__51911),
            .I(\c0.n34190 ));
    CascadeMux I__8584 (
            .O(N__51906),
            .I(N__51902));
    InMux I__8583 (
            .O(N__51905),
            .I(N__51894));
    InMux I__8582 (
            .O(N__51902),
            .I(N__51889));
    InMux I__8581 (
            .O(N__51901),
            .I(N__51889));
    InMux I__8580 (
            .O(N__51900),
            .I(N__51886));
    InMux I__8579 (
            .O(N__51899),
            .I(N__51881));
    InMux I__8578 (
            .O(N__51898),
            .I(N__51881));
    InMux I__8577 (
            .O(N__51897),
            .I(N__51878));
    LocalMux I__8576 (
            .O(N__51894),
            .I(N__51873));
    LocalMux I__8575 (
            .O(N__51889),
            .I(N__51873));
    LocalMux I__8574 (
            .O(N__51886),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    LocalMux I__8573 (
            .O(N__51881),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    LocalMux I__8572 (
            .O(N__51878),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    Odrv4 I__8571 (
            .O(N__51873),
            .I(\c0.data_out_frame_29_7_N_1483_0 ));
    CascadeMux I__8570 (
            .O(N__51864),
            .I(\c0.n12_cascade_ ));
    CascadeMux I__8569 (
            .O(N__51861),
            .I(N__51852));
    InMux I__8568 (
            .O(N__51860),
            .I(N__51847));
    InMux I__8567 (
            .O(N__51859),
            .I(N__51842));
    InMux I__8566 (
            .O(N__51858),
            .I(N__51842));
    InMux I__8565 (
            .O(N__51857),
            .I(N__51839));
    InMux I__8564 (
            .O(N__51856),
            .I(N__51831));
    InMux I__8563 (
            .O(N__51855),
            .I(N__51831));
    InMux I__8562 (
            .O(N__51852),
            .I(N__51828));
    InMux I__8561 (
            .O(N__51851),
            .I(N__51825));
    InMux I__8560 (
            .O(N__51850),
            .I(N__51822));
    LocalMux I__8559 (
            .O(N__51847),
            .I(N__51814));
    LocalMux I__8558 (
            .O(N__51842),
            .I(N__51814));
    LocalMux I__8557 (
            .O(N__51839),
            .I(N__51814));
    InMux I__8556 (
            .O(N__51838),
            .I(N__51811));
    InMux I__8555 (
            .O(N__51837),
            .I(N__51806));
    InMux I__8554 (
            .O(N__51836),
            .I(N__51806));
    LocalMux I__8553 (
            .O(N__51831),
            .I(N__51801));
    LocalMux I__8552 (
            .O(N__51828),
            .I(N__51801));
    LocalMux I__8551 (
            .O(N__51825),
            .I(N__51796));
    LocalMux I__8550 (
            .O(N__51822),
            .I(N__51796));
    InMux I__8549 (
            .O(N__51821),
            .I(N__51793));
    Span4Mux_v I__8548 (
            .O(N__51814),
            .I(N__51790));
    LocalMux I__8547 (
            .O(N__51811),
            .I(N__51787));
    LocalMux I__8546 (
            .O(N__51806),
            .I(N__51782));
    Span4Mux_h I__8545 (
            .O(N__51801),
            .I(N__51782));
    Span4Mux_v I__8544 (
            .O(N__51796),
            .I(N__51777));
    LocalMux I__8543 (
            .O(N__51793),
            .I(N__51777));
    Span4Mux_h I__8542 (
            .O(N__51790),
            .I(N__51774));
    Span4Mux_h I__8541 (
            .O(N__51787),
            .I(N__51769));
    Span4Mux_h I__8540 (
            .O(N__51782),
            .I(N__51769));
    Span4Mux_h I__8539 (
            .O(N__51777),
            .I(N__51766));
    Odrv4 I__8538 (
            .O(N__51774),
            .I(\c0.data_out_frame_29_7_N_1483_1 ));
    Odrv4 I__8537 (
            .O(N__51769),
            .I(\c0.data_out_frame_29_7_N_1483_1 ));
    Odrv4 I__8536 (
            .O(N__51766),
            .I(\c0.data_out_frame_29_7_N_1483_1 ));
    InMux I__8535 (
            .O(N__51759),
            .I(N__51753));
    InMux I__8534 (
            .O(N__51758),
            .I(N__51753));
    LocalMux I__8533 (
            .O(N__51753),
            .I(\c0.n19297 ));
    InMux I__8532 (
            .O(N__51750),
            .I(N__51742));
    InMux I__8531 (
            .O(N__51749),
            .I(N__51737));
    InMux I__8530 (
            .O(N__51748),
            .I(N__51737));
    CascadeMux I__8529 (
            .O(N__51747),
            .I(N__51734));
    InMux I__8528 (
            .O(N__51746),
            .I(N__51729));
    InMux I__8527 (
            .O(N__51745),
            .I(N__51729));
    LocalMux I__8526 (
            .O(N__51742),
            .I(N__51726));
    LocalMux I__8525 (
            .O(N__51737),
            .I(N__51723));
    InMux I__8524 (
            .O(N__51734),
            .I(N__51720));
    LocalMux I__8523 (
            .O(N__51729),
            .I(\c0.n3315 ));
    Odrv4 I__8522 (
            .O(N__51726),
            .I(\c0.n3315 ));
    Odrv4 I__8521 (
            .O(N__51723),
            .I(\c0.n3315 ));
    LocalMux I__8520 (
            .O(N__51720),
            .I(\c0.n3315 ));
    CascadeMux I__8519 (
            .O(N__51711),
            .I(\c0.n19297_cascade_ ));
    CascadeMux I__8518 (
            .O(N__51708),
            .I(N__51704));
    InMux I__8517 (
            .O(N__51707),
            .I(N__51701));
    InMux I__8516 (
            .O(N__51704),
            .I(N__51698));
    LocalMux I__8515 (
            .O(N__51701),
            .I(N__51690));
    LocalMux I__8514 (
            .O(N__51698),
            .I(N__51687));
    InMux I__8513 (
            .O(N__51697),
            .I(N__51679));
    InMux I__8512 (
            .O(N__51696),
            .I(N__51679));
    CascadeMux I__8511 (
            .O(N__51695),
            .I(N__51676));
    InMux I__8510 (
            .O(N__51694),
            .I(N__51673));
    InMux I__8509 (
            .O(N__51693),
            .I(N__51670));
    Span4Mux_h I__8508 (
            .O(N__51690),
            .I(N__51665));
    Span4Mux_h I__8507 (
            .O(N__51687),
            .I(N__51665));
    InMux I__8506 (
            .O(N__51686),
            .I(N__51662));
    InMux I__8505 (
            .O(N__51685),
            .I(N__51657));
    InMux I__8504 (
            .O(N__51684),
            .I(N__51657));
    LocalMux I__8503 (
            .O(N__51679),
            .I(N__51654));
    InMux I__8502 (
            .O(N__51676),
            .I(N__51651));
    LocalMux I__8501 (
            .O(N__51673),
            .I(N__51646));
    LocalMux I__8500 (
            .O(N__51670),
            .I(N__51646));
    Span4Mux_h I__8499 (
            .O(N__51665),
            .I(N__51643));
    LocalMux I__8498 (
            .O(N__51662),
            .I(N__51632));
    LocalMux I__8497 (
            .O(N__51657),
            .I(N__51632));
    Span12Mux_h I__8496 (
            .O(N__51654),
            .I(N__51632));
    LocalMux I__8495 (
            .O(N__51651),
            .I(N__51632));
    Span12Mux_v I__8494 (
            .O(N__51646),
            .I(N__51632));
    Odrv4 I__8493 (
            .O(N__51643),
            .I(\c0.data_out_frame_29_7_N_1483_2 ));
    Odrv12 I__8492 (
            .O(N__51632),
            .I(\c0.data_out_frame_29_7_N_1483_2 ));
    InMux I__8491 (
            .O(N__51627),
            .I(N__51624));
    LocalMux I__8490 (
            .O(N__51624),
            .I(N__51619));
    InMux I__8489 (
            .O(N__51623),
            .I(N__51616));
    CascadeMux I__8488 (
            .O(N__51622),
            .I(N__51613));
    Span4Mux_h I__8487 (
            .O(N__51619),
            .I(N__51610));
    LocalMux I__8486 (
            .O(N__51616),
            .I(N__51607));
    InMux I__8485 (
            .O(N__51613),
            .I(N__51604));
    Span4Mux_v I__8484 (
            .O(N__51610),
            .I(N__51601));
    Sp12to4 I__8483 (
            .O(N__51607),
            .I(N__51598));
    LocalMux I__8482 (
            .O(N__51604),
            .I(\c0.data_in_frame_14_0 ));
    Odrv4 I__8481 (
            .O(N__51601),
            .I(\c0.data_in_frame_14_0 ));
    Odrv12 I__8480 (
            .O(N__51598),
            .I(\c0.data_in_frame_14_0 ));
    InMux I__8479 (
            .O(N__51591),
            .I(N__51587));
    CascadeMux I__8478 (
            .O(N__51590),
            .I(N__51583));
    LocalMux I__8477 (
            .O(N__51587),
            .I(N__51580));
    InMux I__8476 (
            .O(N__51586),
            .I(N__51575));
    InMux I__8475 (
            .O(N__51583),
            .I(N__51575));
    Span4Mux_h I__8474 (
            .O(N__51580),
            .I(N__51572));
    LocalMux I__8473 (
            .O(N__51575),
            .I(N__51569));
    Span4Mux_h I__8472 (
            .O(N__51572),
            .I(N__51564));
    Span4Mux_h I__8471 (
            .O(N__51569),
            .I(N__51564));
    Odrv4 I__8470 (
            .O(N__51564),
            .I(\c0.n29675 ));
    InMux I__8469 (
            .O(N__51561),
            .I(N__51556));
    InMux I__8468 (
            .O(N__51560),
            .I(N__51553));
    InMux I__8467 (
            .O(N__51559),
            .I(N__51547));
    LocalMux I__8466 (
            .O(N__51556),
            .I(N__51544));
    LocalMux I__8465 (
            .O(N__51553),
            .I(N__51541));
    InMux I__8464 (
            .O(N__51552),
            .I(N__51538));
    InMux I__8463 (
            .O(N__51551),
            .I(N__51533));
    InMux I__8462 (
            .O(N__51550),
            .I(N__51533));
    LocalMux I__8461 (
            .O(N__51547),
            .I(\c0.n78 ));
    Odrv12 I__8460 (
            .O(N__51544),
            .I(\c0.n78 ));
    Odrv4 I__8459 (
            .O(N__51541),
            .I(\c0.n78 ));
    LocalMux I__8458 (
            .O(N__51538),
            .I(\c0.n78 ));
    LocalMux I__8457 (
            .O(N__51533),
            .I(\c0.n78 ));
    InMux I__8456 (
            .O(N__51522),
            .I(N__51517));
    InMux I__8455 (
            .O(N__51521),
            .I(N__51514));
    InMux I__8454 (
            .O(N__51520),
            .I(N__51511));
    LocalMux I__8453 (
            .O(N__51517),
            .I(N__51506));
    LocalMux I__8452 (
            .O(N__51514),
            .I(N__51503));
    LocalMux I__8451 (
            .O(N__51511),
            .I(N__51500));
    InMux I__8450 (
            .O(N__51510),
            .I(N__51495));
    InMux I__8449 (
            .O(N__51509),
            .I(N__51495));
    Span4Mux_h I__8448 (
            .O(N__51506),
            .I(N__51492));
    Odrv4 I__8447 (
            .O(N__51503),
            .I(\c0.data_out_frame_0__7__N_2571 ));
    Odrv12 I__8446 (
            .O(N__51500),
            .I(\c0.data_out_frame_0__7__N_2571 ));
    LocalMux I__8445 (
            .O(N__51495),
            .I(\c0.data_out_frame_0__7__N_2571 ));
    Odrv4 I__8444 (
            .O(N__51492),
            .I(\c0.data_out_frame_0__7__N_2571 ));
    CascadeMux I__8443 (
            .O(N__51483),
            .I(N__51480));
    InMux I__8442 (
            .O(N__51480),
            .I(N__51474));
    InMux I__8441 (
            .O(N__51479),
            .I(N__51474));
    LocalMux I__8440 (
            .O(N__51474),
            .I(\c0.data_out_frame_0_2 ));
    CascadeMux I__8439 (
            .O(N__51471),
            .I(\c0.n35960_cascade_ ));
    CascadeMux I__8438 (
            .O(N__51468),
            .I(\c0.n6_adj_4510_cascade_ ));
    InMux I__8437 (
            .O(N__51465),
            .I(N__51459));
    InMux I__8436 (
            .O(N__51464),
            .I(N__51459));
    LocalMux I__8435 (
            .O(N__51459),
            .I(\c0.data_out_frame_0_3 ));
    InMux I__8434 (
            .O(N__51456),
            .I(\c0.n30204 ));
    InMux I__8433 (
            .O(N__51453),
            .I(\c0.n30205 ));
    InMux I__8432 (
            .O(N__51450),
            .I(\c0.n30206 ));
    InMux I__8431 (
            .O(N__51447),
            .I(\c0.n30207 ));
    InMux I__8430 (
            .O(N__51444),
            .I(\c0.n30208 ));
    CEMux I__8429 (
            .O(N__51441),
            .I(N__51438));
    LocalMux I__8428 (
            .O(N__51438),
            .I(N__51434));
    InMux I__8427 (
            .O(N__51437),
            .I(N__51431));
    Span4Mux_v I__8426 (
            .O(N__51434),
            .I(N__51428));
    LocalMux I__8425 (
            .O(N__51431),
            .I(N__51425));
    Span4Mux_h I__8424 (
            .O(N__51428),
            .I(N__51420));
    Span4Mux_v I__8423 (
            .O(N__51425),
            .I(N__51420));
    Span4Mux_h I__8422 (
            .O(N__51420),
            .I(N__51417));
    Odrv4 I__8421 (
            .O(N__51417),
            .I(\c0.n19388 ));
    SRMux I__8420 (
            .O(N__51414),
            .I(N__51411));
    LocalMux I__8419 (
            .O(N__51411),
            .I(N__51408));
    Span4Mux_h I__8418 (
            .O(N__51408),
            .I(N__51405));
    Span4Mux_v I__8417 (
            .O(N__51405),
            .I(N__51402));
    Odrv4 I__8416 (
            .O(N__51402),
            .I(\c0.n29678 ));
    CascadeMux I__8415 (
            .O(N__51399),
            .I(data_out_frame_29__7__N_1482_cascade_));
    InMux I__8414 (
            .O(N__51396),
            .I(N__51393));
    LocalMux I__8413 (
            .O(N__51393),
            .I(N__51390));
    Span4Mux_v I__8412 (
            .O(N__51390),
            .I(N__51387));
    Span4Mux_h I__8411 (
            .O(N__51387),
            .I(N__51384));
    Odrv4 I__8410 (
            .O(N__51384),
            .I(n10_adj_4805));
    InMux I__8409 (
            .O(N__51381),
            .I(N__51378));
    LocalMux I__8408 (
            .O(N__51378),
            .I(N__51374));
    InMux I__8407 (
            .O(N__51377),
            .I(N__51371));
    Span4Mux_v I__8406 (
            .O(N__51374),
            .I(N__51367));
    LocalMux I__8405 (
            .O(N__51371),
            .I(N__51364));
    InMux I__8404 (
            .O(N__51370),
            .I(N__51361));
    Span4Mux_h I__8403 (
            .O(N__51367),
            .I(N__51358));
    Span4Mux_h I__8402 (
            .O(N__51364),
            .I(N__51355));
    LocalMux I__8401 (
            .O(N__51361),
            .I(\c0.n17961 ));
    Odrv4 I__8400 (
            .O(N__51358),
            .I(\c0.n17961 ));
    Odrv4 I__8399 (
            .O(N__51355),
            .I(\c0.n17961 ));
    InMux I__8398 (
            .O(N__51348),
            .I(N__51344));
    InMux I__8397 (
            .O(N__51347),
            .I(N__51341));
    LocalMux I__8396 (
            .O(N__51344),
            .I(N__51335));
    LocalMux I__8395 (
            .O(N__51341),
            .I(N__51335));
    CascadeMux I__8394 (
            .O(N__51340),
            .I(N__51332));
    Span4Mux_h I__8393 (
            .O(N__51335),
            .I(N__51329));
    InMux I__8392 (
            .O(N__51332),
            .I(N__51326));
    Odrv4 I__8391 (
            .O(N__51329),
            .I(\quad_counter0.n2707 ));
    LocalMux I__8390 (
            .O(N__51326),
            .I(\quad_counter0.n2707 ));
    InMux I__8389 (
            .O(N__51321),
            .I(\quad_counter0.n30296 ));
    InMux I__8388 (
            .O(N__51318),
            .I(N__51314));
    InMux I__8387 (
            .O(N__51317),
            .I(N__51311));
    LocalMux I__8386 (
            .O(N__51314),
            .I(N__51306));
    LocalMux I__8385 (
            .O(N__51311),
            .I(N__51306));
    Span4Mux_h I__8384 (
            .O(N__51306),
            .I(N__51302));
    InMux I__8383 (
            .O(N__51305),
            .I(N__51299));
    Odrv4 I__8382 (
            .O(N__51302),
            .I(\quad_counter0.n2706 ));
    LocalMux I__8381 (
            .O(N__51299),
            .I(\quad_counter0.n2706 ));
    InMux I__8380 (
            .O(N__51294),
            .I(\quad_counter0.n30297 ));
    InMux I__8379 (
            .O(N__51291),
            .I(\quad_counter0.n30298 ));
    InMux I__8378 (
            .O(N__51288),
            .I(N__51284));
    InMux I__8377 (
            .O(N__51287),
            .I(N__51281));
    LocalMux I__8376 (
            .O(N__51284),
            .I(N__51276));
    LocalMux I__8375 (
            .O(N__51281),
            .I(N__51276));
    Span4Mux_h I__8374 (
            .O(N__51276),
            .I(N__51272));
    InMux I__8373 (
            .O(N__51275),
            .I(N__51269));
    Odrv4 I__8372 (
            .O(N__51272),
            .I(\quad_counter0.n2705 ));
    LocalMux I__8371 (
            .O(N__51269),
            .I(\quad_counter0.n2705 ));
    InMux I__8370 (
            .O(N__51264),
            .I(N__51261));
    LocalMux I__8369 (
            .O(N__51261),
            .I(N__51258));
    Odrv12 I__8368 (
            .O(N__51258),
            .I(\quad_counter0.n12_adj_4396 ));
    CascadeMux I__8367 (
            .O(N__51255),
            .I(\quad_counter0.n2441_cascade_ ));
    InMux I__8366 (
            .O(N__51252),
            .I(N__51249));
    LocalMux I__8365 (
            .O(N__51249),
            .I(N__51245));
    InMux I__8364 (
            .O(N__51248),
            .I(N__51242));
    Span4Mux_h I__8363 (
            .O(N__51245),
            .I(N__51239));
    LocalMux I__8362 (
            .O(N__51242),
            .I(r_Tx_Data_6));
    Odrv4 I__8361 (
            .O(N__51239),
            .I(r_Tx_Data_6));
    InMux I__8360 (
            .O(N__51234),
            .I(N__51231));
    LocalMux I__8359 (
            .O(N__51231),
            .I(N__51227));
    CascadeMux I__8358 (
            .O(N__51230),
            .I(N__51224));
    Span4Mux_h I__8357 (
            .O(N__51227),
            .I(N__51221));
    InMux I__8356 (
            .O(N__51224),
            .I(N__51218));
    Odrv4 I__8355 (
            .O(N__51221),
            .I(\c0.tx_transmit_N_3651 ));
    LocalMux I__8354 (
            .O(N__51218),
            .I(\c0.tx_transmit_N_3651 ));
    InMux I__8353 (
            .O(N__51213),
            .I(\c0.n30202 ));
    InMux I__8352 (
            .O(N__51210),
            .I(\c0.n30203 ));
    InMux I__8351 (
            .O(N__51207),
            .I(\quad_counter0.n30287 ));
    InMux I__8350 (
            .O(N__51204),
            .I(N__51200));
    InMux I__8349 (
            .O(N__51203),
            .I(N__51197));
    LocalMux I__8348 (
            .O(N__51200),
            .I(N__51192));
    LocalMux I__8347 (
            .O(N__51197),
            .I(N__51192));
    Span4Mux_h I__8346 (
            .O(N__51192),
            .I(N__51188));
    InMux I__8345 (
            .O(N__51191),
            .I(N__51185));
    Odrv4 I__8344 (
            .O(N__51188),
            .I(\quad_counter0.n2715 ));
    LocalMux I__8343 (
            .O(N__51185),
            .I(\quad_counter0.n2715 ));
    InMux I__8342 (
            .O(N__51180),
            .I(\quad_counter0.n30288 ));
    InMux I__8341 (
            .O(N__51177),
            .I(N__51173));
    InMux I__8340 (
            .O(N__51176),
            .I(N__51170));
    LocalMux I__8339 (
            .O(N__51173),
            .I(N__51165));
    LocalMux I__8338 (
            .O(N__51170),
            .I(N__51165));
    Span4Mux_h I__8337 (
            .O(N__51165),
            .I(N__51161));
    InMux I__8336 (
            .O(N__51164),
            .I(N__51158));
    Odrv4 I__8335 (
            .O(N__51161),
            .I(\quad_counter0.n2714 ));
    LocalMux I__8334 (
            .O(N__51158),
            .I(\quad_counter0.n2714 ));
    InMux I__8333 (
            .O(N__51153),
            .I(\quad_counter0.n30289 ));
    InMux I__8332 (
            .O(N__51150),
            .I(N__51146));
    InMux I__8331 (
            .O(N__51149),
            .I(N__51143));
    LocalMux I__8330 (
            .O(N__51146),
            .I(N__51138));
    LocalMux I__8329 (
            .O(N__51143),
            .I(N__51138));
    Span4Mux_h I__8328 (
            .O(N__51138),
            .I(N__51134));
    InMux I__8327 (
            .O(N__51137),
            .I(N__51131));
    Odrv4 I__8326 (
            .O(N__51134),
            .I(\quad_counter0.n2713 ));
    LocalMux I__8325 (
            .O(N__51131),
            .I(\quad_counter0.n2713 ));
    InMux I__8324 (
            .O(N__51126),
            .I(\quad_counter0.n30290 ));
    InMux I__8323 (
            .O(N__51123),
            .I(N__51119));
    InMux I__8322 (
            .O(N__51122),
            .I(N__51116));
    LocalMux I__8321 (
            .O(N__51119),
            .I(N__51111));
    LocalMux I__8320 (
            .O(N__51116),
            .I(N__51111));
    Span4Mux_h I__8319 (
            .O(N__51111),
            .I(N__51107));
    InMux I__8318 (
            .O(N__51110),
            .I(N__51104));
    Odrv4 I__8317 (
            .O(N__51107),
            .I(\quad_counter0.n2712 ));
    LocalMux I__8316 (
            .O(N__51104),
            .I(\quad_counter0.n2712 ));
    InMux I__8315 (
            .O(N__51099),
            .I(\quad_counter0.n30291 ));
    InMux I__8314 (
            .O(N__51096),
            .I(N__51092));
    InMux I__8313 (
            .O(N__51095),
            .I(N__51089));
    LocalMux I__8312 (
            .O(N__51092),
            .I(N__51083));
    LocalMux I__8311 (
            .O(N__51089),
            .I(N__51083));
    CascadeMux I__8310 (
            .O(N__51088),
            .I(N__51080));
    Span4Mux_h I__8309 (
            .O(N__51083),
            .I(N__51077));
    InMux I__8308 (
            .O(N__51080),
            .I(N__51074));
    Odrv4 I__8307 (
            .O(N__51077),
            .I(\quad_counter0.n2711 ));
    LocalMux I__8306 (
            .O(N__51074),
            .I(\quad_counter0.n2711 ));
    InMux I__8305 (
            .O(N__51069),
            .I(bfn_14_12_0_));
    InMux I__8304 (
            .O(N__51066),
            .I(N__51062));
    InMux I__8303 (
            .O(N__51065),
            .I(N__51059));
    LocalMux I__8302 (
            .O(N__51062),
            .I(N__51054));
    LocalMux I__8301 (
            .O(N__51059),
            .I(N__51054));
    Span4Mux_h I__8300 (
            .O(N__51054),
            .I(N__51050));
    InMux I__8299 (
            .O(N__51053),
            .I(N__51047));
    Odrv4 I__8298 (
            .O(N__51050),
            .I(\quad_counter0.n2710 ));
    LocalMux I__8297 (
            .O(N__51047),
            .I(\quad_counter0.n2710 ));
    InMux I__8296 (
            .O(N__51042),
            .I(\quad_counter0.n30293 ));
    InMux I__8295 (
            .O(N__51039),
            .I(N__51035));
    InMux I__8294 (
            .O(N__51038),
            .I(N__51032));
    LocalMux I__8293 (
            .O(N__51035),
            .I(N__51027));
    LocalMux I__8292 (
            .O(N__51032),
            .I(N__51027));
    Span4Mux_v I__8291 (
            .O(N__51027),
            .I(N__51023));
    InMux I__8290 (
            .O(N__51026),
            .I(N__51020));
    Odrv4 I__8289 (
            .O(N__51023),
            .I(\quad_counter0.n2709 ));
    LocalMux I__8288 (
            .O(N__51020),
            .I(\quad_counter0.n2709 ));
    InMux I__8287 (
            .O(N__51015),
            .I(\quad_counter0.n30294 ));
    InMux I__8286 (
            .O(N__51012),
            .I(N__51008));
    InMux I__8285 (
            .O(N__51011),
            .I(N__51005));
    LocalMux I__8284 (
            .O(N__51008),
            .I(N__51000));
    LocalMux I__8283 (
            .O(N__51005),
            .I(N__51000));
    Span4Mux_v I__8282 (
            .O(N__51000),
            .I(N__50996));
    InMux I__8281 (
            .O(N__50999),
            .I(N__50993));
    Odrv4 I__8280 (
            .O(N__50996),
            .I(\quad_counter0.n2708 ));
    LocalMux I__8279 (
            .O(N__50993),
            .I(\quad_counter0.n2708 ));
    InMux I__8278 (
            .O(N__50988),
            .I(\quad_counter0.n30295 ));
    InMux I__8277 (
            .O(N__50985),
            .I(N__50982));
    LocalMux I__8276 (
            .O(N__50982),
            .I(\quad_counter0.n34759 ));
    InMux I__8275 (
            .O(N__50979),
            .I(N__50976));
    LocalMux I__8274 (
            .O(N__50976),
            .I(\quad_counter0.n12 ));
    InMux I__8273 (
            .O(N__50973),
            .I(N__50970));
    LocalMux I__8272 (
            .O(N__50970),
            .I(\quad_counter0.n30_adj_4371 ));
    InMux I__8271 (
            .O(N__50967),
            .I(N__50964));
    LocalMux I__8270 (
            .O(N__50964),
            .I(\quad_counter0.n29_adj_4373 ));
    CascadeMux I__8269 (
            .O(N__50961),
            .I(N__50958));
    InMux I__8268 (
            .O(N__50958),
            .I(N__50955));
    LocalMux I__8267 (
            .O(N__50955),
            .I(\quad_counter0.n28_adj_4372 ));
    InMux I__8266 (
            .O(N__50952),
            .I(N__50949));
    LocalMux I__8265 (
            .O(N__50949),
            .I(\quad_counter0.n27_adj_4374 ));
    InMux I__8264 (
            .O(N__50946),
            .I(N__50942));
    InMux I__8263 (
            .O(N__50945),
            .I(N__50939));
    LocalMux I__8262 (
            .O(N__50942),
            .I(N__50934));
    LocalMux I__8261 (
            .O(N__50939),
            .I(N__50934));
    Span4Mux_h I__8260 (
            .O(N__50934),
            .I(N__50930));
    InMux I__8259 (
            .O(N__50933),
            .I(N__50927));
    Odrv4 I__8258 (
            .O(N__50930),
            .I(\quad_counter0.n2719 ));
    LocalMux I__8257 (
            .O(N__50927),
            .I(\quad_counter0.n2719 ));
    InMux I__8256 (
            .O(N__50922),
            .I(bfn_14_11_0_));
    InMux I__8255 (
            .O(N__50919),
            .I(N__50915));
    InMux I__8254 (
            .O(N__50918),
            .I(N__50912));
    LocalMux I__8253 (
            .O(N__50915),
            .I(N__50907));
    LocalMux I__8252 (
            .O(N__50912),
            .I(N__50907));
    Span4Mux_h I__8251 (
            .O(N__50907),
            .I(N__50903));
    InMux I__8250 (
            .O(N__50906),
            .I(N__50900));
    Odrv4 I__8249 (
            .O(N__50903),
            .I(\quad_counter0.n2718 ));
    LocalMux I__8248 (
            .O(N__50900),
            .I(\quad_counter0.n2718 ));
    InMux I__8247 (
            .O(N__50895),
            .I(\quad_counter0.n30285 ));
    InMux I__8246 (
            .O(N__50892),
            .I(N__50888));
    InMux I__8245 (
            .O(N__50891),
            .I(N__50885));
    LocalMux I__8244 (
            .O(N__50888),
            .I(N__50880));
    LocalMux I__8243 (
            .O(N__50885),
            .I(N__50880));
    Span4Mux_v I__8242 (
            .O(N__50880),
            .I(N__50876));
    InMux I__8241 (
            .O(N__50879),
            .I(N__50873));
    Odrv4 I__8240 (
            .O(N__50876),
            .I(\quad_counter0.n2717 ));
    LocalMux I__8239 (
            .O(N__50873),
            .I(\quad_counter0.n2717 ));
    InMux I__8238 (
            .O(N__50868),
            .I(\quad_counter0.n30286 ));
    InMux I__8237 (
            .O(N__50865),
            .I(N__50861));
    InMux I__8236 (
            .O(N__50864),
            .I(N__50858));
    LocalMux I__8235 (
            .O(N__50861),
            .I(N__50853));
    LocalMux I__8234 (
            .O(N__50858),
            .I(N__50853));
    Span4Mux_v I__8233 (
            .O(N__50853),
            .I(N__50849));
    InMux I__8232 (
            .O(N__50852),
            .I(N__50846));
    Odrv4 I__8231 (
            .O(N__50849),
            .I(\quad_counter0.n2716 ));
    LocalMux I__8230 (
            .O(N__50846),
            .I(\quad_counter0.n2716 ));
    CascadeMux I__8229 (
            .O(N__50841),
            .I(\quad_counter0.n2014_cascade_ ));
    InMux I__8228 (
            .O(N__50838),
            .I(N__50835));
    LocalMux I__8227 (
            .O(N__50835),
            .I(\quad_counter0.n28371 ));
    InMux I__8226 (
            .O(N__50832),
            .I(N__50828));
    InMux I__8225 (
            .O(N__50831),
            .I(N__50825));
    LocalMux I__8224 (
            .O(N__50828),
            .I(\quad_counter0.n2012 ));
    LocalMux I__8223 (
            .O(N__50825),
            .I(\quad_counter0.n2012 ));
    CascadeMux I__8222 (
            .O(N__50820),
            .I(N__50816));
    CascadeMux I__8221 (
            .O(N__50819),
            .I(N__50813));
    InMux I__8220 (
            .O(N__50816),
            .I(N__50809));
    InMux I__8219 (
            .O(N__50813),
            .I(N__50804));
    InMux I__8218 (
            .O(N__50812),
            .I(N__50804));
    LocalMux I__8217 (
            .O(N__50809),
            .I(\quad_counter0.n2013 ));
    LocalMux I__8216 (
            .O(N__50804),
            .I(\quad_counter0.n2013 ));
    CascadeMux I__8215 (
            .O(N__50799),
            .I(\quad_counter0.n10_adj_4378_cascade_ ));
    CascadeMux I__8214 (
            .O(N__50796),
            .I(N__50792));
    InMux I__8213 (
            .O(N__50795),
            .I(N__50789));
    InMux I__8212 (
            .O(N__50792),
            .I(N__50786));
    LocalMux I__8211 (
            .O(N__50789),
            .I(\quad_counter0.n2019 ));
    LocalMux I__8210 (
            .O(N__50786),
            .I(\quad_counter0.n2019 ));
    CascadeMux I__8209 (
            .O(N__50781),
            .I(\quad_counter0.n2045_cascade_ ));
    InMux I__8208 (
            .O(N__50778),
            .I(N__50775));
    LocalMux I__8207 (
            .O(N__50775),
            .I(N__50772));
    Odrv4 I__8206 (
            .O(N__50772),
            .I(\quad_counter0.n2086 ));
    InMux I__8205 (
            .O(N__50769),
            .I(N__50766));
    LocalMux I__8204 (
            .O(N__50766),
            .I(\quad_counter0.n9_adj_4379 ));
    CascadeMux I__8203 (
            .O(N__50763),
            .I(\quad_counter0.n30_cascade_ ));
    CascadeMux I__8202 (
            .O(N__50760),
            .I(\quad_counter0.n28291_cascade_ ));
    CascadeMux I__8201 (
            .O(N__50757),
            .I(\quad_counter0.n10_cascade_ ));
    InMux I__8200 (
            .O(N__50754),
            .I(N__50751));
    LocalMux I__8199 (
            .O(N__50751),
            .I(\quad_counter0.n21 ));
    InMux I__8198 (
            .O(N__50748),
            .I(\quad_counter0.n30226 ));
    InMux I__8197 (
            .O(N__50745),
            .I(\quad_counter0.n30227 ));
    InMux I__8196 (
            .O(N__50742),
            .I(\quad_counter0.n30228 ));
    InMux I__8195 (
            .O(N__50739),
            .I(bfn_14_6_0_));
    InMux I__8194 (
            .O(N__50736),
            .I(N__50733));
    LocalMux I__8193 (
            .O(N__50733),
            .I(\quad_counter0.n2087 ));
    CascadeMux I__8192 (
            .O(N__50730),
            .I(\quad_counter0.n2119_cascade_ ));
    InMux I__8191 (
            .O(N__50727),
            .I(N__50724));
    LocalMux I__8190 (
            .O(N__50724),
            .I(\quad_counter0.n1985 ));
    CascadeMux I__8189 (
            .O(N__50721),
            .I(N__50718));
    InMux I__8188 (
            .O(N__50718),
            .I(N__50715));
    LocalMux I__8187 (
            .O(N__50715),
            .I(N__50711));
    CascadeMux I__8186 (
            .O(N__50714),
            .I(N__50708));
    Span4Mux_v I__8185 (
            .O(N__50711),
            .I(N__50704));
    InMux I__8184 (
            .O(N__50708),
            .I(N__50701));
    InMux I__8183 (
            .O(N__50707),
            .I(N__50698));
    Odrv4 I__8182 (
            .O(N__50704),
            .I(\quad_counter0.n1918 ));
    LocalMux I__8181 (
            .O(N__50701),
            .I(\quad_counter0.n1918 ));
    LocalMux I__8180 (
            .O(N__50698),
            .I(\quad_counter0.n1918 ));
    InMux I__8179 (
            .O(N__50691),
            .I(N__50688));
    LocalMux I__8178 (
            .O(N__50688),
            .I(N__50685));
    Odrv4 I__8177 (
            .O(N__50685),
            .I(\quad_counter0.n2080 ));
    InMux I__8176 (
            .O(N__50682),
            .I(N__50679));
    LocalMux I__8175 (
            .O(N__50679),
            .I(\quad_counter0.n1982 ));
    CascadeMux I__8174 (
            .O(N__50676),
            .I(N__50673));
    InMux I__8173 (
            .O(N__50673),
            .I(N__50669));
    CascadeMux I__8172 (
            .O(N__50672),
            .I(N__50666));
    LocalMux I__8171 (
            .O(N__50669),
            .I(N__50662));
    InMux I__8170 (
            .O(N__50666),
            .I(N__50659));
    InMux I__8169 (
            .O(N__50665),
            .I(N__50656));
    Odrv4 I__8168 (
            .O(N__50662),
            .I(\quad_counter0.n1915 ));
    LocalMux I__8167 (
            .O(N__50659),
            .I(\quad_counter0.n1915 ));
    LocalMux I__8166 (
            .O(N__50656),
            .I(\quad_counter0.n1915 ));
    CascadeMux I__8165 (
            .O(N__50649),
            .I(N__50646));
    InMux I__8164 (
            .O(N__50646),
            .I(N__50642));
    InMux I__8163 (
            .O(N__50645),
            .I(N__50639));
    LocalMux I__8162 (
            .O(N__50642),
            .I(\c0.data_in_frame_23_0 ));
    LocalMux I__8161 (
            .O(N__50639),
            .I(\c0.data_in_frame_23_0 ));
    InMux I__8160 (
            .O(N__50634),
            .I(bfn_14_5_0_));
    InMux I__8159 (
            .O(N__50631),
            .I(\quad_counter0.n30222 ));
    InMux I__8158 (
            .O(N__50628),
            .I(\quad_counter0.n30223 ));
    InMux I__8157 (
            .O(N__50625),
            .I(\quad_counter0.n30224 ));
    InMux I__8156 (
            .O(N__50622),
            .I(\quad_counter0.n30225 ));
    CascadeMux I__8155 (
            .O(N__50619),
            .I(\c0.n33545_cascade_ ));
    CascadeMux I__8154 (
            .O(N__50616),
            .I(\c0.n35505_cascade_ ));
    CascadeMux I__8153 (
            .O(N__50613),
            .I(N__50609));
    InMux I__8152 (
            .O(N__50612),
            .I(N__50605));
    InMux I__8151 (
            .O(N__50609),
            .I(N__50602));
    InMux I__8150 (
            .O(N__50608),
            .I(N__50599));
    LocalMux I__8149 (
            .O(N__50605),
            .I(N__50595));
    LocalMux I__8148 (
            .O(N__50602),
            .I(N__50590));
    LocalMux I__8147 (
            .O(N__50599),
            .I(N__50590));
    InMux I__8146 (
            .O(N__50598),
            .I(N__50587));
    Odrv4 I__8145 (
            .O(N__50595),
            .I(\c0.data_in_frame_18_7 ));
    Odrv4 I__8144 (
            .O(N__50590),
            .I(\c0.data_in_frame_18_7 ));
    LocalMux I__8143 (
            .O(N__50587),
            .I(\c0.data_in_frame_18_7 ));
    CascadeMux I__8142 (
            .O(N__50580),
            .I(N__50574));
    InMux I__8141 (
            .O(N__50579),
            .I(N__50571));
    InMux I__8140 (
            .O(N__50578),
            .I(N__50568));
    InMux I__8139 (
            .O(N__50577),
            .I(N__50565));
    InMux I__8138 (
            .O(N__50574),
            .I(N__50562));
    LocalMux I__8137 (
            .O(N__50571),
            .I(N__50559));
    LocalMux I__8136 (
            .O(N__50568),
            .I(N__50556));
    LocalMux I__8135 (
            .O(N__50565),
            .I(N__50553));
    LocalMux I__8134 (
            .O(N__50562),
            .I(\c0.data_in_frame_18_6 ));
    Odrv12 I__8133 (
            .O(N__50559),
            .I(\c0.data_in_frame_18_6 ));
    Odrv4 I__8132 (
            .O(N__50556),
            .I(\c0.data_in_frame_18_6 ));
    Odrv12 I__8131 (
            .O(N__50553),
            .I(\c0.data_in_frame_18_6 ));
    CascadeMux I__8130 (
            .O(N__50544),
            .I(\c0.n33852_cascade_ ));
    InMux I__8129 (
            .O(N__50541),
            .I(N__50537));
    InMux I__8128 (
            .O(N__50540),
            .I(N__50534));
    LocalMux I__8127 (
            .O(N__50537),
            .I(\c0.n33942 ));
    LocalMux I__8126 (
            .O(N__50534),
            .I(\c0.n33942 ));
    InMux I__8125 (
            .O(N__50529),
            .I(N__50526));
    LocalMux I__8124 (
            .O(N__50526),
            .I(\c0.n10_adj_4575 ));
    InMux I__8123 (
            .O(N__50523),
            .I(N__50518));
    InMux I__8122 (
            .O(N__50522),
            .I(N__50515));
    InMux I__8121 (
            .O(N__50521),
            .I(N__50512));
    LocalMux I__8120 (
            .O(N__50518),
            .I(N__50506));
    LocalMux I__8119 (
            .O(N__50515),
            .I(N__50506));
    LocalMux I__8118 (
            .O(N__50512),
            .I(N__50503));
    InMux I__8117 (
            .O(N__50511),
            .I(N__50500));
    Span4Mux_v I__8116 (
            .O(N__50506),
            .I(N__50497));
    Span4Mux_v I__8115 (
            .O(N__50503),
            .I(N__50492));
    LocalMux I__8114 (
            .O(N__50500),
            .I(N__50492));
    Odrv4 I__8113 (
            .O(N__50497),
            .I(\c0.n33647 ));
    Odrv4 I__8112 (
            .O(N__50492),
            .I(\c0.n33647 ));
    CascadeMux I__8111 (
            .O(N__50487),
            .I(\c0.n10_adj_4575_cascade_ ));
    InMux I__8110 (
            .O(N__50484),
            .I(N__50478));
    InMux I__8109 (
            .O(N__50483),
            .I(N__50473));
    InMux I__8108 (
            .O(N__50482),
            .I(N__50473));
    InMux I__8107 (
            .O(N__50481),
            .I(N__50470));
    LocalMux I__8106 (
            .O(N__50478),
            .I(N__50462));
    LocalMux I__8105 (
            .O(N__50473),
            .I(N__50462));
    LocalMux I__8104 (
            .O(N__50470),
            .I(N__50462));
    InMux I__8103 (
            .O(N__50469),
            .I(N__50459));
    Span4Mux_v I__8102 (
            .O(N__50462),
            .I(N__50454));
    LocalMux I__8101 (
            .O(N__50459),
            .I(N__50454));
    Odrv4 I__8100 (
            .O(N__50454),
            .I(\c0.n32302 ));
    CascadeMux I__8099 (
            .O(N__50451),
            .I(\c0.n32390_cascade_ ));
    InMux I__8098 (
            .O(N__50448),
            .I(N__50445));
    LocalMux I__8097 (
            .O(N__50445),
            .I(N__50442));
    Odrv12 I__8096 (
            .O(N__50442),
            .I(\c0.n18_adj_4563 ));
    CascadeMux I__8095 (
            .O(N__50439),
            .I(N__50435));
    CascadeMux I__8094 (
            .O(N__50438),
            .I(N__50431));
    InMux I__8093 (
            .O(N__50435),
            .I(N__50421));
    InMux I__8092 (
            .O(N__50434),
            .I(N__50421));
    InMux I__8091 (
            .O(N__50431),
            .I(N__50421));
    InMux I__8090 (
            .O(N__50430),
            .I(N__50421));
    LocalMux I__8089 (
            .O(N__50421),
            .I(\c0.data_in_frame_19_4 ));
    InMux I__8088 (
            .O(N__50418),
            .I(N__50414));
    InMux I__8087 (
            .O(N__50417),
            .I(N__50411));
    LocalMux I__8086 (
            .O(N__50414),
            .I(N__50408));
    LocalMux I__8085 (
            .O(N__50411),
            .I(N__50405));
    Span12Mux_s8_v I__8084 (
            .O(N__50408),
            .I(N__50402));
    Span4Mux_h I__8083 (
            .O(N__50405),
            .I(N__50399));
    Odrv12 I__8082 (
            .O(N__50402),
            .I(\c0.n18582 ));
    Odrv4 I__8081 (
            .O(N__50399),
            .I(\c0.n18582 ));
    CascadeMux I__8080 (
            .O(N__50394),
            .I(N__50390));
    InMux I__8079 (
            .O(N__50393),
            .I(N__50385));
    InMux I__8078 (
            .O(N__50390),
            .I(N__50380));
    InMux I__8077 (
            .O(N__50389),
            .I(N__50380));
    CascadeMux I__8076 (
            .O(N__50388),
            .I(N__50377));
    LocalMux I__8075 (
            .O(N__50385),
            .I(N__50372));
    LocalMux I__8074 (
            .O(N__50380),
            .I(N__50369));
    InMux I__8073 (
            .O(N__50377),
            .I(N__50366));
    InMux I__8072 (
            .O(N__50376),
            .I(N__50361));
    InMux I__8071 (
            .O(N__50375),
            .I(N__50361));
    Span12Mux_s8_v I__8070 (
            .O(N__50372),
            .I(N__50358));
    Span4Mux_h I__8069 (
            .O(N__50369),
            .I(N__50355));
    LocalMux I__8068 (
            .O(N__50366),
            .I(N__50350));
    LocalMux I__8067 (
            .O(N__50361),
            .I(N__50350));
    Odrv12 I__8066 (
            .O(N__50358),
            .I(\c0.data_in_frame_17_1 ));
    Odrv4 I__8065 (
            .O(N__50355),
            .I(\c0.data_in_frame_17_1 ));
    Odrv4 I__8064 (
            .O(N__50350),
            .I(\c0.data_in_frame_17_1 ));
    InMux I__8063 (
            .O(N__50343),
            .I(N__50339));
    InMux I__8062 (
            .O(N__50342),
            .I(N__50334));
    LocalMux I__8061 (
            .O(N__50339),
            .I(N__50331));
    InMux I__8060 (
            .O(N__50338),
            .I(N__50326));
    InMux I__8059 (
            .O(N__50337),
            .I(N__50326));
    LocalMux I__8058 (
            .O(N__50334),
            .I(N__50323));
    Span4Mux_v I__8057 (
            .O(N__50331),
            .I(N__50320));
    LocalMux I__8056 (
            .O(N__50326),
            .I(\c0.data_in_frame_12_3 ));
    Odrv4 I__8055 (
            .O(N__50323),
            .I(\c0.data_in_frame_12_3 ));
    Odrv4 I__8054 (
            .O(N__50320),
            .I(\c0.data_in_frame_12_3 ));
    InMux I__8053 (
            .O(N__50313),
            .I(N__50310));
    LocalMux I__8052 (
            .O(N__50310),
            .I(N__50307));
    Span4Mux_h I__8051 (
            .O(N__50307),
            .I(N__50304));
    Odrv4 I__8050 (
            .O(N__50304),
            .I(\c0.n33545 ));
    InMux I__8049 (
            .O(N__50301),
            .I(N__50298));
    LocalMux I__8048 (
            .O(N__50298),
            .I(N__50294));
    InMux I__8047 (
            .O(N__50297),
            .I(N__50291));
    Span4Mux_h I__8046 (
            .O(N__50294),
            .I(N__50288));
    LocalMux I__8045 (
            .O(N__50291),
            .I(\c0.data_in_frame_10_3 ));
    Odrv4 I__8044 (
            .O(N__50288),
            .I(\c0.data_in_frame_10_3 ));
    CascadeMux I__8043 (
            .O(N__50283),
            .I(N__50280));
    InMux I__8042 (
            .O(N__50280),
            .I(N__50277));
    LocalMux I__8041 (
            .O(N__50277),
            .I(N__50274));
    Span4Mux_h I__8040 (
            .O(N__50274),
            .I(N__50271));
    Odrv4 I__8039 (
            .O(N__50271),
            .I(\c0.n5996 ));
    InMux I__8038 (
            .O(N__50268),
            .I(N__50265));
    LocalMux I__8037 (
            .O(N__50265),
            .I(N__50262));
    Odrv4 I__8036 (
            .O(N__50262),
            .I(\c0.n18290 ));
    CascadeMux I__8035 (
            .O(N__50259),
            .I(N__50256));
    InMux I__8034 (
            .O(N__50256),
            .I(N__50253));
    LocalMux I__8033 (
            .O(N__50253),
            .I(N__50247));
    InMux I__8032 (
            .O(N__50252),
            .I(N__50242));
    InMux I__8031 (
            .O(N__50251),
            .I(N__50242));
    CascadeMux I__8030 (
            .O(N__50250),
            .I(N__50239));
    Span4Mux_h I__8029 (
            .O(N__50247),
            .I(N__50234));
    LocalMux I__8028 (
            .O(N__50242),
            .I(N__50234));
    InMux I__8027 (
            .O(N__50239),
            .I(N__50230));
    Span4Mux_h I__8026 (
            .O(N__50234),
            .I(N__50227));
    InMux I__8025 (
            .O(N__50233),
            .I(N__50224));
    LocalMux I__8024 (
            .O(N__50230),
            .I(\c0.data_in_frame_12_6 ));
    Odrv4 I__8023 (
            .O(N__50227),
            .I(\c0.data_in_frame_12_6 ));
    LocalMux I__8022 (
            .O(N__50224),
            .I(\c0.data_in_frame_12_6 ));
    InMux I__8021 (
            .O(N__50217),
            .I(N__50213));
    InMux I__8020 (
            .O(N__50216),
            .I(N__50210));
    LocalMux I__8019 (
            .O(N__50213),
            .I(N__50207));
    LocalMux I__8018 (
            .O(N__50210),
            .I(N__50204));
    Odrv12 I__8017 (
            .O(N__50207),
            .I(\c0.n18147 ));
    Odrv4 I__8016 (
            .O(N__50204),
            .I(\c0.n18147 ));
    InMux I__8015 (
            .O(N__50199),
            .I(N__50194));
    InMux I__8014 (
            .O(N__50198),
            .I(N__50191));
    InMux I__8013 (
            .O(N__50197),
            .I(N__50187));
    LocalMux I__8012 (
            .O(N__50194),
            .I(N__50182));
    LocalMux I__8011 (
            .O(N__50191),
            .I(N__50182));
    InMux I__8010 (
            .O(N__50190),
            .I(N__50179));
    LocalMux I__8009 (
            .O(N__50187),
            .I(N__50176));
    Span4Mux_h I__8008 (
            .O(N__50182),
            .I(N__50173));
    LocalMux I__8007 (
            .O(N__50179),
            .I(\c0.data_in_frame_12_0 ));
    Odrv12 I__8006 (
            .O(N__50176),
            .I(\c0.data_in_frame_12_0 ));
    Odrv4 I__8005 (
            .O(N__50173),
            .I(\c0.data_in_frame_12_0 ));
    InMux I__8004 (
            .O(N__50166),
            .I(N__50163));
    LocalMux I__8003 (
            .O(N__50163),
            .I(N__50160));
    Span4Mux_h I__8002 (
            .O(N__50160),
            .I(N__50157));
    Span4Mux_h I__8001 (
            .O(N__50157),
            .I(N__50154));
    Odrv4 I__8000 (
            .O(N__50154),
            .I(\c0.n33705 ));
    InMux I__7999 (
            .O(N__50151),
            .I(N__50148));
    LocalMux I__7998 (
            .O(N__50148),
            .I(N__50145));
    Span4Mux_h I__7997 (
            .O(N__50145),
            .I(N__50142));
    Odrv4 I__7996 (
            .O(N__50142),
            .I(\c0.n10_adj_4744 ));
    InMux I__7995 (
            .O(N__50139),
            .I(N__50134));
    InMux I__7994 (
            .O(N__50138),
            .I(N__50129));
    InMux I__7993 (
            .O(N__50137),
            .I(N__50129));
    LocalMux I__7992 (
            .O(N__50134),
            .I(N__50121));
    LocalMux I__7991 (
            .O(N__50129),
            .I(N__50121));
    CascadeMux I__7990 (
            .O(N__50128),
            .I(N__50118));
    CascadeMux I__7989 (
            .O(N__50127),
            .I(N__50115));
    InMux I__7988 (
            .O(N__50126),
            .I(N__50112));
    Span4Mux_h I__7987 (
            .O(N__50121),
            .I(N__50109));
    InMux I__7986 (
            .O(N__50118),
            .I(N__50104));
    InMux I__7985 (
            .O(N__50115),
            .I(N__50104));
    LocalMux I__7984 (
            .O(N__50112),
            .I(\c0.data_in_frame_8_3 ));
    Odrv4 I__7983 (
            .O(N__50109),
            .I(\c0.data_in_frame_8_3 ));
    LocalMux I__7982 (
            .O(N__50104),
            .I(\c0.data_in_frame_8_3 ));
    InMux I__7981 (
            .O(N__50097),
            .I(N__50091));
    InMux I__7980 (
            .O(N__50096),
            .I(N__50091));
    LocalMux I__7979 (
            .O(N__50091),
            .I(\c0.n33874 ));
    InMux I__7978 (
            .O(N__50088),
            .I(N__50085));
    LocalMux I__7977 (
            .O(N__50085),
            .I(\c0.n19064 ));
    InMux I__7976 (
            .O(N__50082),
            .I(N__50076));
    InMux I__7975 (
            .O(N__50081),
            .I(N__50073));
    InMux I__7974 (
            .O(N__50080),
            .I(N__50068));
    InMux I__7973 (
            .O(N__50079),
            .I(N__50068));
    LocalMux I__7972 (
            .O(N__50076),
            .I(N__50063));
    LocalMux I__7971 (
            .O(N__50073),
            .I(N__50063));
    LocalMux I__7970 (
            .O(N__50068),
            .I(N__50059));
    Span4Mux_h I__7969 (
            .O(N__50063),
            .I(N__50056));
    CascadeMux I__7968 (
            .O(N__50062),
            .I(N__50053));
    Span4Mux_h I__7967 (
            .O(N__50059),
            .I(N__50048));
    Span4Mux_h I__7966 (
            .O(N__50056),
            .I(N__50048));
    InMux I__7965 (
            .O(N__50053),
            .I(N__50045));
    Span4Mux_v I__7964 (
            .O(N__50048),
            .I(N__50042));
    LocalMux I__7963 (
            .O(N__50045),
            .I(\c0.data_in_frame_13_2 ));
    Odrv4 I__7962 (
            .O(N__50042),
            .I(\c0.data_in_frame_13_2 ));
    InMux I__7961 (
            .O(N__50037),
            .I(N__50033));
    InMux I__7960 (
            .O(N__50036),
            .I(N__50029));
    LocalMux I__7959 (
            .O(N__50033),
            .I(N__50026));
    InMux I__7958 (
            .O(N__50032),
            .I(N__50023));
    LocalMux I__7957 (
            .O(N__50029),
            .I(N__50020));
    Span4Mux_v I__7956 (
            .O(N__50026),
            .I(N__50015));
    LocalMux I__7955 (
            .O(N__50023),
            .I(N__50015));
    Span4Mux_h I__7954 (
            .O(N__50020),
            .I(N__50012));
    Span4Mux_h I__7953 (
            .O(N__50015),
            .I(N__50006));
    Span4Mux_h I__7952 (
            .O(N__50012),
            .I(N__50006));
    InMux I__7951 (
            .O(N__50011),
            .I(N__50003));
    Span4Mux_v I__7950 (
            .O(N__50006),
            .I(N__50000));
    LocalMux I__7949 (
            .O(N__50003),
            .I(\c0.data_in_frame_13_3 ));
    Odrv4 I__7948 (
            .O(N__50000),
            .I(\c0.data_in_frame_13_3 ));
    CascadeMux I__7947 (
            .O(N__49995),
            .I(\c0.n18373_cascade_ ));
    InMux I__7946 (
            .O(N__49992),
            .I(N__49989));
    LocalMux I__7945 (
            .O(N__49989),
            .I(\c0.n5965 ));
    InMux I__7944 (
            .O(N__49986),
            .I(N__49983));
    LocalMux I__7943 (
            .O(N__49983),
            .I(\c0.n4_adj_4734 ));
    CascadeMux I__7942 (
            .O(N__49980),
            .I(\c0.n5965_cascade_ ));
    CascadeMux I__7941 (
            .O(N__49977),
            .I(N__49973));
    InMux I__7940 (
            .O(N__49976),
            .I(N__49970));
    InMux I__7939 (
            .O(N__49973),
            .I(N__49967));
    LocalMux I__7938 (
            .O(N__49970),
            .I(N__49964));
    LocalMux I__7937 (
            .O(N__49967),
            .I(\c0.data_in_frame_17_6 ));
    Odrv4 I__7936 (
            .O(N__49964),
            .I(\c0.data_in_frame_17_6 ));
    InMux I__7935 (
            .O(N__49959),
            .I(N__49955));
    InMux I__7934 (
            .O(N__49958),
            .I(N__49952));
    LocalMux I__7933 (
            .O(N__49955),
            .I(N__49949));
    LocalMux I__7932 (
            .O(N__49952),
            .I(\c0.n33708 ));
    Odrv4 I__7931 (
            .O(N__49949),
            .I(\c0.n33708 ));
    InMux I__7930 (
            .O(N__49944),
            .I(N__49941));
    LocalMux I__7929 (
            .O(N__49941),
            .I(\c0.n33877 ));
    CascadeMux I__7928 (
            .O(N__49938),
            .I(N__49933));
    InMux I__7927 (
            .O(N__49937),
            .I(N__49930));
    InMux I__7926 (
            .O(N__49936),
            .I(N__49927));
    InMux I__7925 (
            .O(N__49933),
            .I(N__49924));
    LocalMux I__7924 (
            .O(N__49930),
            .I(N__49921));
    LocalMux I__7923 (
            .O(N__49927),
            .I(N__49916));
    LocalMux I__7922 (
            .O(N__49924),
            .I(N__49916));
    Odrv4 I__7921 (
            .O(N__49921),
            .I(\c0.data_in_frame_4_2 ));
    Odrv4 I__7920 (
            .O(N__49916),
            .I(\c0.data_in_frame_4_2 ));
    CascadeMux I__7919 (
            .O(N__49911),
            .I(N__49907));
    InMux I__7918 (
            .O(N__49910),
            .I(N__49902));
    InMux I__7917 (
            .O(N__49907),
            .I(N__49902));
    LocalMux I__7916 (
            .O(N__49902),
            .I(\c0.data_in_frame_14_2 ));
    CascadeMux I__7915 (
            .O(N__49899),
            .I(N__49896));
    InMux I__7914 (
            .O(N__49896),
            .I(N__49887));
    InMux I__7913 (
            .O(N__49895),
            .I(N__49887));
    InMux I__7912 (
            .O(N__49894),
            .I(N__49887));
    LocalMux I__7911 (
            .O(N__49887),
            .I(\c0.data_in_frame_8_0 ));
    CascadeMux I__7910 (
            .O(N__49884),
            .I(N__49880));
    InMux I__7909 (
            .O(N__49883),
            .I(N__49876));
    InMux I__7908 (
            .O(N__49880),
            .I(N__49873));
    InMux I__7907 (
            .O(N__49879),
            .I(N__49870));
    LocalMux I__7906 (
            .O(N__49876),
            .I(N__49867));
    LocalMux I__7905 (
            .O(N__49873),
            .I(\c0.data_in_frame_10_4 ));
    LocalMux I__7904 (
            .O(N__49870),
            .I(\c0.data_in_frame_10_4 ));
    Odrv4 I__7903 (
            .O(N__49867),
            .I(\c0.data_in_frame_10_4 ));
    InMux I__7902 (
            .O(N__49860),
            .I(N__49855));
    CascadeMux I__7901 (
            .O(N__49859),
            .I(N__49852));
    CascadeMux I__7900 (
            .O(N__49858),
            .I(N__49849));
    LocalMux I__7899 (
            .O(N__49855),
            .I(N__49846));
    InMux I__7898 (
            .O(N__49852),
            .I(N__49843));
    InMux I__7897 (
            .O(N__49849),
            .I(N__49840));
    Span4Mux_v I__7896 (
            .O(N__49846),
            .I(N__49835));
    LocalMux I__7895 (
            .O(N__49843),
            .I(N__49835));
    LocalMux I__7894 (
            .O(N__49840),
            .I(N__49830));
    Span4Mux_h I__7893 (
            .O(N__49835),
            .I(N__49830));
    Odrv4 I__7892 (
            .O(N__49830),
            .I(\c0.data_in_frame_12_5 ));
    CascadeMux I__7891 (
            .O(N__49827),
            .I(\c0.n33874_cascade_ ));
    InMux I__7890 (
            .O(N__49824),
            .I(N__49820));
    CascadeMux I__7889 (
            .O(N__49823),
            .I(N__49817));
    LocalMux I__7888 (
            .O(N__49820),
            .I(N__49813));
    InMux I__7887 (
            .O(N__49817),
            .I(N__49808));
    InMux I__7886 (
            .O(N__49816),
            .I(N__49808));
    Span4Mux_v I__7885 (
            .O(N__49813),
            .I(N__49805));
    LocalMux I__7884 (
            .O(N__49808),
            .I(N__49802));
    Odrv4 I__7883 (
            .O(N__49805),
            .I(\c0.data_out_frame_0__7__N_2580 ));
    Odrv4 I__7882 (
            .O(N__49802),
            .I(\c0.data_out_frame_0__7__N_2580 ));
    CascadeMux I__7881 (
            .O(N__49797),
            .I(N__49794));
    InMux I__7880 (
            .O(N__49794),
            .I(N__49790));
    InMux I__7879 (
            .O(N__49793),
            .I(N__49787));
    LocalMux I__7878 (
            .O(N__49790),
            .I(\c0.n5_adj_4742 ));
    LocalMux I__7877 (
            .O(N__49787),
            .I(\c0.n5_adj_4742 ));
    InMux I__7876 (
            .O(N__49782),
            .I(N__49778));
    InMux I__7875 (
            .O(N__49781),
            .I(N__49775));
    LocalMux I__7874 (
            .O(N__49778),
            .I(N__49772));
    LocalMux I__7873 (
            .O(N__49775),
            .I(N__49769));
    Span4Mux_v I__7872 (
            .O(N__49772),
            .I(N__49766));
    Odrv12 I__7871 (
            .O(N__49769),
            .I(\c0.n33288 ));
    Odrv4 I__7870 (
            .O(N__49766),
            .I(\c0.n33288 ));
    InMux I__7869 (
            .O(N__49761),
            .I(N__49758));
    LocalMux I__7868 (
            .O(N__49758),
            .I(N__49755));
    Span4Mux_v I__7867 (
            .O(N__49755),
            .I(N__49751));
    InMux I__7866 (
            .O(N__49754),
            .I(N__49748));
    Odrv4 I__7865 (
            .O(N__49751),
            .I(\c0.n18705 ));
    LocalMux I__7864 (
            .O(N__49748),
            .I(\c0.n18705 ));
    InMux I__7863 (
            .O(N__49743),
            .I(N__49740));
    LocalMux I__7862 (
            .O(N__49740),
            .I(N__49736));
    CascadeMux I__7861 (
            .O(N__49739),
            .I(N__49733));
    Span4Mux_h I__7860 (
            .O(N__49736),
            .I(N__49729));
    InMux I__7859 (
            .O(N__49733),
            .I(N__49724));
    InMux I__7858 (
            .O(N__49732),
            .I(N__49724));
    Odrv4 I__7857 (
            .O(N__49729),
            .I(\c0.data_in_frame_8_2 ));
    LocalMux I__7856 (
            .O(N__49724),
            .I(\c0.data_in_frame_8_2 ));
    CascadeMux I__7855 (
            .O(N__49719),
            .I(\c0.n18705_cascade_ ));
    InMux I__7854 (
            .O(N__49716),
            .I(N__49713));
    LocalMux I__7853 (
            .O(N__49713),
            .I(N__49708));
    InMux I__7852 (
            .O(N__49712),
            .I(N__49705));
    InMux I__7851 (
            .O(N__49711),
            .I(N__49702));
    Odrv4 I__7850 (
            .O(N__49708),
            .I(\c0.n33291 ));
    LocalMux I__7849 (
            .O(N__49705),
            .I(\c0.n33291 ));
    LocalMux I__7848 (
            .O(N__49702),
            .I(\c0.n33291 ));
    InMux I__7847 (
            .O(N__49695),
            .I(N__49692));
    LocalMux I__7846 (
            .O(N__49692),
            .I(\c0.n10_adj_4743 ));
    InMux I__7845 (
            .O(N__49689),
            .I(N__49683));
    InMux I__7844 (
            .O(N__49688),
            .I(N__49679));
    InMux I__7843 (
            .O(N__49687),
            .I(N__49676));
    InMux I__7842 (
            .O(N__49686),
            .I(N__49673));
    LocalMux I__7841 (
            .O(N__49683),
            .I(N__49670));
    InMux I__7840 (
            .O(N__49682),
            .I(N__49667));
    LocalMux I__7839 (
            .O(N__49679),
            .I(\c0.n18709 ));
    LocalMux I__7838 (
            .O(N__49676),
            .I(\c0.n18709 ));
    LocalMux I__7837 (
            .O(N__49673),
            .I(\c0.n18709 ));
    Odrv4 I__7836 (
            .O(N__49670),
            .I(\c0.n18709 ));
    LocalMux I__7835 (
            .O(N__49667),
            .I(\c0.n18709 ));
    CascadeMux I__7834 (
            .O(N__49656),
            .I(N__49652));
    InMux I__7833 (
            .O(N__49655),
            .I(N__49649));
    InMux I__7832 (
            .O(N__49652),
            .I(N__49644));
    LocalMux I__7831 (
            .O(N__49649),
            .I(N__49641));
    InMux I__7830 (
            .O(N__49648),
            .I(N__49638));
    InMux I__7829 (
            .O(N__49647),
            .I(N__49635));
    LocalMux I__7828 (
            .O(N__49644),
            .I(N__49628));
    Span4Mux_h I__7827 (
            .O(N__49641),
            .I(N__49628));
    LocalMux I__7826 (
            .O(N__49638),
            .I(N__49628));
    LocalMux I__7825 (
            .O(N__49635),
            .I(N__49625));
    Odrv4 I__7824 (
            .O(N__49628),
            .I(\c0.data_in_frame_7_4 ));
    Odrv12 I__7823 (
            .O(N__49625),
            .I(\c0.data_in_frame_7_4 ));
    InMux I__7822 (
            .O(N__49620),
            .I(N__49617));
    LocalMux I__7821 (
            .O(N__49617),
            .I(N__49613));
    CascadeMux I__7820 (
            .O(N__49616),
            .I(N__49610));
    Span4Mux_h I__7819 (
            .O(N__49613),
            .I(N__49606));
    InMux I__7818 (
            .O(N__49610),
            .I(N__49601));
    InMux I__7817 (
            .O(N__49609),
            .I(N__49601));
    Odrv4 I__7816 (
            .O(N__49606),
            .I(\c0.data_in_frame_10_0 ));
    LocalMux I__7815 (
            .O(N__49601),
            .I(\c0.data_in_frame_10_0 ));
    CascadeMux I__7814 (
            .O(N__49596),
            .I(\c0.n8_adj_4555_cascade_ ));
    InMux I__7813 (
            .O(N__49593),
            .I(N__49590));
    LocalMux I__7812 (
            .O(N__49590),
            .I(N__49587));
    Odrv4 I__7811 (
            .O(N__49587),
            .I(\c0.n7_adj_4554 ));
    CascadeMux I__7810 (
            .O(N__49584),
            .I(\c0.n33441_cascade_ ));
    InMux I__7809 (
            .O(N__49581),
            .I(N__49577));
    InMux I__7808 (
            .O(N__49580),
            .I(N__49574));
    LocalMux I__7807 (
            .O(N__49577),
            .I(\c0.data_in_frame_7_7 ));
    LocalMux I__7806 (
            .O(N__49574),
            .I(\c0.data_in_frame_7_7 ));
    InMux I__7805 (
            .O(N__49569),
            .I(N__49565));
    InMux I__7804 (
            .O(N__49568),
            .I(N__49561));
    LocalMux I__7803 (
            .O(N__49565),
            .I(N__49558));
    InMux I__7802 (
            .O(N__49564),
            .I(N__49555));
    LocalMux I__7801 (
            .O(N__49561),
            .I(\c0.n18141 ));
    Odrv4 I__7800 (
            .O(N__49558),
            .I(\c0.n18141 ));
    LocalMux I__7799 (
            .O(N__49555),
            .I(\c0.n18141 ));
    CascadeMux I__7798 (
            .O(N__49548),
            .I(N__49545));
    InMux I__7797 (
            .O(N__49545),
            .I(N__49538));
    InMux I__7796 (
            .O(N__49544),
            .I(N__49538));
    InMux I__7795 (
            .O(N__49543),
            .I(N__49535));
    LocalMux I__7794 (
            .O(N__49538),
            .I(\c0.data_in_frame_7_6 ));
    LocalMux I__7793 (
            .O(N__49535),
            .I(\c0.data_in_frame_7_6 ));
    InMux I__7792 (
            .O(N__49530),
            .I(N__49527));
    LocalMux I__7791 (
            .O(N__49527),
            .I(\c0.n6_adj_4733 ));
    InMux I__7790 (
            .O(N__49524),
            .I(N__49519));
    InMux I__7789 (
            .O(N__49523),
            .I(N__49514));
    InMux I__7788 (
            .O(N__49522),
            .I(N__49514));
    LocalMux I__7787 (
            .O(N__49519),
            .I(N__49511));
    LocalMux I__7786 (
            .O(N__49514),
            .I(N__49508));
    Span4Mux_h I__7785 (
            .O(N__49511),
            .I(N__49505));
    Odrv4 I__7784 (
            .O(N__49508),
            .I(\c0.n32298 ));
    Odrv4 I__7783 (
            .O(N__49505),
            .I(\c0.n32298 ));
    InMux I__7782 (
            .O(N__49500),
            .I(N__49495));
    InMux I__7781 (
            .O(N__49499),
            .I(N__49490));
    InMux I__7780 (
            .O(N__49498),
            .I(N__49490));
    LocalMux I__7779 (
            .O(N__49495),
            .I(\c0.data_in_frame_9_7 ));
    LocalMux I__7778 (
            .O(N__49490),
            .I(\c0.data_in_frame_9_7 ));
    CascadeMux I__7777 (
            .O(N__49485),
            .I(N__49481));
    CascadeMux I__7776 (
            .O(N__49484),
            .I(N__49478));
    InMux I__7775 (
            .O(N__49481),
            .I(N__49475));
    InMux I__7774 (
            .O(N__49478),
            .I(N__49472));
    LocalMux I__7773 (
            .O(N__49475),
            .I(\c0.data_in_frame_10_1 ));
    LocalMux I__7772 (
            .O(N__49472),
            .I(\c0.data_in_frame_10_1 ));
    InMux I__7771 (
            .O(N__49467),
            .I(N__49464));
    LocalMux I__7770 (
            .O(N__49464),
            .I(N__49460));
    InMux I__7769 (
            .O(N__49463),
            .I(N__49457));
    Odrv4 I__7768 (
            .O(N__49460),
            .I(\c0.n33698 ));
    LocalMux I__7767 (
            .O(N__49457),
            .I(\c0.n33698 ));
    CascadeMux I__7766 (
            .O(N__49452),
            .I(N__49449));
    InMux I__7765 (
            .O(N__49449),
            .I(N__49446));
    LocalMux I__7764 (
            .O(N__49446),
            .I(N__49443));
    Odrv4 I__7763 (
            .O(N__49443),
            .I(\c0.n10_adj_4736 ));
    InMux I__7762 (
            .O(N__49440),
            .I(N__49435));
    CascadeMux I__7761 (
            .O(N__49439),
            .I(N__49430));
    CascadeMux I__7760 (
            .O(N__49438),
            .I(N__49425));
    LocalMux I__7759 (
            .O(N__49435),
            .I(N__49421));
    InMux I__7758 (
            .O(N__49434),
            .I(N__49418));
    InMux I__7757 (
            .O(N__49433),
            .I(N__49415));
    InMux I__7756 (
            .O(N__49430),
            .I(N__49406));
    InMux I__7755 (
            .O(N__49429),
            .I(N__49406));
    InMux I__7754 (
            .O(N__49428),
            .I(N__49406));
    InMux I__7753 (
            .O(N__49425),
            .I(N__49406));
    InMux I__7752 (
            .O(N__49424),
            .I(N__49403));
    Span4Mux_h I__7751 (
            .O(N__49421),
            .I(N__49400));
    LocalMux I__7750 (
            .O(N__49418),
            .I(N__49395));
    LocalMux I__7749 (
            .O(N__49415),
            .I(N__49395));
    LocalMux I__7748 (
            .O(N__49406),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__7747 (
            .O(N__49403),
            .I(\c0.data_in_frame_0_6 ));
    Odrv4 I__7746 (
            .O(N__49400),
            .I(\c0.data_in_frame_0_6 ));
    Odrv4 I__7745 (
            .O(N__49395),
            .I(\c0.data_in_frame_0_6 ));
    InMux I__7744 (
            .O(N__49386),
            .I(N__49383));
    LocalMux I__7743 (
            .O(N__49383),
            .I(\c0.n18354 ));
    InMux I__7742 (
            .O(N__49380),
            .I(N__49376));
    InMux I__7741 (
            .O(N__49379),
            .I(N__49373));
    LocalMux I__7740 (
            .O(N__49376),
            .I(N__49370));
    LocalMux I__7739 (
            .O(N__49373),
            .I(\c0.n33326 ));
    Odrv4 I__7738 (
            .O(N__49370),
            .I(\c0.n33326 ));
    InMux I__7737 (
            .O(N__49365),
            .I(N__49361));
    InMux I__7736 (
            .O(N__49364),
            .I(N__49358));
    LocalMux I__7735 (
            .O(N__49361),
            .I(N__49353));
    LocalMux I__7734 (
            .O(N__49358),
            .I(N__49353));
    Odrv12 I__7733 (
            .O(N__49353),
            .I(\c0.n33804 ));
    CascadeMux I__7732 (
            .O(N__49350),
            .I(\c0.n18354_cascade_ ));
    InMux I__7731 (
            .O(N__49347),
            .I(N__49344));
    LocalMux I__7730 (
            .O(N__49344),
            .I(N__49341));
    Span4Mux_h I__7729 (
            .O(N__49341),
            .I(N__49338));
    Odrv4 I__7728 (
            .O(N__49338),
            .I(\c0.n31_adj_4766 ));
    InMux I__7727 (
            .O(N__49335),
            .I(N__49332));
    LocalMux I__7726 (
            .O(N__49332),
            .I(N__49329));
    Span4Mux_h I__7725 (
            .O(N__49329),
            .I(N__49326));
    Odrv4 I__7724 (
            .O(N__49326),
            .I(\c0.n30_adj_4765 ));
    CascadeMux I__7723 (
            .O(N__49323),
            .I(\c0.n29_adj_4767_cascade_ ));
    InMux I__7722 (
            .O(N__49320),
            .I(N__49317));
    LocalMux I__7721 (
            .O(N__49317),
            .I(\c0.n33830 ));
    InMux I__7720 (
            .O(N__49314),
            .I(N__49311));
    LocalMux I__7719 (
            .O(N__49311),
            .I(N__49306));
    InMux I__7718 (
            .O(N__49310),
            .I(N__49303));
    InMux I__7717 (
            .O(N__49309),
            .I(N__49300));
    Span4Mux_h I__7716 (
            .O(N__49306),
            .I(N__49297));
    LocalMux I__7715 (
            .O(N__49303),
            .I(N__49294));
    LocalMux I__7714 (
            .O(N__49300),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__7713 (
            .O(N__49297),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__7712 (
            .O(N__49294),
            .I(\c0.data_in_frame_3_5 ));
    CascadeMux I__7711 (
            .O(N__49287),
            .I(\c0.n33830_cascade_ ));
    InMux I__7710 (
            .O(N__49284),
            .I(N__49281));
    LocalMux I__7709 (
            .O(N__49281),
            .I(\c0.n6_adj_4535 ));
    InMux I__7708 (
            .O(N__49278),
            .I(N__49265));
    InMux I__7707 (
            .O(N__49277),
            .I(N__49255));
    InMux I__7706 (
            .O(N__49276),
            .I(N__49255));
    InMux I__7705 (
            .O(N__49275),
            .I(N__49255));
    InMux I__7704 (
            .O(N__49274),
            .I(N__49250));
    InMux I__7703 (
            .O(N__49273),
            .I(N__49250));
    InMux I__7702 (
            .O(N__49272),
            .I(N__49247));
    InMux I__7701 (
            .O(N__49271),
            .I(N__49238));
    InMux I__7700 (
            .O(N__49270),
            .I(N__49238));
    InMux I__7699 (
            .O(N__49269),
            .I(N__49238));
    InMux I__7698 (
            .O(N__49268),
            .I(N__49238));
    LocalMux I__7697 (
            .O(N__49265),
            .I(N__49233));
    InMux I__7696 (
            .O(N__49264),
            .I(N__49228));
    InMux I__7695 (
            .O(N__49263),
            .I(N__49228));
    InMux I__7694 (
            .O(N__49262),
            .I(N__49225));
    LocalMux I__7693 (
            .O(N__49255),
            .I(N__49216));
    LocalMux I__7692 (
            .O(N__49250),
            .I(N__49216));
    LocalMux I__7691 (
            .O(N__49247),
            .I(N__49216));
    LocalMux I__7690 (
            .O(N__49238),
            .I(N__49216));
    InMux I__7689 (
            .O(N__49237),
            .I(N__49211));
    InMux I__7688 (
            .O(N__49236),
            .I(N__49211));
    Span4Mux_v I__7687 (
            .O(N__49233),
            .I(N__49206));
    LocalMux I__7686 (
            .O(N__49228),
            .I(N__49206));
    LocalMux I__7685 (
            .O(N__49225),
            .I(N__49203));
    Span4Mux_v I__7684 (
            .O(N__49216),
            .I(N__49200));
    LocalMux I__7683 (
            .O(N__49211),
            .I(N__49195));
    Span4Mux_h I__7682 (
            .O(N__49206),
            .I(N__49195));
    Span4Mux_v I__7681 (
            .O(N__49203),
            .I(N__49190));
    Span4Mux_h I__7680 (
            .O(N__49200),
            .I(N__49190));
    Odrv4 I__7679 (
            .O(N__49195),
            .I(\c0.n29668 ));
    Odrv4 I__7678 (
            .O(N__49190),
            .I(\c0.n29668 ));
    InMux I__7677 (
            .O(N__49185),
            .I(N__49181));
    CascadeMux I__7676 (
            .O(N__49184),
            .I(N__49177));
    LocalMux I__7675 (
            .O(N__49181),
            .I(N__49174));
    InMux I__7674 (
            .O(N__49180),
            .I(N__49168));
    InMux I__7673 (
            .O(N__49177),
            .I(N__49168));
    Span4Mux_v I__7672 (
            .O(N__49174),
            .I(N__49164));
    CascadeMux I__7671 (
            .O(N__49173),
            .I(N__49161));
    LocalMux I__7670 (
            .O(N__49168),
            .I(N__49157));
    CascadeMux I__7669 (
            .O(N__49167),
            .I(N__49153));
    Span4Mux_h I__7668 (
            .O(N__49164),
            .I(N__49150));
    InMux I__7667 (
            .O(N__49161),
            .I(N__49147));
    InMux I__7666 (
            .O(N__49160),
            .I(N__49144));
    Span4Mux_h I__7665 (
            .O(N__49157),
            .I(N__49141));
    InMux I__7664 (
            .O(N__49156),
            .I(N__49136));
    InMux I__7663 (
            .O(N__49153),
            .I(N__49136));
    Odrv4 I__7662 (
            .O(N__49150),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7661 (
            .O(N__49147),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7660 (
            .O(N__49144),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__7659 (
            .O(N__49141),
            .I(\c0.FRAME_MATCHER_state_0 ));
    LocalMux I__7658 (
            .O(N__49136),
            .I(\c0.FRAME_MATCHER_state_0 ));
    CascadeMux I__7657 (
            .O(N__49125),
            .I(\c0.n72_cascade_ ));
    InMux I__7656 (
            .O(N__49122),
            .I(N__49117));
    CascadeMux I__7655 (
            .O(N__49121),
            .I(N__49112));
    CascadeMux I__7654 (
            .O(N__49120),
            .I(N__49108));
    LocalMux I__7653 (
            .O(N__49117),
            .I(N__49105));
    InMux I__7652 (
            .O(N__49116),
            .I(N__49096));
    InMux I__7651 (
            .O(N__49115),
            .I(N__49096));
    InMux I__7650 (
            .O(N__49112),
            .I(N__49096));
    InMux I__7649 (
            .O(N__49111),
            .I(N__49096));
    InMux I__7648 (
            .O(N__49108),
            .I(N__49088));
    Span4Mux_v I__7647 (
            .O(N__49105),
            .I(N__49085));
    LocalMux I__7646 (
            .O(N__49096),
            .I(N__49082));
    InMux I__7645 (
            .O(N__49095),
            .I(N__49079));
    InMux I__7644 (
            .O(N__49094),
            .I(N__49074));
    InMux I__7643 (
            .O(N__49093),
            .I(N__49074));
    InMux I__7642 (
            .O(N__49092),
            .I(N__49067));
    InMux I__7641 (
            .O(N__49091),
            .I(N__49064));
    LocalMux I__7640 (
            .O(N__49088),
            .I(N__49061));
    Span4Mux_v I__7639 (
            .O(N__49085),
            .I(N__49056));
    Span4Mux_v I__7638 (
            .O(N__49082),
            .I(N__49056));
    LocalMux I__7637 (
            .O(N__49079),
            .I(N__49051));
    LocalMux I__7636 (
            .O(N__49074),
            .I(N__49051));
    InMux I__7635 (
            .O(N__49073),
            .I(N__49047));
    InMux I__7634 (
            .O(N__49072),
            .I(N__49040));
    InMux I__7633 (
            .O(N__49071),
            .I(N__49040));
    InMux I__7632 (
            .O(N__49070),
            .I(N__49040));
    LocalMux I__7631 (
            .O(N__49067),
            .I(N__49035));
    LocalMux I__7630 (
            .O(N__49064),
            .I(N__49035));
    Span4Mux_v I__7629 (
            .O(N__49061),
            .I(N__49028));
    Span4Mux_h I__7628 (
            .O(N__49056),
            .I(N__49028));
    Span4Mux_h I__7627 (
            .O(N__49051),
            .I(N__49028));
    InMux I__7626 (
            .O(N__49050),
            .I(N__49025));
    LocalMux I__7625 (
            .O(N__49047),
            .I(N__49020));
    LocalMux I__7624 (
            .O(N__49040),
            .I(N__49020));
    Span4Mux_h I__7623 (
            .O(N__49035),
            .I(N__49015));
    Span4Mux_h I__7622 (
            .O(N__49028),
            .I(N__49015));
    LocalMux I__7621 (
            .O(N__49025),
            .I(\c0.n11851 ));
    Odrv12 I__7620 (
            .O(N__49020),
            .I(\c0.n11851 ));
    Odrv4 I__7619 (
            .O(N__49015),
            .I(\c0.n11851 ));
    InMux I__7618 (
            .O(N__49008),
            .I(N__49004));
    InMux I__7617 (
            .O(N__49007),
            .I(N__49000));
    LocalMux I__7616 (
            .O(N__49004),
            .I(N__48997));
    InMux I__7615 (
            .O(N__49003),
            .I(N__48994));
    LocalMux I__7614 (
            .O(N__49000),
            .I(N__48991));
    Span4Mux_h I__7613 (
            .O(N__48997),
            .I(N__48988));
    LocalMux I__7612 (
            .O(N__48994),
            .I(N__48985));
    Odrv12 I__7611 (
            .O(N__48991),
            .I(\c0.data_out_frame_0__7__N_2570 ));
    Odrv4 I__7610 (
            .O(N__48988),
            .I(\c0.data_out_frame_0__7__N_2570 ));
    Odrv4 I__7609 (
            .O(N__48985),
            .I(\c0.data_out_frame_0__7__N_2570 ));
    CascadeMux I__7608 (
            .O(N__48978),
            .I(\c0.n18675_cascade_ ));
    InMux I__7607 (
            .O(N__48975),
            .I(N__48966));
    InMux I__7606 (
            .O(N__48974),
            .I(N__48966));
    InMux I__7605 (
            .O(N__48973),
            .I(N__48966));
    LocalMux I__7604 (
            .O(N__48966),
            .I(N__48962));
    InMux I__7603 (
            .O(N__48965),
            .I(N__48959));
    Span4Mux_v I__7602 (
            .O(N__48962),
            .I(N__48953));
    LocalMux I__7601 (
            .O(N__48959),
            .I(N__48953));
    CascadeMux I__7600 (
            .O(N__48958),
            .I(N__48950));
    Span4Mux_v I__7599 (
            .O(N__48953),
            .I(N__48947));
    InMux I__7598 (
            .O(N__48950),
            .I(N__48944));
    Span4Mux_h I__7597 (
            .O(N__48947),
            .I(N__48941));
    LocalMux I__7596 (
            .O(N__48944),
            .I(\c0.n5_adj_4545 ));
    Odrv4 I__7595 (
            .O(N__48941),
            .I(\c0.n5_adj_4545 ));
    InMux I__7594 (
            .O(N__48936),
            .I(N__48933));
    LocalMux I__7593 (
            .O(N__48933),
            .I(\c0.n18667 ));
    CascadeMux I__7592 (
            .O(N__48930),
            .I(\c0.n18667_cascade_ ));
    CascadeMux I__7591 (
            .O(N__48927),
            .I(N__48924));
    InMux I__7590 (
            .O(N__48924),
            .I(N__48921));
    LocalMux I__7589 (
            .O(N__48921),
            .I(N__48918));
    Span4Mux_v I__7588 (
            .O(N__48918),
            .I(N__48914));
    InMux I__7587 (
            .O(N__48917),
            .I(N__48911));
    Odrv4 I__7586 (
            .O(N__48914),
            .I(\c0.n33347 ));
    LocalMux I__7585 (
            .O(N__48911),
            .I(\c0.n33347 ));
    InMux I__7584 (
            .O(N__48906),
            .I(N__48901));
    InMux I__7583 (
            .O(N__48905),
            .I(N__48898));
    InMux I__7582 (
            .O(N__48904),
            .I(N__48894));
    LocalMux I__7581 (
            .O(N__48901),
            .I(N__48891));
    LocalMux I__7580 (
            .O(N__48898),
            .I(N__48888));
    InMux I__7579 (
            .O(N__48897),
            .I(N__48885));
    LocalMux I__7578 (
            .O(N__48894),
            .I(N__48882));
    Span4Mux_v I__7577 (
            .O(N__48891),
            .I(N__48879));
    Span4Mux_v I__7576 (
            .O(N__48888),
            .I(N__48874));
    LocalMux I__7575 (
            .O(N__48885),
            .I(N__48874));
    Span4Mux_v I__7574 (
            .O(N__48882),
            .I(N__48869));
    Span4Mux_v I__7573 (
            .O(N__48879),
            .I(N__48869));
    Span4Mux_h I__7572 (
            .O(N__48874),
            .I(N__48866));
    Odrv4 I__7571 (
            .O(N__48869),
            .I(\c0.n18319 ));
    Odrv4 I__7570 (
            .O(N__48866),
            .I(\c0.n18319 ));
    CascadeMux I__7569 (
            .O(N__48861),
            .I(N__48858));
    InMux I__7568 (
            .O(N__48858),
            .I(N__48855));
    LocalMux I__7567 (
            .O(N__48855),
            .I(N__48850));
    CascadeMux I__7566 (
            .O(N__48854),
            .I(N__48846));
    CascadeMux I__7565 (
            .O(N__48853),
            .I(N__48842));
    Span4Mux_v I__7564 (
            .O(N__48850),
            .I(N__48839));
    CascadeMux I__7563 (
            .O(N__48849),
            .I(N__48835));
    InMux I__7562 (
            .O(N__48846),
            .I(N__48829));
    InMux I__7561 (
            .O(N__48845),
            .I(N__48829));
    InMux I__7560 (
            .O(N__48842),
            .I(N__48826));
    Span4Mux_h I__7559 (
            .O(N__48839),
            .I(N__48823));
    InMux I__7558 (
            .O(N__48838),
            .I(N__48820));
    InMux I__7557 (
            .O(N__48835),
            .I(N__48815));
    InMux I__7556 (
            .O(N__48834),
            .I(N__48815));
    LocalMux I__7555 (
            .O(N__48829),
            .I(N__48810));
    LocalMux I__7554 (
            .O(N__48826),
            .I(N__48810));
    Odrv4 I__7553 (
            .O(N__48823),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__7552 (
            .O(N__48820),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__7551 (
            .O(N__48815),
            .I(\c0.data_in_frame_0_0 ));
    Odrv12 I__7550 (
            .O(N__48810),
            .I(\c0.data_in_frame_0_0 ));
    CascadeMux I__7549 (
            .O(N__48801),
            .I(N__48797));
    CascadeMux I__7548 (
            .O(N__48800),
            .I(N__48793));
    InMux I__7547 (
            .O(N__48797),
            .I(N__48788));
    InMux I__7546 (
            .O(N__48796),
            .I(N__48788));
    InMux I__7545 (
            .O(N__48793),
            .I(N__48784));
    LocalMux I__7544 (
            .O(N__48788),
            .I(N__48781));
    InMux I__7543 (
            .O(N__48787),
            .I(N__48778));
    LocalMux I__7542 (
            .O(N__48784),
            .I(\c0.data_in_frame_2_2 ));
    Odrv12 I__7541 (
            .O(N__48781),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__7540 (
            .O(N__48778),
            .I(\c0.data_in_frame_2_2 ));
    InMux I__7539 (
            .O(N__48771),
            .I(N__48768));
    LocalMux I__7538 (
            .O(N__48768),
            .I(\c0.n35806 ));
    CascadeMux I__7537 (
            .O(N__48765),
            .I(\c0.n4_adj_4537_cascade_ ));
    CascadeMux I__7536 (
            .O(N__48762),
            .I(\c0.n18020_cascade_ ));
    CascadeMux I__7535 (
            .O(N__48759),
            .I(\c0.n35757_cascade_ ));
    InMux I__7534 (
            .O(N__48756),
            .I(N__48752));
    CascadeMux I__7533 (
            .O(N__48755),
            .I(N__48749));
    LocalMux I__7532 (
            .O(N__48752),
            .I(N__48746));
    InMux I__7531 (
            .O(N__48749),
            .I(N__48743));
    Span4Mux_h I__7530 (
            .O(N__48746),
            .I(N__48738));
    LocalMux I__7529 (
            .O(N__48743),
            .I(N__48738));
    Span4Mux_h I__7528 (
            .O(N__48738),
            .I(N__48735));
    Odrv4 I__7527 (
            .O(N__48735),
            .I(\c0.n79 ));
    CascadeMux I__7526 (
            .O(N__48732),
            .I(\c0.n47_adj_4611_cascade_ ));
    InMux I__7525 (
            .O(N__48729),
            .I(N__48726));
    LocalMux I__7524 (
            .O(N__48726),
            .I(N__48723));
    Odrv4 I__7523 (
            .O(N__48723),
            .I(\c0.n58 ));
    InMux I__7522 (
            .O(N__48720),
            .I(N__48717));
    LocalMux I__7521 (
            .O(N__48717),
            .I(\c0.n4_adj_4612 ));
    InMux I__7520 (
            .O(N__48714),
            .I(N__48708));
    InMux I__7519 (
            .O(N__48713),
            .I(N__48708));
    LocalMux I__7518 (
            .O(N__48708),
            .I(N__48704));
    InMux I__7517 (
            .O(N__48707),
            .I(N__48700));
    Span4Mux_v I__7516 (
            .O(N__48704),
            .I(N__48697));
    InMux I__7515 (
            .O(N__48703),
            .I(N__48694));
    LocalMux I__7514 (
            .O(N__48700),
            .I(N__48691));
    Span4Mux_h I__7513 (
            .O(N__48697),
            .I(N__48688));
    LocalMux I__7512 (
            .O(N__48694),
            .I(data_in_3_1));
    Odrv12 I__7511 (
            .O(N__48691),
            .I(data_in_3_1));
    Odrv4 I__7510 (
            .O(N__48688),
            .I(data_in_3_1));
    InMux I__7509 (
            .O(N__48681),
            .I(N__48677));
    InMux I__7508 (
            .O(N__48680),
            .I(N__48674));
    LocalMux I__7507 (
            .O(N__48677),
            .I(\c0.n19909 ));
    LocalMux I__7506 (
            .O(N__48674),
            .I(\c0.n19909 ));
    InMux I__7505 (
            .O(N__48669),
            .I(N__48666));
    LocalMux I__7504 (
            .O(N__48666),
            .I(\c0.n30862 ));
    InMux I__7503 (
            .O(N__48663),
            .I(N__48657));
    InMux I__7502 (
            .O(N__48662),
            .I(N__48652));
    InMux I__7501 (
            .O(N__48661),
            .I(N__48652));
    InMux I__7500 (
            .O(N__48660),
            .I(N__48649));
    LocalMux I__7499 (
            .O(N__48657),
            .I(N__48646));
    LocalMux I__7498 (
            .O(N__48652),
            .I(N__48643));
    LocalMux I__7497 (
            .O(N__48649),
            .I(\c0.n4_adj_4537 ));
    Odrv4 I__7496 (
            .O(N__48646),
            .I(\c0.n4_adj_4537 ));
    Odrv4 I__7495 (
            .O(N__48643),
            .I(\c0.n4_adj_4537 ));
    CascadeMux I__7494 (
            .O(N__48636),
            .I(\c0.n30862_cascade_ ));
    InMux I__7493 (
            .O(N__48633),
            .I(N__48630));
    LocalMux I__7492 (
            .O(N__48630),
            .I(\c0.n72 ));
    CascadeMux I__7491 (
            .O(N__48627),
            .I(\c0.n14779_cascade_ ));
    InMux I__7490 (
            .O(N__48624),
            .I(N__48621));
    LocalMux I__7489 (
            .O(N__48621),
            .I(N__48618));
    Span4Mux_v I__7488 (
            .O(N__48618),
            .I(N__48615));
    Odrv4 I__7487 (
            .O(N__48615),
            .I(\c0.n6_adj_4617 ));
    CascadeMux I__7486 (
            .O(N__48612),
            .I(N__48609));
    InMux I__7485 (
            .O(N__48609),
            .I(N__48603));
    InMux I__7484 (
            .O(N__48608),
            .I(N__48603));
    LocalMux I__7483 (
            .O(N__48603),
            .I(\c0.n18115 ));
    InMux I__7482 (
            .O(N__48600),
            .I(N__48596));
    InMux I__7481 (
            .O(N__48599),
            .I(N__48593));
    LocalMux I__7480 (
            .O(N__48596),
            .I(N__48586));
    LocalMux I__7479 (
            .O(N__48593),
            .I(N__48586));
    InMux I__7478 (
            .O(N__48592),
            .I(N__48581));
    InMux I__7477 (
            .O(N__48591),
            .I(N__48581));
    Span4Mux_h I__7476 (
            .O(N__48586),
            .I(N__48578));
    LocalMux I__7475 (
            .O(N__48581),
            .I(N__48575));
    Span4Mux_h I__7474 (
            .O(N__48578),
            .I(N__48572));
    Span4Mux_v I__7473 (
            .O(N__48575),
            .I(N__48569));
    Span4Mux_h I__7472 (
            .O(N__48572),
            .I(N__48566));
    Odrv4 I__7471 (
            .O(N__48569),
            .I(\c0.n33166 ));
    Odrv4 I__7470 (
            .O(N__48566),
            .I(\c0.n33166 ));
    CascadeMux I__7469 (
            .O(N__48561),
            .I(N__48558));
    InMux I__7468 (
            .O(N__48558),
            .I(N__48552));
    InMux I__7467 (
            .O(N__48557),
            .I(N__48552));
    LocalMux I__7466 (
            .O(N__48552),
            .I(N__48549));
    Span4Mux_h I__7465 (
            .O(N__48549),
            .I(N__48546));
    Span4Mux_h I__7464 (
            .O(N__48546),
            .I(N__48543));
    Odrv4 I__7463 (
            .O(N__48543),
            .I(\c0.n19820 ));
    InMux I__7462 (
            .O(N__48540),
            .I(N__48535));
    InMux I__7461 (
            .O(N__48539),
            .I(N__48532));
    InMux I__7460 (
            .O(N__48538),
            .I(N__48528));
    LocalMux I__7459 (
            .O(N__48535),
            .I(N__48525));
    LocalMux I__7458 (
            .O(N__48532),
            .I(N__48522));
    InMux I__7457 (
            .O(N__48531),
            .I(N__48519));
    LocalMux I__7456 (
            .O(N__48528),
            .I(N__48516));
    Span4Mux_v I__7455 (
            .O(N__48525),
            .I(N__48509));
    Span4Mux_h I__7454 (
            .O(N__48522),
            .I(N__48509));
    LocalMux I__7453 (
            .O(N__48519),
            .I(N__48509));
    Span4Mux_v I__7452 (
            .O(N__48516),
            .I(N__48502));
    Span4Mux_h I__7451 (
            .O(N__48509),
            .I(N__48502));
    InMux I__7450 (
            .O(N__48508),
            .I(N__48497));
    InMux I__7449 (
            .O(N__48507),
            .I(N__48497));
    Odrv4 I__7448 (
            .O(N__48502),
            .I(\c0.n14779 ));
    LocalMux I__7447 (
            .O(N__48497),
            .I(\c0.n14779 ));
    InMux I__7446 (
            .O(N__48492),
            .I(N__48487));
    CascadeMux I__7445 (
            .O(N__48491),
            .I(N__48484));
    InMux I__7444 (
            .O(N__48490),
            .I(N__48481));
    LocalMux I__7443 (
            .O(N__48487),
            .I(N__48477));
    InMux I__7442 (
            .O(N__48484),
            .I(N__48474));
    LocalMux I__7441 (
            .O(N__48481),
            .I(N__48470));
    InMux I__7440 (
            .O(N__48480),
            .I(N__48467));
    Span4Mux_v I__7439 (
            .O(N__48477),
            .I(N__48462));
    LocalMux I__7438 (
            .O(N__48474),
            .I(N__48462));
    InMux I__7437 (
            .O(N__48473),
            .I(N__48459));
    Span12Mux_v I__7436 (
            .O(N__48470),
            .I(N__48454));
    LocalMux I__7435 (
            .O(N__48467),
            .I(N__48454));
    Odrv4 I__7434 (
            .O(N__48462),
            .I(\c0.data_out_frame_0__7__N_2569 ));
    LocalMux I__7433 (
            .O(N__48459),
            .I(\c0.data_out_frame_0__7__N_2569 ));
    Odrv12 I__7432 (
            .O(N__48454),
            .I(\c0.data_out_frame_0__7__N_2569 ));
    InMux I__7431 (
            .O(N__48447),
            .I(N__48444));
    LocalMux I__7430 (
            .O(N__48444),
            .I(N__48440));
    InMux I__7429 (
            .O(N__48443),
            .I(N__48437));
    Span4Mux_v I__7428 (
            .O(N__48440),
            .I(N__48433));
    LocalMux I__7427 (
            .O(N__48437),
            .I(N__48430));
    CascadeMux I__7426 (
            .O(N__48436),
            .I(N__48427));
    Span4Mux_h I__7425 (
            .O(N__48433),
            .I(N__48424));
    Span4Mux_h I__7424 (
            .O(N__48430),
            .I(N__48421));
    InMux I__7423 (
            .O(N__48427),
            .I(N__48418));
    Sp12to4 I__7422 (
            .O(N__48424),
            .I(N__48415));
    Odrv4 I__7421 (
            .O(N__48421),
            .I(\c0.n688 ));
    LocalMux I__7420 (
            .O(N__48418),
            .I(\c0.n688 ));
    Odrv12 I__7419 (
            .O(N__48415),
            .I(\c0.n688 ));
    InMux I__7418 (
            .O(N__48408),
            .I(N__48405));
    LocalMux I__7417 (
            .O(N__48405),
            .I(\c0.n118 ));
    InMux I__7416 (
            .O(N__48402),
            .I(N__48395));
    InMux I__7415 (
            .O(N__48401),
            .I(N__48395));
    InMux I__7414 (
            .O(N__48400),
            .I(N__48392));
    LocalMux I__7413 (
            .O(N__48395),
            .I(N__48389));
    LocalMux I__7412 (
            .O(N__48392),
            .I(N__48386));
    Span4Mux_h I__7411 (
            .O(N__48389),
            .I(N__48383));
    Span4Mux_h I__7410 (
            .O(N__48386),
            .I(N__48380));
    Span4Mux_h I__7409 (
            .O(N__48383),
            .I(N__48377));
    Odrv4 I__7408 (
            .O(N__48380),
            .I(\c0.n30958 ));
    Odrv4 I__7407 (
            .O(N__48377),
            .I(\c0.n30958 ));
    InMux I__7406 (
            .O(N__48372),
            .I(N__48369));
    LocalMux I__7405 (
            .O(N__48369),
            .I(N__48366));
    Odrv12 I__7404 (
            .O(N__48366),
            .I(\c0.n18100 ));
    CascadeMux I__7403 (
            .O(N__48363),
            .I(\c0.n18100_cascade_ ));
    InMux I__7402 (
            .O(N__48360),
            .I(N__48355));
    InMux I__7401 (
            .O(N__48359),
            .I(N__48350));
    InMux I__7400 (
            .O(N__48358),
            .I(N__48350));
    LocalMux I__7399 (
            .O(N__48355),
            .I(\c0.n18045 ));
    LocalMux I__7398 (
            .O(N__48350),
            .I(\c0.n18045 ));
    InMux I__7397 (
            .O(N__48345),
            .I(N__48341));
    CascadeMux I__7396 (
            .O(N__48344),
            .I(N__48338));
    LocalMux I__7395 (
            .O(N__48341),
            .I(N__48335));
    InMux I__7394 (
            .O(N__48338),
            .I(N__48332));
    Span4Mux_h I__7393 (
            .O(N__48335),
            .I(N__48329));
    LocalMux I__7392 (
            .O(N__48332),
            .I(\c0.n31012 ));
    Odrv4 I__7391 (
            .O(N__48329),
            .I(\c0.n31012 ));
    InMux I__7390 (
            .O(N__48324),
            .I(N__48321));
    LocalMux I__7389 (
            .O(N__48321),
            .I(N__48318));
    Odrv4 I__7388 (
            .O(N__48318),
            .I(\c0.n111 ));
    CascadeMux I__7387 (
            .O(N__48315),
            .I(\c0.data_out_frame_0__7__N_2569_cascade_ ));
    InMux I__7386 (
            .O(N__48312),
            .I(N__48309));
    LocalMux I__7385 (
            .O(N__48309),
            .I(N__48305));
    InMux I__7384 (
            .O(N__48308),
            .I(N__48302));
    Span4Mux_h I__7383 (
            .O(N__48305),
            .I(N__48299));
    LocalMux I__7382 (
            .O(N__48302),
            .I(\c0.n33170 ));
    Odrv4 I__7381 (
            .O(N__48299),
            .I(\c0.n33170 ));
    CascadeMux I__7380 (
            .O(N__48294),
            .I(N__48290));
    InMux I__7379 (
            .O(N__48293),
            .I(N__48284));
    InMux I__7378 (
            .O(N__48290),
            .I(N__48284));
    InMux I__7377 (
            .O(N__48289),
            .I(N__48278));
    LocalMux I__7376 (
            .O(N__48284),
            .I(N__48275));
    InMux I__7375 (
            .O(N__48283),
            .I(N__48272));
    InMux I__7374 (
            .O(N__48282),
            .I(N__48267));
    InMux I__7373 (
            .O(N__48281),
            .I(N__48267));
    LocalMux I__7372 (
            .O(N__48278),
            .I(N__48264));
    Span4Mux_v I__7371 (
            .O(N__48275),
            .I(N__48261));
    LocalMux I__7370 (
            .O(N__48272),
            .I(N__48256));
    LocalMux I__7369 (
            .O(N__48267),
            .I(N__48256));
    Span12Mux_s11_h I__7368 (
            .O(N__48264),
            .I(N__48253));
    Span4Mux_h I__7367 (
            .O(N__48261),
            .I(N__48250));
    Span4Mux_v I__7366 (
            .O(N__48256),
            .I(N__48247));
    Odrv12 I__7365 (
            .O(N__48253),
            .I(r_SM_Main_2_N_3755_0));
    Odrv4 I__7364 (
            .O(N__48250),
            .I(r_SM_Main_2_N_3755_0));
    Odrv4 I__7363 (
            .O(N__48247),
            .I(r_SM_Main_2_N_3755_0));
    CascadeMux I__7362 (
            .O(N__48240),
            .I(N__48235));
    InMux I__7361 (
            .O(N__48239),
            .I(N__48228));
    InMux I__7360 (
            .O(N__48238),
            .I(N__48228));
    InMux I__7359 (
            .O(N__48235),
            .I(N__48228));
    LocalMux I__7358 (
            .O(N__48228),
            .I(N__48225));
    Span4Mux_v I__7357 (
            .O(N__48225),
            .I(N__48222));
    Span4Mux_h I__7356 (
            .O(N__48222),
            .I(N__48218));
    InMux I__7355 (
            .O(N__48221),
            .I(N__48215));
    Span4Mux_h I__7354 (
            .O(N__48218),
            .I(N__48212));
    LocalMux I__7353 (
            .O(N__48215),
            .I(\c0.tx_active ));
    Odrv4 I__7352 (
            .O(N__48212),
            .I(\c0.tx_active ));
    InMux I__7351 (
            .O(N__48207),
            .I(N__48204));
    LocalMux I__7350 (
            .O(N__48204),
            .I(\c0.n35938 ));
    InMux I__7349 (
            .O(N__48201),
            .I(N__48198));
    LocalMux I__7348 (
            .O(N__48198),
            .I(N__48195));
    Odrv12 I__7347 (
            .O(N__48195),
            .I(\c0.n6_adj_4638 ));
    InMux I__7346 (
            .O(N__48192),
            .I(N__48187));
    InMux I__7345 (
            .O(N__48191),
            .I(N__48184));
    InMux I__7344 (
            .O(N__48190),
            .I(N__48181));
    LocalMux I__7343 (
            .O(N__48187),
            .I(N__48178));
    LocalMux I__7342 (
            .O(N__48184),
            .I(N__48175));
    LocalMux I__7341 (
            .O(N__48181),
            .I(N__48172));
    Span4Mux_v I__7340 (
            .O(N__48178),
            .I(N__48169));
    Span4Mux_v I__7339 (
            .O(N__48175),
            .I(N__48164));
    Span4Mux_h I__7338 (
            .O(N__48172),
            .I(N__48164));
    Sp12to4 I__7337 (
            .O(N__48169),
            .I(N__48161));
    Span4Mux_h I__7336 (
            .O(N__48164),
            .I(N__48158));
    Odrv12 I__7335 (
            .O(N__48161),
            .I(\c0.n35339 ));
    Odrv4 I__7334 (
            .O(N__48158),
            .I(\c0.n35339 ));
    CascadeMux I__7333 (
            .O(N__48153),
            .I(\quad_counter0.n28331_cascade_ ));
    CascadeMux I__7332 (
            .O(N__48150),
            .I(\quad_counter0.n10_adj_4402_cascade_ ));
    InMux I__7331 (
            .O(N__48147),
            .I(N__48144));
    LocalMux I__7330 (
            .O(N__48144),
            .I(\quad_counter0.n16_adj_4403 ));
    InMux I__7329 (
            .O(N__48141),
            .I(N__48138));
    LocalMux I__7328 (
            .O(N__48138),
            .I(\quad_counter0.n14_adj_4404 ));
    CascadeMux I__7327 (
            .O(N__48135),
            .I(\quad_counter0.n18_adj_4405_cascade_ ));
    CascadeMux I__7326 (
            .O(N__48132),
            .I(N__48120));
    CascadeMux I__7325 (
            .O(N__48131),
            .I(N__48117));
    CascadeMux I__7324 (
            .O(N__48130),
            .I(N__48114));
    CascadeMux I__7323 (
            .O(N__48129),
            .I(N__48111));
    CascadeMux I__7322 (
            .O(N__48128),
            .I(N__48108));
    CascadeMux I__7321 (
            .O(N__48127),
            .I(N__48105));
    CascadeMux I__7320 (
            .O(N__48126),
            .I(N__48102));
    CascadeMux I__7319 (
            .O(N__48125),
            .I(N__48099));
    CascadeMux I__7318 (
            .O(N__48124),
            .I(N__48096));
    CascadeMux I__7317 (
            .O(N__48123),
            .I(N__48093));
    InMux I__7316 (
            .O(N__48120),
            .I(N__48084));
    InMux I__7315 (
            .O(N__48117),
            .I(N__48084));
    InMux I__7314 (
            .O(N__48114),
            .I(N__48084));
    InMux I__7313 (
            .O(N__48111),
            .I(N__48084));
    InMux I__7312 (
            .O(N__48108),
            .I(N__48075));
    InMux I__7311 (
            .O(N__48105),
            .I(N__48075));
    InMux I__7310 (
            .O(N__48102),
            .I(N__48075));
    InMux I__7309 (
            .O(N__48099),
            .I(N__48075));
    InMux I__7308 (
            .O(N__48096),
            .I(N__48070));
    InMux I__7307 (
            .O(N__48093),
            .I(N__48070));
    LocalMux I__7306 (
            .O(N__48084),
            .I(\quad_counter0.n2738 ));
    LocalMux I__7305 (
            .O(N__48075),
            .I(\quad_counter0.n2738 ));
    LocalMux I__7304 (
            .O(N__48070),
            .I(\quad_counter0.n2738 ));
    CascadeMux I__7303 (
            .O(N__48063),
            .I(\quad_counter0.n2738_cascade_ ));
    CascadeMux I__7302 (
            .O(N__48060),
            .I(N__48052));
    CascadeMux I__7301 (
            .O(N__48059),
            .I(N__48049));
    CascadeMux I__7300 (
            .O(N__48058),
            .I(N__48046));
    CascadeMux I__7299 (
            .O(N__48057),
            .I(N__48043));
    CascadeMux I__7298 (
            .O(N__48056),
            .I(N__48040));
    CascadeMux I__7297 (
            .O(N__48055),
            .I(N__48037));
    InMux I__7296 (
            .O(N__48052),
            .I(N__48032));
    InMux I__7295 (
            .O(N__48049),
            .I(N__48032));
    InMux I__7294 (
            .O(N__48046),
            .I(N__48023));
    InMux I__7293 (
            .O(N__48043),
            .I(N__48023));
    InMux I__7292 (
            .O(N__48040),
            .I(N__48023));
    InMux I__7291 (
            .O(N__48037),
            .I(N__48023));
    LocalMux I__7290 (
            .O(N__48032),
            .I(\quad_counter0.n36149 ));
    LocalMux I__7289 (
            .O(N__48023),
            .I(\quad_counter0.n36149 ));
    CascadeMux I__7288 (
            .O(N__48018),
            .I(\quad_counter0.n8_adj_4369_cascade_ ));
    InMux I__7287 (
            .O(N__48015),
            .I(N__48010));
    InMux I__7286 (
            .O(N__48014),
            .I(N__48007));
    InMux I__7285 (
            .O(N__48013),
            .I(N__48004));
    LocalMux I__7284 (
            .O(N__48010),
            .I(N__47999));
    LocalMux I__7283 (
            .O(N__48007),
            .I(N__47999));
    LocalMux I__7282 (
            .O(N__48004),
            .I(N__47996));
    Odrv12 I__7281 (
            .O(N__47999),
            .I(\quad_counter0.n3319 ));
    Odrv4 I__7280 (
            .O(N__47996),
            .I(\quad_counter0.n3319 ));
    InMux I__7279 (
            .O(N__47991),
            .I(N__47986));
    InMux I__7278 (
            .O(N__47990),
            .I(N__47983));
    InMux I__7277 (
            .O(N__47989),
            .I(N__47980));
    LocalMux I__7276 (
            .O(N__47986),
            .I(N__47975));
    LocalMux I__7275 (
            .O(N__47983),
            .I(N__47975));
    LocalMux I__7274 (
            .O(N__47980),
            .I(N__47972));
    Odrv12 I__7273 (
            .O(N__47975),
            .I(\quad_counter0.n3318 ));
    Odrv4 I__7272 (
            .O(N__47972),
            .I(\quad_counter0.n3318 ));
    InMux I__7271 (
            .O(N__47967),
            .I(N__47964));
    LocalMux I__7270 (
            .O(N__47964),
            .I(\quad_counter0.n7_adj_4363 ));
    InMux I__7269 (
            .O(N__47961),
            .I(N__47958));
    LocalMux I__7268 (
            .O(N__47958),
            .I(\quad_counter0.n7_adj_4370 ));
    CascadeMux I__7267 (
            .O(N__47955),
            .I(\quad_counter0.n18_adj_4368_cascade_ ));
    InMux I__7266 (
            .O(N__47952),
            .I(N__47949));
    LocalMux I__7265 (
            .O(N__47949),
            .I(\quad_counter0.n34805 ));
    InMux I__7264 (
            .O(N__47946),
            .I(N__47943));
    LocalMux I__7263 (
            .O(N__47943),
            .I(N__47940));
    Odrv4 I__7262 (
            .O(N__47940),
            .I(\quad_counter0.n7_adj_4395 ));
    CascadeMux I__7261 (
            .O(N__47937),
            .I(N__47933));
    InMux I__7260 (
            .O(N__47936),
            .I(N__47929));
    InMux I__7259 (
            .O(N__47933),
            .I(N__47926));
    InMux I__7258 (
            .O(N__47932),
            .I(N__47923));
    LocalMux I__7257 (
            .O(N__47929),
            .I(\quad_counter0.n1917 ));
    LocalMux I__7256 (
            .O(N__47926),
            .I(\quad_counter0.n1917 ));
    LocalMux I__7255 (
            .O(N__47923),
            .I(\quad_counter0.n1917 ));
    InMux I__7254 (
            .O(N__47916),
            .I(N__47913));
    LocalMux I__7253 (
            .O(N__47913),
            .I(\quad_counter0.n1984 ));
    InMux I__7252 (
            .O(N__47910),
            .I(\quad_counter0.n30217 ));
    CascadeMux I__7251 (
            .O(N__47907),
            .I(N__47903));
    CascadeMux I__7250 (
            .O(N__47906),
            .I(N__47899));
    InMux I__7249 (
            .O(N__47903),
            .I(N__47896));
    InMux I__7248 (
            .O(N__47902),
            .I(N__47891));
    InMux I__7247 (
            .O(N__47899),
            .I(N__47891));
    LocalMux I__7246 (
            .O(N__47896),
            .I(\quad_counter0.n1916 ));
    LocalMux I__7245 (
            .O(N__47891),
            .I(\quad_counter0.n1916 ));
    InMux I__7244 (
            .O(N__47886),
            .I(N__47883));
    LocalMux I__7243 (
            .O(N__47883),
            .I(\quad_counter0.n1983 ));
    InMux I__7242 (
            .O(N__47880),
            .I(\quad_counter0.n30218 ));
    InMux I__7241 (
            .O(N__47877),
            .I(\quad_counter0.n30219 ));
    CascadeMux I__7240 (
            .O(N__47874),
            .I(N__47870));
    CascadeMux I__7239 (
            .O(N__47873),
            .I(N__47867));
    InMux I__7238 (
            .O(N__47870),
            .I(N__47863));
    InMux I__7237 (
            .O(N__47867),
            .I(N__47860));
    InMux I__7236 (
            .O(N__47866),
            .I(N__47857));
    LocalMux I__7235 (
            .O(N__47863),
            .I(\quad_counter0.n1914 ));
    LocalMux I__7234 (
            .O(N__47860),
            .I(\quad_counter0.n1914 ));
    LocalMux I__7233 (
            .O(N__47857),
            .I(\quad_counter0.n1914 ));
    InMux I__7232 (
            .O(N__47850),
            .I(N__47847));
    LocalMux I__7231 (
            .O(N__47847),
            .I(\quad_counter0.n1981 ));
    InMux I__7230 (
            .O(N__47844),
            .I(\quad_counter0.n30220 ));
    InMux I__7229 (
            .O(N__47841),
            .I(N__47837));
    InMux I__7228 (
            .O(N__47840),
            .I(N__47834));
    LocalMux I__7227 (
            .O(N__47837),
            .I(\quad_counter0.n1913 ));
    LocalMux I__7226 (
            .O(N__47834),
            .I(\quad_counter0.n1913 ));
    InMux I__7225 (
            .O(N__47829),
            .I(\quad_counter0.n30221 ));
    InMux I__7224 (
            .O(N__47826),
            .I(N__47821));
    InMux I__7223 (
            .O(N__47825),
            .I(N__47818));
    InMux I__7222 (
            .O(N__47824),
            .I(N__47815));
    LocalMux I__7221 (
            .O(N__47821),
            .I(N__47808));
    LocalMux I__7220 (
            .O(N__47818),
            .I(N__47808));
    LocalMux I__7219 (
            .O(N__47815),
            .I(N__47808));
    Odrv4 I__7218 (
            .O(N__47808),
            .I(\quad_counter0.n3316 ));
    CascadeMux I__7217 (
            .O(N__47805),
            .I(N__47800));
    InMux I__7216 (
            .O(N__47804),
            .I(N__47797));
    InMux I__7215 (
            .O(N__47803),
            .I(N__47794));
    InMux I__7214 (
            .O(N__47800),
            .I(N__47791));
    LocalMux I__7213 (
            .O(N__47797),
            .I(N__47784));
    LocalMux I__7212 (
            .O(N__47794),
            .I(N__47784));
    LocalMux I__7211 (
            .O(N__47791),
            .I(N__47784));
    Odrv4 I__7210 (
            .O(N__47784),
            .I(\quad_counter0.n3315 ));
    InMux I__7209 (
            .O(N__47781),
            .I(N__47778));
    LocalMux I__7208 (
            .O(N__47778),
            .I(N__47775));
    Span4Mux_h I__7207 (
            .O(N__47775),
            .I(N__47772));
    Odrv4 I__7206 (
            .O(N__47772),
            .I(\quad_counter0.n35311 ));
    InMux I__7205 (
            .O(N__47769),
            .I(N__47764));
    InMux I__7204 (
            .O(N__47768),
            .I(N__47761));
    InMux I__7203 (
            .O(N__47767),
            .I(N__47758));
    LocalMux I__7202 (
            .O(N__47764),
            .I(N__47751));
    LocalMux I__7201 (
            .O(N__47761),
            .I(N__47751));
    LocalMux I__7200 (
            .O(N__47758),
            .I(N__47751));
    Odrv4 I__7199 (
            .O(N__47751),
            .I(\quad_counter0.n3317 ));
    InMux I__7198 (
            .O(N__47748),
            .I(N__47743));
    InMux I__7197 (
            .O(N__47747),
            .I(N__47740));
    InMux I__7196 (
            .O(N__47746),
            .I(N__47737));
    LocalMux I__7195 (
            .O(N__47743),
            .I(N__47730));
    LocalMux I__7194 (
            .O(N__47740),
            .I(N__47730));
    LocalMux I__7193 (
            .O(N__47737),
            .I(N__47730));
    Odrv4 I__7192 (
            .O(N__47730),
            .I(\quad_counter0.n3314 ));
    InMux I__7191 (
            .O(N__47727),
            .I(N__47724));
    LocalMux I__7190 (
            .O(N__47724),
            .I(\quad_counter0.n8_adj_4362 ));
    InMux I__7189 (
            .O(N__47721),
            .I(N__47718));
    LocalMux I__7188 (
            .O(N__47718),
            .I(\quad_counter0.n10_adj_4377 ));
    CascadeMux I__7187 (
            .O(N__47715),
            .I(\quad_counter0.n1946_cascade_ ));
    CascadeMux I__7186 (
            .O(N__47712),
            .I(\quad_counter0.n2019_cascade_ ));
    CascadeMux I__7185 (
            .O(N__47709),
            .I(N__47706));
    InMux I__7184 (
            .O(N__47706),
            .I(N__47703));
    LocalMux I__7183 (
            .O(N__47703),
            .I(\quad_counter0.n1987 ));
    InMux I__7182 (
            .O(N__47700),
            .I(bfn_13_7_0_));
    InMux I__7181 (
            .O(N__47697),
            .I(\quad_counter0.n30215 ));
    InMux I__7180 (
            .O(N__47694),
            .I(\quad_counter0.n30216 ));
    InMux I__7179 (
            .O(N__47691),
            .I(N__47688));
    LocalMux I__7178 (
            .O(N__47688),
            .I(\c0.n33308 ));
    InMux I__7177 (
            .O(N__47685),
            .I(N__47680));
    InMux I__7176 (
            .O(N__47684),
            .I(N__47677));
    InMux I__7175 (
            .O(N__47683),
            .I(N__47674));
    LocalMux I__7174 (
            .O(N__47680),
            .I(N__47669));
    LocalMux I__7173 (
            .O(N__47677),
            .I(N__47669));
    LocalMux I__7172 (
            .O(N__47674),
            .I(\c0.n33735 ));
    Odrv4 I__7171 (
            .O(N__47669),
            .I(\c0.n33735 ));
    CascadeMux I__7170 (
            .O(N__47664),
            .I(\c0.n33308_cascade_ ));
    InMux I__7169 (
            .O(N__47661),
            .I(N__47658));
    LocalMux I__7168 (
            .O(N__47658),
            .I(N__47655));
    Odrv4 I__7167 (
            .O(N__47655),
            .I(\c0.n36 ));
    InMux I__7166 (
            .O(N__47652),
            .I(N__47649));
    LocalMux I__7165 (
            .O(N__47649),
            .I(N__47646));
    Span4Mux_v I__7164 (
            .O(N__47646),
            .I(N__47641));
    InMux I__7163 (
            .O(N__47645),
            .I(N__47638));
    InMux I__7162 (
            .O(N__47644),
            .I(N__47635));
    Span4Mux_h I__7161 (
            .O(N__47641),
            .I(N__47630));
    LocalMux I__7160 (
            .O(N__47638),
            .I(N__47630));
    LocalMux I__7159 (
            .O(N__47635),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__7158 (
            .O(N__47630),
            .I(\c0.data_in_frame_19_7 ));
    CascadeMux I__7157 (
            .O(N__47625),
            .I(N__47622));
    InMux I__7156 (
            .O(N__47622),
            .I(N__47619));
    LocalMux I__7155 (
            .O(N__47619),
            .I(N__47616));
    Span4Mux_h I__7154 (
            .O(N__47616),
            .I(N__47613));
    Odrv4 I__7153 (
            .O(N__47613),
            .I(\c0.n22_adj_4574 ));
    CascadeMux I__7152 (
            .O(N__47610),
            .I(N__47606));
    CascadeMux I__7151 (
            .O(N__47609),
            .I(N__47603));
    InMux I__7150 (
            .O(N__47606),
            .I(N__47600));
    InMux I__7149 (
            .O(N__47603),
            .I(N__47597));
    LocalMux I__7148 (
            .O(N__47600),
            .I(N__47594));
    LocalMux I__7147 (
            .O(N__47597),
            .I(\c0.data_in_frame_20_1 ));
    Odrv12 I__7146 (
            .O(N__47594),
            .I(\c0.data_in_frame_20_1 ));
    InMux I__7145 (
            .O(N__47589),
            .I(N__47586));
    LocalMux I__7144 (
            .O(N__47586),
            .I(N__47583));
    Span4Mux_h I__7143 (
            .O(N__47583),
            .I(N__47579));
    InMux I__7142 (
            .O(N__47582),
            .I(N__47576));
    Odrv4 I__7141 (
            .O(N__47579),
            .I(\c0.n33945 ));
    LocalMux I__7140 (
            .O(N__47576),
            .I(\c0.n33945 ));
    InMux I__7139 (
            .O(N__47571),
            .I(N__47568));
    LocalMux I__7138 (
            .O(N__47568),
            .I(N__47565));
    Odrv12 I__7137 (
            .O(N__47565),
            .I(\c0.n18431 ));
    InMux I__7136 (
            .O(N__47562),
            .I(N__47558));
    InMux I__7135 (
            .O(N__47561),
            .I(N__47555));
    LocalMux I__7134 (
            .O(N__47558),
            .I(N__47552));
    LocalMux I__7133 (
            .O(N__47555),
            .I(\c0.n33886 ));
    Odrv4 I__7132 (
            .O(N__47552),
            .I(\c0.n33886 ));
    CascadeMux I__7131 (
            .O(N__47547),
            .I(N__47544));
    InMux I__7130 (
            .O(N__47544),
            .I(N__47540));
    CascadeMux I__7129 (
            .O(N__47543),
            .I(N__47537));
    LocalMux I__7128 (
            .O(N__47540),
            .I(N__47533));
    InMux I__7127 (
            .O(N__47537),
            .I(N__47528));
    InMux I__7126 (
            .O(N__47536),
            .I(N__47525));
    Span4Mux_v I__7125 (
            .O(N__47533),
            .I(N__47522));
    InMux I__7124 (
            .O(N__47532),
            .I(N__47519));
    InMux I__7123 (
            .O(N__47531),
            .I(N__47516));
    LocalMux I__7122 (
            .O(N__47528),
            .I(\c0.data_in_frame_17_5 ));
    LocalMux I__7121 (
            .O(N__47525),
            .I(\c0.data_in_frame_17_5 ));
    Odrv4 I__7120 (
            .O(N__47522),
            .I(\c0.data_in_frame_17_5 ));
    LocalMux I__7119 (
            .O(N__47519),
            .I(\c0.data_in_frame_17_5 ));
    LocalMux I__7118 (
            .O(N__47516),
            .I(\c0.data_in_frame_17_5 ));
    InMux I__7117 (
            .O(N__47505),
            .I(N__47502));
    LocalMux I__7116 (
            .O(N__47502),
            .I(\c0.n8_adj_4745 ));
    CascadeMux I__7115 (
            .O(N__47499),
            .I(\c0.n6242_cascade_ ));
    CascadeMux I__7114 (
            .O(N__47496),
            .I(\c0.n33665_cascade_ ));
    CascadeMux I__7113 (
            .O(N__47493),
            .I(N__47490));
    InMux I__7112 (
            .O(N__47490),
            .I(N__47486));
    InMux I__7111 (
            .O(N__47489),
            .I(N__47483));
    LocalMux I__7110 (
            .O(N__47486),
            .I(\c0.data_in_frame_19_0 ));
    LocalMux I__7109 (
            .O(N__47483),
            .I(\c0.data_in_frame_19_0 ));
    CascadeMux I__7108 (
            .O(N__47478),
            .I(N__47475));
    InMux I__7107 (
            .O(N__47475),
            .I(N__47471));
    InMux I__7106 (
            .O(N__47474),
            .I(N__47468));
    LocalMux I__7105 (
            .O(N__47471),
            .I(\c0.data_in_frame_20_0 ));
    LocalMux I__7104 (
            .O(N__47468),
            .I(\c0.data_in_frame_20_0 ));
    CascadeMux I__7103 (
            .O(N__47463),
            .I(N__47460));
    InMux I__7102 (
            .O(N__47460),
            .I(N__47457));
    LocalMux I__7101 (
            .O(N__47457),
            .I(N__47454));
    Span4Mux_h I__7100 (
            .O(N__47454),
            .I(N__47451));
    Odrv4 I__7099 (
            .O(N__47451),
            .I(\c0.n19199 ));
    InMux I__7098 (
            .O(N__47448),
            .I(N__47444));
    InMux I__7097 (
            .O(N__47447),
            .I(N__47441));
    LocalMux I__7096 (
            .O(N__47444),
            .I(\c0.n31589 ));
    LocalMux I__7095 (
            .O(N__47441),
            .I(\c0.n31589 ));
    CascadeMux I__7094 (
            .O(N__47436),
            .I(\c0.n33514_cascade_ ));
    InMux I__7093 (
            .O(N__47433),
            .I(N__47427));
    InMux I__7092 (
            .O(N__47432),
            .I(N__47427));
    LocalMux I__7091 (
            .O(N__47427),
            .I(\c0.n19226 ));
    InMux I__7090 (
            .O(N__47424),
            .I(N__47421));
    LocalMux I__7089 (
            .O(N__47421),
            .I(\c0.n12_adj_4696 ));
    InMux I__7088 (
            .O(N__47418),
            .I(N__47412));
    InMux I__7087 (
            .O(N__47417),
            .I(N__47412));
    LocalMux I__7086 (
            .O(N__47412),
            .I(\c0.n33717 ));
    InMux I__7085 (
            .O(N__47409),
            .I(N__47405));
    InMux I__7084 (
            .O(N__47408),
            .I(N__47402));
    LocalMux I__7083 (
            .O(N__47405),
            .I(N__47399));
    LocalMux I__7082 (
            .O(N__47402),
            .I(\c0.data_in_frame_19_1 ));
    Odrv4 I__7081 (
            .O(N__47399),
            .I(\c0.data_in_frame_19_1 ));
    InMux I__7080 (
            .O(N__47394),
            .I(N__47391));
    LocalMux I__7079 (
            .O(N__47391),
            .I(N__47388));
    Odrv4 I__7078 (
            .O(N__47388),
            .I(\c0.n34003 ));
    InMux I__7077 (
            .O(N__47385),
            .I(N__47382));
    LocalMux I__7076 (
            .O(N__47382),
            .I(\c0.n24_adj_4717 ));
    CascadeMux I__7075 (
            .O(N__47379),
            .I(N__47375));
    InMux I__7074 (
            .O(N__47378),
            .I(N__47369));
    InMux I__7073 (
            .O(N__47375),
            .I(N__47369));
    InMux I__7072 (
            .O(N__47374),
            .I(N__47366));
    LocalMux I__7071 (
            .O(N__47369),
            .I(\c0.data_in_frame_18_0 ));
    LocalMux I__7070 (
            .O(N__47366),
            .I(\c0.data_in_frame_18_0 ));
    InMux I__7069 (
            .O(N__47361),
            .I(N__47357));
    InMux I__7068 (
            .O(N__47360),
            .I(N__47354));
    LocalMux I__7067 (
            .O(N__47357),
            .I(N__47351));
    LocalMux I__7066 (
            .O(N__47354),
            .I(N__47348));
    Span4Mux_v I__7065 (
            .O(N__47351),
            .I(N__47345));
    Odrv4 I__7064 (
            .O(N__47348),
            .I(\c0.n33371 ));
    Odrv4 I__7063 (
            .O(N__47345),
            .I(\c0.n33371 ));
    InMux I__7062 (
            .O(N__47340),
            .I(N__47337));
    LocalMux I__7061 (
            .O(N__47337),
            .I(N__47334));
    Odrv4 I__7060 (
            .O(N__47334),
            .I(\c0.n10_adj_4697 ));
    InMux I__7059 (
            .O(N__47331),
            .I(N__47327));
    InMux I__7058 (
            .O(N__47330),
            .I(N__47324));
    LocalMux I__7057 (
            .O(N__47327),
            .I(\c0.n33356 ));
    LocalMux I__7056 (
            .O(N__47324),
            .I(\c0.n33356 ));
    CascadeMux I__7055 (
            .O(N__47319),
            .I(\c0.n18588_cascade_ ));
    InMux I__7054 (
            .O(N__47316),
            .I(N__47313));
    LocalMux I__7053 (
            .O(N__47313),
            .I(\c0.n33789 ));
    CascadeMux I__7052 (
            .O(N__47310),
            .I(\c0.n33789_cascade_ ));
    CascadeMux I__7051 (
            .O(N__47307),
            .I(\c0.n19108_cascade_ ));
    InMux I__7050 (
            .O(N__47304),
            .I(N__47301));
    LocalMux I__7049 (
            .O(N__47301),
            .I(N__47297));
    CascadeMux I__7048 (
            .O(N__47300),
            .I(N__47294));
    Span4Mux_h I__7047 (
            .O(N__47297),
            .I(N__47291));
    InMux I__7046 (
            .O(N__47294),
            .I(N__47288));
    Span4Mux_h I__7045 (
            .O(N__47291),
            .I(N__47285));
    LocalMux I__7044 (
            .O(N__47288),
            .I(\c0.data_in_frame_18_2 ));
    Odrv4 I__7043 (
            .O(N__47285),
            .I(\c0.data_in_frame_18_2 ));
    CascadeMux I__7042 (
            .O(N__47280),
            .I(\c0.n12_adj_4716_cascade_ ));
    InMux I__7041 (
            .O(N__47277),
            .I(N__47274));
    LocalMux I__7040 (
            .O(N__47274),
            .I(N__47271));
    Span4Mux_v I__7039 (
            .O(N__47271),
            .I(N__47268));
    Odrv4 I__7038 (
            .O(N__47268),
            .I(\c0.n33741 ));
    InMux I__7037 (
            .O(N__47265),
            .I(N__47259));
    InMux I__7036 (
            .O(N__47264),
            .I(N__47259));
    LocalMux I__7035 (
            .O(N__47259),
            .I(N__47256));
    Span4Mux_h I__7034 (
            .O(N__47256),
            .I(N__47253));
    Span4Mux_h I__7033 (
            .O(N__47253),
            .I(N__47250));
    Odrv4 I__7032 (
            .O(N__47250),
            .I(\c0.n18368 ));
    CascadeMux I__7031 (
            .O(N__47247),
            .I(\c0.n33741_cascade_ ));
    InMux I__7030 (
            .O(N__47244),
            .I(N__47241));
    LocalMux I__7029 (
            .O(N__47241),
            .I(\c0.n33880 ));
    CascadeMux I__7028 (
            .O(N__47238),
            .I(N__47234));
    InMux I__7027 (
            .O(N__47237),
            .I(N__47230));
    InMux I__7026 (
            .O(N__47234),
            .I(N__47225));
    InMux I__7025 (
            .O(N__47233),
            .I(N__47225));
    LocalMux I__7024 (
            .O(N__47230),
            .I(\c0.data_in_frame_17_7 ));
    LocalMux I__7023 (
            .O(N__47225),
            .I(\c0.data_in_frame_17_7 ));
    InMux I__7022 (
            .O(N__47220),
            .I(N__47216));
    InMux I__7021 (
            .O(N__47219),
            .I(N__47213));
    LocalMux I__7020 (
            .O(N__47216),
            .I(\c0.n33711 ));
    LocalMux I__7019 (
            .O(N__47213),
            .I(\c0.n33711 ));
    InMux I__7018 (
            .O(N__47208),
            .I(N__47204));
    InMux I__7017 (
            .O(N__47207),
            .I(N__47201));
    LocalMux I__7016 (
            .O(N__47204),
            .I(N__47196));
    LocalMux I__7015 (
            .O(N__47201),
            .I(N__47196));
    Odrv12 I__7014 (
            .O(N__47196),
            .I(\c0.n5896 ));
    CascadeMux I__7013 (
            .O(N__47193),
            .I(\c0.n34_adj_4718_cascade_ ));
    InMux I__7012 (
            .O(N__47190),
            .I(N__47187));
    LocalMux I__7011 (
            .O(N__47187),
            .I(N__47184));
    Span4Mux_h I__7010 (
            .O(N__47184),
            .I(N__47181));
    Odrv4 I__7009 (
            .O(N__47181),
            .I(\c0.n37_adj_4720 ));
    InMux I__7008 (
            .O(N__47178),
            .I(N__47175));
    LocalMux I__7007 (
            .O(N__47175),
            .I(\c0.n35_adj_4721 ));
    CascadeMux I__7006 (
            .O(N__47172),
            .I(\c0.n38_adj_4719_cascade_ ));
    CascadeMux I__7005 (
            .O(N__47169),
            .I(N__47165));
    InMux I__7004 (
            .O(N__47168),
            .I(N__47161));
    InMux I__7003 (
            .O(N__47165),
            .I(N__47158));
    InMux I__7002 (
            .O(N__47164),
            .I(N__47155));
    LocalMux I__7001 (
            .O(N__47161),
            .I(N__47152));
    LocalMux I__7000 (
            .O(N__47158),
            .I(\c0.data_in_frame_16_1 ));
    LocalMux I__6999 (
            .O(N__47155),
            .I(\c0.data_in_frame_16_1 ));
    Odrv4 I__6998 (
            .O(N__47152),
            .I(\c0.data_in_frame_16_1 ));
    CascadeMux I__6997 (
            .O(N__47145),
            .I(\c0.n2_adj_4741_cascade_ ));
    InMux I__6996 (
            .O(N__47142),
            .I(N__47136));
    InMux I__6995 (
            .O(N__47141),
            .I(N__47136));
    LocalMux I__6994 (
            .O(N__47136),
            .I(N__47133));
    Span4Mux_v I__6993 (
            .O(N__47133),
            .I(N__47130));
    Odrv4 I__6992 (
            .O(N__47130),
            .I(\c0.n33283 ));
    CascadeMux I__6991 (
            .O(N__47127),
            .I(N__47124));
    InMux I__6990 (
            .O(N__47124),
            .I(N__47117));
    InMux I__6989 (
            .O(N__47123),
            .I(N__47117));
    InMux I__6988 (
            .O(N__47122),
            .I(N__47114));
    LocalMux I__6987 (
            .O(N__47117),
            .I(N__47111));
    LocalMux I__6986 (
            .O(N__47114),
            .I(\c0.data_in_frame_8_1 ));
    Odrv4 I__6985 (
            .O(N__47111),
            .I(\c0.data_in_frame_8_1 ));
    CascadeMux I__6984 (
            .O(N__47106),
            .I(\c0.n33283_cascade_ ));
    InMux I__6983 (
            .O(N__47103),
            .I(N__47099));
    InMux I__6982 (
            .O(N__47102),
            .I(N__47096));
    LocalMux I__6981 (
            .O(N__47099),
            .I(N__47093));
    LocalMux I__6980 (
            .O(N__47096),
            .I(N__47090));
    Span4Mux_v I__6979 (
            .O(N__47093),
            .I(N__47087));
    Odrv4 I__6978 (
            .O(N__47090),
            .I(\c0.n33871 ));
    Odrv4 I__6977 (
            .O(N__47087),
            .I(\c0.n33871 ));
    CascadeMux I__6976 (
            .O(N__47082),
            .I(N__47079));
    InMux I__6975 (
            .O(N__47079),
            .I(N__47073));
    InMux I__6974 (
            .O(N__47078),
            .I(N__47073));
    LocalMux I__6973 (
            .O(N__47073),
            .I(\c0.data_in_frame_18_3 ));
    CascadeMux I__6972 (
            .O(N__47070),
            .I(N__47066));
    InMux I__6971 (
            .O(N__47069),
            .I(N__47063));
    InMux I__6970 (
            .O(N__47066),
            .I(N__47059));
    LocalMux I__6969 (
            .O(N__47063),
            .I(N__47056));
    CascadeMux I__6968 (
            .O(N__47062),
            .I(N__47053));
    LocalMux I__6967 (
            .O(N__47059),
            .I(N__47050));
    Span4Mux_h I__6966 (
            .O(N__47056),
            .I(N__47047));
    InMux I__6965 (
            .O(N__47053),
            .I(N__47044));
    Odrv4 I__6964 (
            .O(N__47050),
            .I(\c0.data_in_frame_14_5 ));
    Odrv4 I__6963 (
            .O(N__47047),
            .I(\c0.data_in_frame_14_5 ));
    LocalMux I__6962 (
            .O(N__47044),
            .I(\c0.data_in_frame_14_5 ));
    CascadeMux I__6961 (
            .O(N__47037),
            .I(N__47033));
    CascadeMux I__6960 (
            .O(N__47036),
            .I(N__47030));
    InMux I__6959 (
            .O(N__47033),
            .I(N__47025));
    InMux I__6958 (
            .O(N__47030),
            .I(N__47025));
    LocalMux I__6957 (
            .O(N__47025),
            .I(\c0.data_in_frame_6_1 ));
    InMux I__6956 (
            .O(N__47022),
            .I(N__47019));
    LocalMux I__6955 (
            .O(N__47019),
            .I(N__47016));
    Odrv12 I__6954 (
            .O(N__47016),
            .I(\c0.n18364 ));
    CascadeMux I__6953 (
            .O(N__47013),
            .I(\c0.n33880_cascade_ ));
    CascadeMux I__6952 (
            .O(N__47010),
            .I(\c0.n33927_cascade_ ));
    CascadeMux I__6951 (
            .O(N__47007),
            .I(N__47004));
    InMux I__6950 (
            .O(N__47004),
            .I(N__46998));
    InMux I__6949 (
            .O(N__47003),
            .I(N__46998));
    LocalMux I__6948 (
            .O(N__46998),
            .I(\c0.data_in_frame_10_2 ));
    InMux I__6947 (
            .O(N__46995),
            .I(N__46991));
    CascadeMux I__6946 (
            .O(N__46994),
            .I(N__46987));
    LocalMux I__6945 (
            .O(N__46991),
            .I(N__46983));
    InMux I__6944 (
            .O(N__46990),
            .I(N__46980));
    InMux I__6943 (
            .O(N__46987),
            .I(N__46975));
    InMux I__6942 (
            .O(N__46986),
            .I(N__46975));
    Odrv12 I__6941 (
            .O(N__46983),
            .I(\c0.n31439 ));
    LocalMux I__6940 (
            .O(N__46980),
            .I(\c0.n31439 ));
    LocalMux I__6939 (
            .O(N__46975),
            .I(\c0.n31439 ));
    CascadeMux I__6938 (
            .O(N__46968),
            .I(N__46964));
    InMux I__6937 (
            .O(N__46967),
            .I(N__46961));
    InMux I__6936 (
            .O(N__46964),
            .I(N__46958));
    LocalMux I__6935 (
            .O(N__46961),
            .I(N__46955));
    LocalMux I__6934 (
            .O(N__46958),
            .I(\c0.data_in_frame_14_1 ));
    Odrv4 I__6933 (
            .O(N__46955),
            .I(\c0.data_in_frame_14_1 ));
    InMux I__6932 (
            .O(N__46950),
            .I(N__46947));
    LocalMux I__6931 (
            .O(N__46947),
            .I(N__46944));
    Odrv12 I__6930 (
            .O(N__46944),
            .I(\c0.n2_adj_4741 ));
    InMux I__6929 (
            .O(N__46941),
            .I(N__46937));
    InMux I__6928 (
            .O(N__46940),
            .I(N__46932));
    LocalMux I__6927 (
            .O(N__46937),
            .I(N__46929));
    InMux I__6926 (
            .O(N__46936),
            .I(N__46925));
    InMux I__6925 (
            .O(N__46935),
            .I(N__46922));
    LocalMux I__6924 (
            .O(N__46932),
            .I(N__46919));
    Span4Mux_v I__6923 (
            .O(N__46929),
            .I(N__46915));
    InMux I__6922 (
            .O(N__46928),
            .I(N__46912));
    LocalMux I__6921 (
            .O(N__46925),
            .I(N__46909));
    LocalMux I__6920 (
            .O(N__46922),
            .I(N__46906));
    Span4Mux_h I__6919 (
            .O(N__46919),
            .I(N__46903));
    InMux I__6918 (
            .O(N__46918),
            .I(N__46900));
    Span4Mux_h I__6917 (
            .O(N__46915),
            .I(N__46897));
    LocalMux I__6916 (
            .O(N__46912),
            .I(N__46892));
    Span4Mux_v I__6915 (
            .O(N__46909),
            .I(N__46892));
    Span4Mux_h I__6914 (
            .O(N__46906),
            .I(N__46889));
    Span4Mux_h I__6913 (
            .O(N__46903),
            .I(N__46886));
    LocalMux I__6912 (
            .O(N__46900),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__6911 (
            .O(N__46897),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__6910 (
            .O(N__46892),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__6909 (
            .O(N__46889),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__6908 (
            .O(N__46886),
            .I(\c0.data_in_frame_6_7 ));
    CascadeMux I__6907 (
            .O(N__46875),
            .I(\c0.n6_adj_4501_cascade_ ));
    InMux I__6906 (
            .O(N__46872),
            .I(N__46869));
    LocalMux I__6905 (
            .O(N__46869),
            .I(N__46865));
    CascadeMux I__6904 (
            .O(N__46868),
            .I(N__46861));
    Span4Mux_h I__6903 (
            .O(N__46865),
            .I(N__46858));
    InMux I__6902 (
            .O(N__46864),
            .I(N__46855));
    InMux I__6901 (
            .O(N__46861),
            .I(N__46852));
    Span4Mux_v I__6900 (
            .O(N__46858),
            .I(N__46849));
    LocalMux I__6899 (
            .O(N__46855),
            .I(N__46846));
    LocalMux I__6898 (
            .O(N__46852),
            .I(\c0.data_in_frame_3_2 ));
    Odrv4 I__6897 (
            .O(N__46849),
            .I(\c0.data_in_frame_3_2 ));
    Odrv12 I__6896 (
            .O(N__46846),
            .I(\c0.data_in_frame_3_2 ));
    CascadeMux I__6895 (
            .O(N__46839),
            .I(N__46836));
    InMux I__6894 (
            .O(N__46836),
            .I(N__46832));
    InMux I__6893 (
            .O(N__46835),
            .I(N__46829));
    LocalMux I__6892 (
            .O(N__46832),
            .I(\c0.data_in_frame_5_5 ));
    LocalMux I__6891 (
            .O(N__46829),
            .I(\c0.data_in_frame_5_5 ));
    CascadeMux I__6890 (
            .O(N__46824),
            .I(\c0.n6_cascade_ ));
    CascadeMux I__6889 (
            .O(N__46821),
            .I(\c0.n18141_cascade_ ));
    InMux I__6888 (
            .O(N__46818),
            .I(N__46815));
    LocalMux I__6887 (
            .O(N__46815),
            .I(N__46809));
    InMux I__6886 (
            .O(N__46814),
            .I(N__46804));
    InMux I__6885 (
            .O(N__46813),
            .I(N__46804));
    InMux I__6884 (
            .O(N__46812),
            .I(N__46801));
    Odrv12 I__6883 (
            .O(N__46809),
            .I(\c0.data_in_frame_3_3 ));
    LocalMux I__6882 (
            .O(N__46804),
            .I(\c0.data_in_frame_3_3 ));
    LocalMux I__6881 (
            .O(N__46801),
            .I(\c0.data_in_frame_3_3 ));
    InMux I__6880 (
            .O(N__46794),
            .I(N__46790));
    InMux I__6879 (
            .O(N__46793),
            .I(N__46786));
    LocalMux I__6878 (
            .O(N__46790),
            .I(N__46782));
    InMux I__6877 (
            .O(N__46789),
            .I(N__46779));
    LocalMux I__6876 (
            .O(N__46786),
            .I(N__46776));
    InMux I__6875 (
            .O(N__46785),
            .I(N__46773));
    Span4Mux_v I__6874 (
            .O(N__46782),
            .I(N__46770));
    LocalMux I__6873 (
            .O(N__46779),
            .I(N__46765));
    Span4Mux_h I__6872 (
            .O(N__46776),
            .I(N__46765));
    LocalMux I__6871 (
            .O(N__46773),
            .I(\c0.data_in_frame_2_7 ));
    Odrv4 I__6870 (
            .O(N__46770),
            .I(\c0.data_in_frame_2_7 ));
    Odrv4 I__6869 (
            .O(N__46765),
            .I(\c0.data_in_frame_2_7 ));
    InMux I__6868 (
            .O(N__46758),
            .I(N__46755));
    LocalMux I__6867 (
            .O(N__46755),
            .I(\c0.n39_adj_4781 ));
    InMux I__6866 (
            .O(N__46752),
            .I(N__46749));
    LocalMux I__6865 (
            .O(N__46749),
            .I(\c0.n37_adj_4782 ));
    InMux I__6864 (
            .O(N__46746),
            .I(N__46737));
    CascadeMux I__6863 (
            .O(N__46745),
            .I(N__46734));
    CascadeMux I__6862 (
            .O(N__46744),
            .I(N__46731));
    InMux I__6861 (
            .O(N__46743),
            .I(N__46726));
    InMux I__6860 (
            .O(N__46742),
            .I(N__46726));
    InMux I__6859 (
            .O(N__46741),
            .I(N__46721));
    InMux I__6858 (
            .O(N__46740),
            .I(N__46721));
    LocalMux I__6857 (
            .O(N__46737),
            .I(N__46717));
    InMux I__6856 (
            .O(N__46734),
            .I(N__46714));
    InMux I__6855 (
            .O(N__46731),
            .I(N__46711));
    LocalMux I__6854 (
            .O(N__46726),
            .I(N__46706));
    LocalMux I__6853 (
            .O(N__46721),
            .I(N__46706));
    InMux I__6852 (
            .O(N__46720),
            .I(N__46703));
    Span4Mux_v I__6851 (
            .O(N__46717),
            .I(N__46698));
    LocalMux I__6850 (
            .O(N__46714),
            .I(N__46698));
    LocalMux I__6849 (
            .O(N__46711),
            .I(\c0.data_in_frame_0_5 ));
    Odrv4 I__6848 (
            .O(N__46706),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__6847 (
            .O(N__46703),
            .I(\c0.data_in_frame_0_5 ));
    Odrv4 I__6846 (
            .O(N__46698),
            .I(\c0.data_in_frame_0_5 ));
    InMux I__6845 (
            .O(N__46689),
            .I(N__46686));
    LocalMux I__6844 (
            .O(N__46686),
            .I(N__46683));
    Span4Mux_h I__6843 (
            .O(N__46683),
            .I(N__46680));
    Odrv4 I__6842 (
            .O(N__46680),
            .I(\c0.n10_adj_4768 ));
    InMux I__6841 (
            .O(N__46677),
            .I(N__46674));
    LocalMux I__6840 (
            .O(N__46674),
            .I(N__46671));
    Span4Mux_v I__6839 (
            .O(N__46671),
            .I(N__46668));
    Span4Mux_h I__6838 (
            .O(N__46668),
            .I(N__46662));
    InMux I__6837 (
            .O(N__46667),
            .I(N__46659));
    InMux I__6836 (
            .O(N__46666),
            .I(N__46654));
    InMux I__6835 (
            .O(N__46665),
            .I(N__46654));
    Odrv4 I__6834 (
            .O(N__46662),
            .I(n18026));
    LocalMux I__6833 (
            .O(N__46659),
            .I(n18026));
    LocalMux I__6832 (
            .O(N__46654),
            .I(n18026));
    InMux I__6831 (
            .O(N__46647),
            .I(N__46641));
    InMux I__6830 (
            .O(N__46646),
            .I(N__46638));
    CascadeMux I__6829 (
            .O(N__46645),
            .I(N__46635));
    InMux I__6828 (
            .O(N__46644),
            .I(N__46632));
    LocalMux I__6827 (
            .O(N__46641),
            .I(N__46629));
    LocalMux I__6826 (
            .O(N__46638),
            .I(N__46626));
    InMux I__6825 (
            .O(N__46635),
            .I(N__46622));
    LocalMux I__6824 (
            .O(N__46632),
            .I(N__46619));
    Span4Mux_v I__6823 (
            .O(N__46629),
            .I(N__46615));
    Span4Mux_v I__6822 (
            .O(N__46626),
            .I(N__46612));
    InMux I__6821 (
            .O(N__46625),
            .I(N__46609));
    LocalMux I__6820 (
            .O(N__46622),
            .I(N__46604));
    Span4Mux_v I__6819 (
            .O(N__46619),
            .I(N__46604));
    InMux I__6818 (
            .O(N__46618),
            .I(N__46601));
    Span4Mux_h I__6817 (
            .O(N__46615),
            .I(N__46598));
    Span4Mux_v I__6816 (
            .O(N__46612),
            .I(N__46595));
    LocalMux I__6815 (
            .O(N__46609),
            .I(N__46592));
    Span4Mux_h I__6814 (
            .O(N__46604),
            .I(N__46589));
    LocalMux I__6813 (
            .O(N__46601),
            .I(\c0.data_in_frame_6_6 ));
    Odrv4 I__6812 (
            .O(N__46598),
            .I(\c0.data_in_frame_6_6 ));
    Odrv4 I__6811 (
            .O(N__46595),
            .I(\c0.data_in_frame_6_6 ));
    Odrv4 I__6810 (
            .O(N__46592),
            .I(\c0.data_in_frame_6_6 ));
    Odrv4 I__6809 (
            .O(N__46589),
            .I(\c0.data_in_frame_6_6 ));
    CascadeMux I__6808 (
            .O(N__46578),
            .I(N__46575));
    InMux I__6807 (
            .O(N__46575),
            .I(N__46572));
    LocalMux I__6806 (
            .O(N__46572),
            .I(N__46569));
    Odrv12 I__6805 (
            .O(N__46569),
            .I(\c0.data_out_frame_0__7__N_2747 ));
    InMux I__6804 (
            .O(N__46566),
            .I(N__46563));
    LocalMux I__6803 (
            .O(N__46563),
            .I(N__46560));
    Odrv4 I__6802 (
            .O(N__46560),
            .I(\c0.n26_adj_4775 ));
    CascadeMux I__6801 (
            .O(N__46557),
            .I(N__46553));
    InMux I__6800 (
            .O(N__46556),
            .I(N__46550));
    InMux I__6799 (
            .O(N__46553),
            .I(N__46547));
    LocalMux I__6798 (
            .O(N__46550),
            .I(\c0.n33582 ));
    LocalMux I__6797 (
            .O(N__46547),
            .I(\c0.n33582 ));
    CascadeMux I__6796 (
            .O(N__46542),
            .I(\c0.n33291_cascade_ ));
    InMux I__6795 (
            .O(N__46539),
            .I(N__46536));
    LocalMux I__6794 (
            .O(N__46536),
            .I(N__46533));
    Odrv4 I__6793 (
            .O(N__46533),
            .I(\c0.n19_adj_4779 ));
    InMux I__6792 (
            .O(N__46530),
            .I(N__46525));
    CascadeMux I__6791 (
            .O(N__46529),
            .I(N__46521));
    InMux I__6790 (
            .O(N__46528),
            .I(N__46518));
    LocalMux I__6789 (
            .O(N__46525),
            .I(N__46515));
    InMux I__6788 (
            .O(N__46524),
            .I(N__46512));
    InMux I__6787 (
            .O(N__46521),
            .I(N__46509));
    LocalMux I__6786 (
            .O(N__46518),
            .I(N__46506));
    Span4Mux_h I__6785 (
            .O(N__46515),
            .I(N__46503));
    LocalMux I__6784 (
            .O(N__46512),
            .I(N__46500));
    LocalMux I__6783 (
            .O(N__46509),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__6782 (
            .O(N__46506),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__6781 (
            .O(N__46503),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__6780 (
            .O(N__46500),
            .I(\c0.data_in_frame_2_6 ));
    CascadeMux I__6779 (
            .O(N__46491),
            .I(N__46487));
    InMux I__6778 (
            .O(N__46490),
            .I(N__46482));
    InMux I__6777 (
            .O(N__46487),
            .I(N__46482));
    LocalMux I__6776 (
            .O(N__46482),
            .I(\c0.data_in_frame_5_6 ));
    InMux I__6775 (
            .O(N__46479),
            .I(N__46476));
    LocalMux I__6774 (
            .O(N__46476),
            .I(N__46473));
    Odrv4 I__6773 (
            .O(N__46473),
            .I(\c0.n29_adj_4776 ));
    CascadeMux I__6772 (
            .O(N__46470),
            .I(N__46467));
    InMux I__6771 (
            .O(N__46467),
            .I(N__46464));
    LocalMux I__6770 (
            .O(N__46464),
            .I(N__46460));
    InMux I__6769 (
            .O(N__46463),
            .I(N__46457));
    Span4Mux_h I__6768 (
            .O(N__46460),
            .I(N__46454));
    LocalMux I__6767 (
            .O(N__46457),
            .I(N__46451));
    Span4Mux_h I__6766 (
            .O(N__46454),
            .I(N__46448));
    Span4Mux_h I__6765 (
            .O(N__46451),
            .I(N__46445));
    Odrv4 I__6764 (
            .O(N__46448),
            .I(\c0.n9_adj_4509 ));
    Odrv4 I__6763 (
            .O(N__46445),
            .I(\c0.n9_adj_4509 ));
    InMux I__6762 (
            .O(N__46440),
            .I(N__46437));
    LocalMux I__6761 (
            .O(N__46437),
            .I(N__46434));
    Span4Mux_v I__6760 (
            .O(N__46434),
            .I(N__46431));
    Odrv4 I__6759 (
            .O(N__46431),
            .I(\c0.n34 ));
    InMux I__6758 (
            .O(N__46428),
            .I(N__46425));
    LocalMux I__6757 (
            .O(N__46425),
            .I(N__46420));
    InMux I__6756 (
            .O(N__46424),
            .I(N__46415));
    InMux I__6755 (
            .O(N__46423),
            .I(N__46415));
    Span12Mux_v I__6754 (
            .O(N__46420),
            .I(N__46410));
    LocalMux I__6753 (
            .O(N__46415),
            .I(N__46407));
    InMux I__6752 (
            .O(N__46414),
            .I(N__46404));
    InMux I__6751 (
            .O(N__46413),
            .I(N__46401));
    Odrv12 I__6750 (
            .O(N__46410),
            .I(\c0.n18330 ));
    Odrv4 I__6749 (
            .O(N__46407),
            .I(\c0.n18330 ));
    LocalMux I__6748 (
            .O(N__46404),
            .I(\c0.n18330 ));
    LocalMux I__6747 (
            .O(N__46401),
            .I(\c0.n18330 ));
    InMux I__6746 (
            .O(N__46392),
            .I(N__46389));
    LocalMux I__6745 (
            .O(N__46389),
            .I(N__46386));
    Odrv4 I__6744 (
            .O(N__46386),
            .I(\c0.n20_adj_4534 ));
    CascadeMux I__6743 (
            .O(N__46383),
            .I(\c0.n28_adj_4777_cascade_ ));
    InMux I__6742 (
            .O(N__46380),
            .I(N__46377));
    LocalMux I__6741 (
            .O(N__46377),
            .I(\c0.n32_adj_4778 ));
    CascadeMux I__6740 (
            .O(N__46374),
            .I(\c0.n27710_cascade_ ));
    CascadeMux I__6739 (
            .O(N__46371),
            .I(\c0.n35947_cascade_ ));
    InMux I__6738 (
            .O(N__46368),
            .I(N__46365));
    LocalMux I__6737 (
            .O(N__46365),
            .I(N__46362));
    Span4Mux_v I__6736 (
            .O(N__46362),
            .I(N__46359));
    Odrv4 I__6735 (
            .O(N__46359),
            .I(\c0.n35808 ));
    CascadeMux I__6734 (
            .O(N__46356),
            .I(\c0.n38_adj_4780_cascade_ ));
    InMux I__6733 (
            .O(N__46353),
            .I(N__46350));
    LocalMux I__6732 (
            .O(N__46350),
            .I(\c0.n35804 ));
    CascadeMux I__6731 (
            .O(N__46347),
            .I(\c0.n46_adj_4783_cascade_ ));
    SRMux I__6730 (
            .O(N__46344),
            .I(N__46341));
    LocalMux I__6729 (
            .O(N__46341),
            .I(N__46338));
    Span4Mux_v I__6728 (
            .O(N__46338),
            .I(N__46335));
    Odrv4 I__6727 (
            .O(N__46335),
            .I(\c0.n32740 ));
    InMux I__6726 (
            .O(N__46332),
            .I(N__46328));
    CascadeMux I__6725 (
            .O(N__46331),
            .I(N__46324));
    LocalMux I__6724 (
            .O(N__46328),
            .I(N__46320));
    InMux I__6723 (
            .O(N__46327),
            .I(N__46313));
    InMux I__6722 (
            .O(N__46324),
            .I(N__46313));
    InMux I__6721 (
            .O(N__46323),
            .I(N__46313));
    Odrv12 I__6720 (
            .O(N__46320),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__6719 (
            .O(N__46313),
            .I(\c0.FRAME_MATCHER_state_10 ));
    InMux I__6718 (
            .O(N__46308),
            .I(N__46304));
    InMux I__6717 (
            .O(N__46307),
            .I(N__46301));
    LocalMux I__6716 (
            .O(N__46304),
            .I(N__46297));
    LocalMux I__6715 (
            .O(N__46301),
            .I(N__46294));
    CascadeMux I__6714 (
            .O(N__46300),
            .I(N__46290));
    Span4Mux_v I__6713 (
            .O(N__46297),
            .I(N__46285));
    Span4Mux_v I__6712 (
            .O(N__46294),
            .I(N__46285));
    InMux I__6711 (
            .O(N__46293),
            .I(N__46282));
    InMux I__6710 (
            .O(N__46290),
            .I(N__46279));
    Sp12to4 I__6709 (
            .O(N__46285),
            .I(N__46276));
    LocalMux I__6708 (
            .O(N__46282),
            .I(\c0.FRAME_MATCHER_state_12 ));
    LocalMux I__6707 (
            .O(N__46279),
            .I(\c0.FRAME_MATCHER_state_12 ));
    Odrv12 I__6706 (
            .O(N__46276),
            .I(\c0.FRAME_MATCHER_state_12 ));
    CascadeMux I__6705 (
            .O(N__46269),
            .I(N__46266));
    InMux I__6704 (
            .O(N__46266),
            .I(N__46262));
    InMux I__6703 (
            .O(N__46265),
            .I(N__46259));
    LocalMux I__6702 (
            .O(N__46262),
            .I(N__46254));
    LocalMux I__6701 (
            .O(N__46259),
            .I(N__46254));
    Span12Mux_h I__6700 (
            .O(N__46254),
            .I(N__46251));
    Odrv12 I__6699 (
            .O(N__46251),
            .I(\c0.n33160 ));
    CascadeMux I__6698 (
            .O(N__46248),
            .I(\c0.n19909_cascade_ ));
    InMux I__6697 (
            .O(N__46245),
            .I(N__46242));
    LocalMux I__6696 (
            .O(N__46242),
            .I(N__46238));
    InMux I__6695 (
            .O(N__46241),
            .I(N__46235));
    Span4Mux_h I__6694 (
            .O(N__46238),
            .I(N__46232));
    LocalMux I__6693 (
            .O(N__46235),
            .I(N__46228));
    Span4Mux_h I__6692 (
            .O(N__46232),
            .I(N__46225));
    InMux I__6691 (
            .O(N__46231),
            .I(N__46222));
    Odrv4 I__6690 (
            .O(N__46228),
            .I(\c0.data_out_frame_29_7_N_2879_2 ));
    Odrv4 I__6689 (
            .O(N__46225),
            .I(\c0.data_out_frame_29_7_N_2879_2 ));
    LocalMux I__6688 (
            .O(N__46222),
            .I(\c0.data_out_frame_29_7_N_2879_2 ));
    CascadeMux I__6687 (
            .O(N__46215),
            .I(\c0.n34017_cascade_ ));
    CascadeMux I__6686 (
            .O(N__46212),
            .I(\c0.n29675_cascade_ ));
    CascadeMux I__6685 (
            .O(N__46209),
            .I(\c0.n81_cascade_ ));
    InMux I__6684 (
            .O(N__46206),
            .I(N__46170));
    InMux I__6683 (
            .O(N__46205),
            .I(N__46170));
    InMux I__6682 (
            .O(N__46204),
            .I(N__46170));
    InMux I__6681 (
            .O(N__46203),
            .I(N__46170));
    InMux I__6680 (
            .O(N__46202),
            .I(N__46170));
    InMux I__6679 (
            .O(N__46201),
            .I(N__46163));
    InMux I__6678 (
            .O(N__46200),
            .I(N__46163));
    InMux I__6677 (
            .O(N__46199),
            .I(N__46163));
    InMux I__6676 (
            .O(N__46198),
            .I(N__46154));
    InMux I__6675 (
            .O(N__46197),
            .I(N__46154));
    InMux I__6674 (
            .O(N__46196),
            .I(N__46154));
    InMux I__6673 (
            .O(N__46195),
            .I(N__46154));
    InMux I__6672 (
            .O(N__46194),
            .I(N__46149));
    InMux I__6671 (
            .O(N__46193),
            .I(N__46149));
    InMux I__6670 (
            .O(N__46192),
            .I(N__46145));
    InMux I__6669 (
            .O(N__46191),
            .I(N__46142));
    InMux I__6668 (
            .O(N__46190),
            .I(N__46129));
    InMux I__6667 (
            .O(N__46189),
            .I(N__46129));
    InMux I__6666 (
            .O(N__46188),
            .I(N__46129));
    InMux I__6665 (
            .O(N__46187),
            .I(N__46129));
    InMux I__6664 (
            .O(N__46186),
            .I(N__46129));
    InMux I__6663 (
            .O(N__46185),
            .I(N__46129));
    InMux I__6662 (
            .O(N__46184),
            .I(N__46124));
    InMux I__6661 (
            .O(N__46183),
            .I(N__46124));
    InMux I__6660 (
            .O(N__46182),
            .I(N__46119));
    InMux I__6659 (
            .O(N__46181),
            .I(N__46119));
    LocalMux I__6658 (
            .O(N__46170),
            .I(N__46116));
    LocalMux I__6657 (
            .O(N__46163),
            .I(N__46109));
    LocalMux I__6656 (
            .O(N__46154),
            .I(N__46109));
    LocalMux I__6655 (
            .O(N__46149),
            .I(N__46109));
    InMux I__6654 (
            .O(N__46148),
            .I(N__46106));
    LocalMux I__6653 (
            .O(N__46145),
            .I(N__46101));
    LocalMux I__6652 (
            .O(N__46142),
            .I(N__46101));
    LocalMux I__6651 (
            .O(N__46129),
            .I(N__46098));
    LocalMux I__6650 (
            .O(N__46124),
            .I(N__46095));
    LocalMux I__6649 (
            .O(N__46119),
            .I(N__46088));
    Span4Mux_v I__6648 (
            .O(N__46116),
            .I(N__46088));
    Span4Mux_h I__6647 (
            .O(N__46109),
            .I(N__46088));
    LocalMux I__6646 (
            .O(N__46106),
            .I(N__46085));
    Span4Mux_v I__6645 (
            .O(N__46101),
            .I(N__46082));
    Span12Mux_s9_h I__6644 (
            .O(N__46098),
            .I(N__46079));
    Span4Mux_h I__6643 (
            .O(N__46095),
            .I(N__46076));
    Span4Mux_h I__6642 (
            .O(N__46088),
            .I(N__46073));
    Odrv12 I__6641 (
            .O(N__46085),
            .I(\c0.n99 ));
    Odrv4 I__6640 (
            .O(N__46082),
            .I(\c0.n99 ));
    Odrv12 I__6639 (
            .O(N__46079),
            .I(\c0.n99 ));
    Odrv4 I__6638 (
            .O(N__46076),
            .I(\c0.n99 ));
    Odrv4 I__6637 (
            .O(N__46073),
            .I(\c0.n99 ));
    CascadeMux I__6636 (
            .O(N__46062),
            .I(N__46055));
    InMux I__6635 (
            .O(N__46061),
            .I(N__46050));
    CascadeMux I__6634 (
            .O(N__46060),
            .I(N__46042));
    CascadeMux I__6633 (
            .O(N__46059),
            .I(N__46039));
    InMux I__6632 (
            .O(N__46058),
            .I(N__46033));
    InMux I__6631 (
            .O(N__46055),
            .I(N__46033));
    CascadeMux I__6630 (
            .O(N__46054),
            .I(N__46023));
    CascadeMux I__6629 (
            .O(N__46053),
            .I(N__46020));
    LocalMux I__6628 (
            .O(N__46050),
            .I(N__46016));
    InMux I__6627 (
            .O(N__46049),
            .I(N__46005));
    InMux I__6626 (
            .O(N__46048),
            .I(N__46005));
    InMux I__6625 (
            .O(N__46047),
            .I(N__46005));
    InMux I__6624 (
            .O(N__46046),
            .I(N__46005));
    InMux I__6623 (
            .O(N__46045),
            .I(N__46005));
    InMux I__6622 (
            .O(N__46042),
            .I(N__45998));
    InMux I__6621 (
            .O(N__46039),
            .I(N__45998));
    InMux I__6620 (
            .O(N__46038),
            .I(N__45998));
    LocalMux I__6619 (
            .O(N__46033),
            .I(N__45995));
    CascadeMux I__6618 (
            .O(N__46032),
            .I(N__45992));
    CascadeMux I__6617 (
            .O(N__46031),
            .I(N__45988));
    InMux I__6616 (
            .O(N__46030),
            .I(N__45982));
    InMux I__6615 (
            .O(N__46029),
            .I(N__45975));
    InMux I__6614 (
            .O(N__46028),
            .I(N__45975));
    InMux I__6613 (
            .O(N__46027),
            .I(N__45975));
    InMux I__6612 (
            .O(N__46026),
            .I(N__45966));
    InMux I__6611 (
            .O(N__46023),
            .I(N__45966));
    InMux I__6610 (
            .O(N__46020),
            .I(N__45966));
    InMux I__6609 (
            .O(N__46019),
            .I(N__45966));
    Span4Mux_v I__6608 (
            .O(N__46016),
            .I(N__45963));
    LocalMux I__6607 (
            .O(N__46005),
            .I(N__45958));
    LocalMux I__6606 (
            .O(N__45998),
            .I(N__45958));
    Span4Mux_h I__6605 (
            .O(N__45995),
            .I(N__45955));
    InMux I__6604 (
            .O(N__45992),
            .I(N__45944));
    InMux I__6603 (
            .O(N__45991),
            .I(N__45944));
    InMux I__6602 (
            .O(N__45988),
            .I(N__45944));
    InMux I__6601 (
            .O(N__45987),
            .I(N__45944));
    InMux I__6600 (
            .O(N__45986),
            .I(N__45944));
    InMux I__6599 (
            .O(N__45985),
            .I(N__45941));
    LocalMux I__6598 (
            .O(N__45982),
            .I(N__45938));
    LocalMux I__6597 (
            .O(N__45975),
            .I(N__45933));
    LocalMux I__6596 (
            .O(N__45966),
            .I(N__45933));
    Span4Mux_h I__6595 (
            .O(N__45963),
            .I(N__45926));
    Span4Mux_v I__6594 (
            .O(N__45958),
            .I(N__45926));
    Span4Mux_h I__6593 (
            .O(N__45955),
            .I(N__45926));
    LocalMux I__6592 (
            .O(N__45944),
            .I(\c0.n3_adj_4636 ));
    LocalMux I__6591 (
            .O(N__45941),
            .I(\c0.n3_adj_4636 ));
    Odrv4 I__6590 (
            .O(N__45938),
            .I(\c0.n3_adj_4636 ));
    Odrv4 I__6589 (
            .O(N__45933),
            .I(\c0.n3_adj_4636 ));
    Odrv4 I__6588 (
            .O(N__45926),
            .I(\c0.n3_adj_4636 ));
    CascadeMux I__6587 (
            .O(N__45915),
            .I(N__45912));
    InMux I__6586 (
            .O(N__45912),
            .I(N__45887));
    InMux I__6585 (
            .O(N__45911),
            .I(N__45887));
    InMux I__6584 (
            .O(N__45910),
            .I(N__45887));
    InMux I__6583 (
            .O(N__45909),
            .I(N__45874));
    InMux I__6582 (
            .O(N__45908),
            .I(N__45874));
    InMux I__6581 (
            .O(N__45907),
            .I(N__45874));
    InMux I__6580 (
            .O(N__45906),
            .I(N__45874));
    InMux I__6579 (
            .O(N__45905),
            .I(N__45874));
    InMux I__6578 (
            .O(N__45904),
            .I(N__45874));
    InMux I__6577 (
            .O(N__45903),
            .I(N__45869));
    InMux I__6576 (
            .O(N__45902),
            .I(N__45869));
    CascadeMux I__6575 (
            .O(N__45901),
            .I(N__45866));
    CascadeMux I__6574 (
            .O(N__45900),
            .I(N__45863));
    InMux I__6573 (
            .O(N__45899),
            .I(N__45853));
    InMux I__6572 (
            .O(N__45898),
            .I(N__45853));
    InMux I__6571 (
            .O(N__45897),
            .I(N__45853));
    InMux I__6570 (
            .O(N__45896),
            .I(N__45853));
    CascadeMux I__6569 (
            .O(N__45895),
            .I(N__45850));
    InMux I__6568 (
            .O(N__45894),
            .I(N__45847));
    LocalMux I__6567 (
            .O(N__45887),
            .I(N__45844));
    LocalMux I__6566 (
            .O(N__45874),
            .I(N__45841));
    LocalMux I__6565 (
            .O(N__45869),
            .I(N__45838));
    InMux I__6564 (
            .O(N__45866),
            .I(N__45826));
    InMux I__6563 (
            .O(N__45863),
            .I(N__45826));
    InMux I__6562 (
            .O(N__45862),
            .I(N__45826));
    LocalMux I__6561 (
            .O(N__45853),
            .I(N__45823));
    InMux I__6560 (
            .O(N__45850),
            .I(N__45820));
    LocalMux I__6559 (
            .O(N__45847),
            .I(N__45815));
    Span4Mux_v I__6558 (
            .O(N__45844),
            .I(N__45815));
    Span4Mux_h I__6557 (
            .O(N__45841),
            .I(N__45810));
    Span4Mux_h I__6556 (
            .O(N__45838),
            .I(N__45810));
    InMux I__6555 (
            .O(N__45837),
            .I(N__45806));
    InMux I__6554 (
            .O(N__45836),
            .I(N__45803));
    InMux I__6553 (
            .O(N__45835),
            .I(N__45796));
    InMux I__6552 (
            .O(N__45834),
            .I(N__45796));
    InMux I__6551 (
            .O(N__45833),
            .I(N__45796));
    LocalMux I__6550 (
            .O(N__45826),
            .I(N__45791));
    Span4Mux_v I__6549 (
            .O(N__45823),
            .I(N__45791));
    LocalMux I__6548 (
            .O(N__45820),
            .I(N__45786));
    Span4Mux_h I__6547 (
            .O(N__45815),
            .I(N__45786));
    Span4Mux_h I__6546 (
            .O(N__45810),
            .I(N__45783));
    InMux I__6545 (
            .O(N__45809),
            .I(N__45780));
    LocalMux I__6544 (
            .O(N__45806),
            .I(\c0.n45_adj_4637 ));
    LocalMux I__6543 (
            .O(N__45803),
            .I(\c0.n45_adj_4637 ));
    LocalMux I__6542 (
            .O(N__45796),
            .I(\c0.n45_adj_4637 ));
    Odrv4 I__6541 (
            .O(N__45791),
            .I(\c0.n45_adj_4637 ));
    Odrv4 I__6540 (
            .O(N__45786),
            .I(\c0.n45_adj_4637 ));
    Odrv4 I__6539 (
            .O(N__45783),
            .I(\c0.n45_adj_4637 ));
    LocalMux I__6538 (
            .O(N__45780),
            .I(\c0.n45_adj_4637 ));
    InMux I__6537 (
            .O(N__45765),
            .I(\quad_counter0.n30312 ));
    InMux I__6536 (
            .O(N__45762),
            .I(\quad_counter0.n30313 ));
    InMux I__6535 (
            .O(N__45759),
            .I(N__45754));
    InMux I__6534 (
            .O(N__45758),
            .I(N__45751));
    InMux I__6533 (
            .O(N__45757),
            .I(N__45748));
    LocalMux I__6532 (
            .O(N__45754),
            .I(N__45745));
    LocalMux I__6531 (
            .O(N__45751),
            .I(\quad_counter0.n2813 ));
    LocalMux I__6530 (
            .O(N__45748),
            .I(\quad_counter0.n2813 ));
    Odrv4 I__6529 (
            .O(N__45745),
            .I(\quad_counter0.n2813 ));
    InMux I__6528 (
            .O(N__45738),
            .I(N__45733));
    InMux I__6527 (
            .O(N__45737),
            .I(N__45730));
    InMux I__6526 (
            .O(N__45736),
            .I(N__45727));
    LocalMux I__6525 (
            .O(N__45733),
            .I(\quad_counter0.n2811 ));
    LocalMux I__6524 (
            .O(N__45730),
            .I(\quad_counter0.n2811 ));
    LocalMux I__6523 (
            .O(N__45727),
            .I(\quad_counter0.n2811 ));
    CascadeMux I__6522 (
            .O(N__45720),
            .I(N__45715));
    InMux I__6521 (
            .O(N__45719),
            .I(N__45712));
    InMux I__6520 (
            .O(N__45718),
            .I(N__45709));
    InMux I__6519 (
            .O(N__45715),
            .I(N__45706));
    LocalMux I__6518 (
            .O(N__45712),
            .I(\quad_counter0.n2810 ));
    LocalMux I__6517 (
            .O(N__45709),
            .I(\quad_counter0.n2810 ));
    LocalMux I__6516 (
            .O(N__45706),
            .I(\quad_counter0.n2810 ));
    InMux I__6515 (
            .O(N__45699),
            .I(N__45694));
    InMux I__6514 (
            .O(N__45698),
            .I(N__45691));
    InMux I__6513 (
            .O(N__45697),
            .I(N__45688));
    LocalMux I__6512 (
            .O(N__45694),
            .I(\quad_counter0.n2807 ));
    LocalMux I__6511 (
            .O(N__45691),
            .I(\quad_counter0.n2807 ));
    LocalMux I__6510 (
            .O(N__45688),
            .I(\quad_counter0.n2807 ));
    InMux I__6509 (
            .O(N__45681),
            .I(N__45676));
    InMux I__6508 (
            .O(N__45680),
            .I(N__45673));
    InMux I__6507 (
            .O(N__45679),
            .I(N__45670));
    LocalMux I__6506 (
            .O(N__45676),
            .I(\quad_counter0.n2808 ));
    LocalMux I__6505 (
            .O(N__45673),
            .I(\quad_counter0.n2808 ));
    LocalMux I__6504 (
            .O(N__45670),
            .I(\quad_counter0.n2808 ));
    InMux I__6503 (
            .O(N__45663),
            .I(N__45660));
    LocalMux I__6502 (
            .O(N__45660),
            .I(N__45655));
    InMux I__6501 (
            .O(N__45659),
            .I(N__45652));
    InMux I__6500 (
            .O(N__45658),
            .I(N__45649));
    Span4Mux_h I__6499 (
            .O(N__45655),
            .I(N__45646));
    LocalMux I__6498 (
            .O(N__45652),
            .I(N__45643));
    LocalMux I__6497 (
            .O(N__45649),
            .I(N__45640));
    Odrv4 I__6496 (
            .O(N__45646),
            .I(\quad_counter0.n2812 ));
    Odrv4 I__6495 (
            .O(N__45643),
            .I(\quad_counter0.n2812 ));
    Odrv4 I__6494 (
            .O(N__45640),
            .I(\quad_counter0.n2812 ));
    CascadeMux I__6493 (
            .O(N__45633),
            .I(N__45628));
    InMux I__6492 (
            .O(N__45632),
            .I(N__45625));
    InMux I__6491 (
            .O(N__45631),
            .I(N__45622));
    InMux I__6490 (
            .O(N__45628),
            .I(N__45619));
    LocalMux I__6489 (
            .O(N__45625),
            .I(\quad_counter0.n2805 ));
    LocalMux I__6488 (
            .O(N__45622),
            .I(\quad_counter0.n2805 ));
    LocalMux I__6487 (
            .O(N__45619),
            .I(\quad_counter0.n2805 ));
    InMux I__6486 (
            .O(N__45612),
            .I(N__45608));
    InMux I__6485 (
            .O(N__45611),
            .I(N__45605));
    LocalMux I__6484 (
            .O(N__45608),
            .I(N__45602));
    LocalMux I__6483 (
            .O(N__45605),
            .I(N__45596));
    Span4Mux_h I__6482 (
            .O(N__45602),
            .I(N__45596));
    InMux I__6481 (
            .O(N__45601),
            .I(N__45593));
    Odrv4 I__6480 (
            .O(N__45596),
            .I(\quad_counter0.n2804 ));
    LocalMux I__6479 (
            .O(N__45593),
            .I(\quad_counter0.n2804 ));
    InMux I__6478 (
            .O(N__45588),
            .I(N__45583));
    InMux I__6477 (
            .O(N__45587),
            .I(N__45580));
    InMux I__6476 (
            .O(N__45586),
            .I(N__45577));
    LocalMux I__6475 (
            .O(N__45583),
            .I(\quad_counter0.n2806 ));
    LocalMux I__6474 (
            .O(N__45580),
            .I(\quad_counter0.n2806 ));
    LocalMux I__6473 (
            .O(N__45577),
            .I(\quad_counter0.n2806 ));
    CascadeMux I__6472 (
            .O(N__45570),
            .I(\quad_counter0.n19_adj_4409_cascade_ ));
    InMux I__6471 (
            .O(N__45567),
            .I(N__45564));
    LocalMux I__6470 (
            .O(N__45564),
            .I(\quad_counter0.n18_adj_4408 ));
    CascadeMux I__6469 (
            .O(N__45561),
            .I(N__45549));
    CascadeMux I__6468 (
            .O(N__45560),
            .I(N__45546));
    CascadeMux I__6467 (
            .O(N__45559),
            .I(N__45542));
    CascadeMux I__6466 (
            .O(N__45558),
            .I(N__45539));
    CascadeMux I__6465 (
            .O(N__45557),
            .I(N__45536));
    CascadeMux I__6464 (
            .O(N__45556),
            .I(N__45533));
    CascadeMux I__6463 (
            .O(N__45555),
            .I(N__45530));
    CascadeMux I__6462 (
            .O(N__45554),
            .I(N__45527));
    CascadeMux I__6461 (
            .O(N__45553),
            .I(N__45524));
    CascadeMux I__6460 (
            .O(N__45552),
            .I(N__45521));
    InMux I__6459 (
            .O(N__45549),
            .I(N__45516));
    InMux I__6458 (
            .O(N__45546),
            .I(N__45516));
    CascadeMux I__6457 (
            .O(N__45545),
            .I(N__45513));
    InMux I__6456 (
            .O(N__45542),
            .I(N__45503));
    InMux I__6455 (
            .O(N__45539),
            .I(N__45503));
    InMux I__6454 (
            .O(N__45536),
            .I(N__45503));
    InMux I__6453 (
            .O(N__45533),
            .I(N__45503));
    InMux I__6452 (
            .O(N__45530),
            .I(N__45494));
    InMux I__6451 (
            .O(N__45527),
            .I(N__45494));
    InMux I__6450 (
            .O(N__45524),
            .I(N__45494));
    InMux I__6449 (
            .O(N__45521),
            .I(N__45494));
    LocalMux I__6448 (
            .O(N__45516),
            .I(N__45491));
    InMux I__6447 (
            .O(N__45513),
            .I(N__45486));
    InMux I__6446 (
            .O(N__45512),
            .I(N__45486));
    LocalMux I__6445 (
            .O(N__45503),
            .I(\quad_counter0.n2837 ));
    LocalMux I__6444 (
            .O(N__45494),
            .I(\quad_counter0.n2837 ));
    Odrv4 I__6443 (
            .O(N__45491),
            .I(\quad_counter0.n2837 ));
    LocalMux I__6442 (
            .O(N__45486),
            .I(\quad_counter0.n2837 ));
    CascadeMux I__6441 (
            .O(N__45477),
            .I(N__45474));
    InMux I__6440 (
            .O(N__45474),
            .I(N__45469));
    InMux I__6439 (
            .O(N__45473),
            .I(N__45466));
    InMux I__6438 (
            .O(N__45472),
            .I(N__45463));
    LocalMux I__6437 (
            .O(N__45469),
            .I(N__45460));
    LocalMux I__6436 (
            .O(N__45466),
            .I(\quad_counter0.n2819 ));
    LocalMux I__6435 (
            .O(N__45463),
            .I(\quad_counter0.n2819 ));
    Odrv4 I__6434 (
            .O(N__45460),
            .I(\quad_counter0.n2819 ));
    InMux I__6433 (
            .O(N__45453),
            .I(N__45448));
    InMux I__6432 (
            .O(N__45452),
            .I(N__45445));
    InMux I__6431 (
            .O(N__45451),
            .I(N__45442));
    LocalMux I__6430 (
            .O(N__45448),
            .I(N__45439));
    LocalMux I__6429 (
            .O(N__45445),
            .I(\quad_counter0.n2817 ));
    LocalMux I__6428 (
            .O(N__45442),
            .I(\quad_counter0.n2817 ));
    Odrv4 I__6427 (
            .O(N__45439),
            .I(\quad_counter0.n2817 ));
    InMux I__6426 (
            .O(N__45432),
            .I(N__45427));
    InMux I__6425 (
            .O(N__45431),
            .I(N__45424));
    InMux I__6424 (
            .O(N__45430),
            .I(N__45421));
    LocalMux I__6423 (
            .O(N__45427),
            .I(N__45418));
    LocalMux I__6422 (
            .O(N__45424),
            .I(\quad_counter0.n2818 ));
    LocalMux I__6421 (
            .O(N__45421),
            .I(\quad_counter0.n2818 ));
    Odrv4 I__6420 (
            .O(N__45418),
            .I(\quad_counter0.n2818 ));
    CascadeMux I__6419 (
            .O(N__45411),
            .I(\quad_counter0.n28323_cascade_ ));
    InMux I__6418 (
            .O(N__45408),
            .I(N__45403));
    InMux I__6417 (
            .O(N__45407),
            .I(N__45400));
    InMux I__6416 (
            .O(N__45406),
            .I(N__45397));
    LocalMux I__6415 (
            .O(N__45403),
            .I(N__45394));
    LocalMux I__6414 (
            .O(N__45400),
            .I(\quad_counter0.n2814 ));
    LocalMux I__6413 (
            .O(N__45397),
            .I(\quad_counter0.n2814 ));
    Odrv4 I__6412 (
            .O(N__45394),
            .I(\quad_counter0.n2814 ));
    InMux I__6411 (
            .O(N__45387),
            .I(N__45382));
    InMux I__6410 (
            .O(N__45386),
            .I(N__45379));
    InMux I__6409 (
            .O(N__45385),
            .I(N__45376));
    LocalMux I__6408 (
            .O(N__45382),
            .I(N__45373));
    LocalMux I__6407 (
            .O(N__45379),
            .I(\quad_counter0.n2816 ));
    LocalMux I__6406 (
            .O(N__45376),
            .I(\quad_counter0.n2816 ));
    Odrv4 I__6405 (
            .O(N__45373),
            .I(\quad_counter0.n2816 ));
    InMux I__6404 (
            .O(N__45366),
            .I(N__45361));
    InMux I__6403 (
            .O(N__45365),
            .I(N__45358));
    InMux I__6402 (
            .O(N__45364),
            .I(N__45355));
    LocalMux I__6401 (
            .O(N__45361),
            .I(N__45352));
    LocalMux I__6400 (
            .O(N__45358),
            .I(\quad_counter0.n2815 ));
    LocalMux I__6399 (
            .O(N__45355),
            .I(\quad_counter0.n2815 ));
    Odrv4 I__6398 (
            .O(N__45352),
            .I(\quad_counter0.n2815 ));
    CascadeMux I__6397 (
            .O(N__45345),
            .I(\quad_counter0.n10_adj_4406_cascade_ ));
    InMux I__6396 (
            .O(N__45342),
            .I(N__45337));
    InMux I__6395 (
            .O(N__45341),
            .I(N__45334));
    InMux I__6394 (
            .O(N__45340),
            .I(N__45331));
    LocalMux I__6393 (
            .O(N__45337),
            .I(\quad_counter0.n2809 ));
    LocalMux I__6392 (
            .O(N__45334),
            .I(\quad_counter0.n2809 ));
    LocalMux I__6391 (
            .O(N__45331),
            .I(\quad_counter0.n2809 ));
    InMux I__6390 (
            .O(N__45324),
            .I(N__45321));
    LocalMux I__6389 (
            .O(N__45321),
            .I(\quad_counter0.n12_adj_4407 ));
    InMux I__6388 (
            .O(N__45318),
            .I(\quad_counter0.n30303 ));
    InMux I__6387 (
            .O(N__45315),
            .I(\quad_counter0.n30304 ));
    InMux I__6386 (
            .O(N__45312),
            .I(\quad_counter0.n30305 ));
    InMux I__6385 (
            .O(N__45309),
            .I(bfn_12_14_0_));
    InMux I__6384 (
            .O(N__45306),
            .I(\quad_counter0.n30307 ));
    InMux I__6383 (
            .O(N__45303),
            .I(\quad_counter0.n30308 ));
    InMux I__6382 (
            .O(N__45300),
            .I(\quad_counter0.n30309 ));
    InMux I__6381 (
            .O(N__45297),
            .I(\quad_counter0.n30310 ));
    InMux I__6380 (
            .O(N__45294),
            .I(\quad_counter0.n30311 ));
    InMux I__6379 (
            .O(N__45291),
            .I(N__45287));
    InMux I__6378 (
            .O(N__45290),
            .I(N__45284));
    LocalMux I__6377 (
            .O(N__45287),
            .I(N__45278));
    LocalMux I__6376 (
            .O(N__45284),
            .I(N__45278));
    InMux I__6375 (
            .O(N__45283),
            .I(N__45275));
    Odrv4 I__6374 (
            .O(N__45278),
            .I(\quad_counter0.n3301 ));
    LocalMux I__6373 (
            .O(N__45275),
            .I(\quad_counter0.n3301 ));
    InMux I__6372 (
            .O(N__45270),
            .I(\quad_counter0.n30422 ));
    InMux I__6371 (
            .O(N__45267),
            .I(N__45263));
    InMux I__6370 (
            .O(N__45266),
            .I(N__45260));
    LocalMux I__6369 (
            .O(N__45263),
            .I(N__45254));
    LocalMux I__6368 (
            .O(N__45260),
            .I(N__45254));
    InMux I__6367 (
            .O(N__45259),
            .I(N__45251));
    Odrv4 I__6366 (
            .O(N__45254),
            .I(\quad_counter0.n3300 ));
    LocalMux I__6365 (
            .O(N__45251),
            .I(\quad_counter0.n3300 ));
    InMux I__6364 (
            .O(N__45246),
            .I(\quad_counter0.n30423 ));
    InMux I__6363 (
            .O(N__45243),
            .I(N__45239));
    InMux I__6362 (
            .O(N__45242),
            .I(N__45236));
    LocalMux I__6361 (
            .O(N__45239),
            .I(N__45230));
    LocalMux I__6360 (
            .O(N__45236),
            .I(N__45230));
    InMux I__6359 (
            .O(N__45235),
            .I(N__45227));
    Odrv4 I__6358 (
            .O(N__45230),
            .I(\quad_counter0.n3299 ));
    LocalMux I__6357 (
            .O(N__45227),
            .I(\quad_counter0.n3299 ));
    CascadeMux I__6356 (
            .O(N__45222),
            .I(N__45204));
    CascadeMux I__6355 (
            .O(N__45221),
            .I(N__45201));
    CascadeMux I__6354 (
            .O(N__45220),
            .I(N__45198));
    CascadeMux I__6353 (
            .O(N__45219),
            .I(N__45195));
    CascadeMux I__6352 (
            .O(N__45218),
            .I(N__45192));
    CascadeMux I__6351 (
            .O(N__45217),
            .I(N__45189));
    CascadeMux I__6350 (
            .O(N__45216),
            .I(N__45186));
    CascadeMux I__6349 (
            .O(N__45215),
            .I(N__45183));
    CascadeMux I__6348 (
            .O(N__45214),
            .I(N__45180));
    CascadeMux I__6347 (
            .O(N__45213),
            .I(N__45177));
    CascadeMux I__6346 (
            .O(N__45212),
            .I(N__45174));
    CascadeMux I__6345 (
            .O(N__45211),
            .I(N__45171));
    CascadeMux I__6344 (
            .O(N__45210),
            .I(N__45168));
    CascadeMux I__6343 (
            .O(N__45209),
            .I(N__45165));
    CascadeMux I__6342 (
            .O(N__45208),
            .I(N__45162));
    CascadeMux I__6341 (
            .O(N__45207),
            .I(N__45159));
    InMux I__6340 (
            .O(N__45204),
            .I(N__45152));
    InMux I__6339 (
            .O(N__45201),
            .I(N__45152));
    InMux I__6338 (
            .O(N__45198),
            .I(N__45152));
    InMux I__6337 (
            .O(N__45195),
            .I(N__45145));
    InMux I__6336 (
            .O(N__45192),
            .I(N__45145));
    InMux I__6335 (
            .O(N__45189),
            .I(N__45145));
    InMux I__6334 (
            .O(N__45186),
            .I(N__45136));
    InMux I__6333 (
            .O(N__45183),
            .I(N__45136));
    InMux I__6332 (
            .O(N__45180),
            .I(N__45136));
    InMux I__6331 (
            .O(N__45177),
            .I(N__45136));
    InMux I__6330 (
            .O(N__45174),
            .I(N__45127));
    InMux I__6329 (
            .O(N__45171),
            .I(N__45127));
    InMux I__6328 (
            .O(N__45168),
            .I(N__45127));
    InMux I__6327 (
            .O(N__45165),
            .I(N__45127));
    InMux I__6326 (
            .O(N__45162),
            .I(N__45122));
    InMux I__6325 (
            .O(N__45159),
            .I(N__45122));
    LocalMux I__6324 (
            .O(N__45152),
            .I(N__45116));
    LocalMux I__6323 (
            .O(N__45145),
            .I(N__45116));
    LocalMux I__6322 (
            .O(N__45136),
            .I(N__45111));
    LocalMux I__6321 (
            .O(N__45127),
            .I(N__45111));
    LocalMux I__6320 (
            .O(N__45122),
            .I(N__45108));
    InMux I__6319 (
            .O(N__45121),
            .I(N__45105));
    Span4Mux_v I__6318 (
            .O(N__45116),
            .I(N__45096));
    Span4Mux_h I__6317 (
            .O(N__45111),
            .I(N__45096));
    Span4Mux_v I__6316 (
            .O(N__45108),
            .I(N__45096));
    LocalMux I__6315 (
            .O(N__45105),
            .I(N__45096));
    Odrv4 I__6314 (
            .O(N__45096),
            .I(\quad_counter0.n3332 ));
    InMux I__6313 (
            .O(N__45093),
            .I(\quad_counter0.n30424 ));
    InMux I__6312 (
            .O(N__45090),
            .I(N__45087));
    LocalMux I__6311 (
            .O(N__45087),
            .I(N__45084));
    Span4Mux_h I__6310 (
            .O(N__45084),
            .I(N__45079));
    InMux I__6309 (
            .O(N__45083),
            .I(N__45076));
    InMux I__6308 (
            .O(N__45082),
            .I(N__45073));
    Span4Mux_h I__6307 (
            .O(N__45079),
            .I(N__45070));
    LocalMux I__6306 (
            .O(N__45076),
            .I(\c0.FRAME_MATCHER_state_5 ));
    LocalMux I__6305 (
            .O(N__45073),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv4 I__6304 (
            .O(N__45070),
            .I(\c0.FRAME_MATCHER_state_5 ));
    SRMux I__6303 (
            .O(N__45063),
            .I(N__45060));
    LocalMux I__6302 (
            .O(N__45060),
            .I(\c0.n32730 ));
    InMux I__6301 (
            .O(N__45057),
            .I(bfn_12_13_0_));
    InMux I__6300 (
            .O(N__45054),
            .I(\quad_counter0.n30299 ));
    InMux I__6299 (
            .O(N__45051),
            .I(\quad_counter0.n30300 ));
    InMux I__6298 (
            .O(N__45048),
            .I(\quad_counter0.n30301 ));
    InMux I__6297 (
            .O(N__45045),
            .I(\quad_counter0.n30302 ));
    InMux I__6296 (
            .O(N__45042),
            .I(N__45037));
    InMux I__6295 (
            .O(N__45041),
            .I(N__45034));
    CascadeMux I__6294 (
            .O(N__45040),
            .I(N__45031));
    LocalMux I__6293 (
            .O(N__45037),
            .I(N__45026));
    LocalMux I__6292 (
            .O(N__45034),
            .I(N__45026));
    InMux I__6291 (
            .O(N__45031),
            .I(N__45023));
    Odrv12 I__6290 (
            .O(N__45026),
            .I(\quad_counter0.n3309 ));
    LocalMux I__6289 (
            .O(N__45023),
            .I(\quad_counter0.n3309 ));
    InMux I__6288 (
            .O(N__45018),
            .I(\quad_counter0.n30414 ));
    InMux I__6287 (
            .O(N__45015),
            .I(N__45011));
    InMux I__6286 (
            .O(N__45014),
            .I(N__45008));
    LocalMux I__6285 (
            .O(N__45011),
            .I(N__45002));
    LocalMux I__6284 (
            .O(N__45008),
            .I(N__45002));
    InMux I__6283 (
            .O(N__45007),
            .I(N__44999));
    Odrv4 I__6282 (
            .O(N__45002),
            .I(\quad_counter0.n3308 ));
    LocalMux I__6281 (
            .O(N__44999),
            .I(\quad_counter0.n3308 ));
    InMux I__6280 (
            .O(N__44994),
            .I(\quad_counter0.n30415 ));
    InMux I__6279 (
            .O(N__44991),
            .I(N__44987));
    InMux I__6278 (
            .O(N__44990),
            .I(N__44984));
    LocalMux I__6277 (
            .O(N__44987),
            .I(N__44978));
    LocalMux I__6276 (
            .O(N__44984),
            .I(N__44978));
    InMux I__6275 (
            .O(N__44983),
            .I(N__44975));
    Odrv4 I__6274 (
            .O(N__44978),
            .I(\quad_counter0.n3307 ));
    LocalMux I__6273 (
            .O(N__44975),
            .I(\quad_counter0.n3307 ));
    InMux I__6272 (
            .O(N__44970),
            .I(\quad_counter0.n30416 ));
    InMux I__6271 (
            .O(N__44967),
            .I(N__44963));
    InMux I__6270 (
            .O(N__44966),
            .I(N__44960));
    LocalMux I__6269 (
            .O(N__44963),
            .I(N__44954));
    LocalMux I__6268 (
            .O(N__44960),
            .I(N__44954));
    InMux I__6267 (
            .O(N__44959),
            .I(N__44951));
    Odrv12 I__6266 (
            .O(N__44954),
            .I(\quad_counter0.n3306 ));
    LocalMux I__6265 (
            .O(N__44951),
            .I(\quad_counter0.n3306 ));
    InMux I__6264 (
            .O(N__44946),
            .I(\quad_counter0.n30417 ));
    InMux I__6263 (
            .O(N__44943),
            .I(N__44939));
    InMux I__6262 (
            .O(N__44942),
            .I(N__44936));
    LocalMux I__6261 (
            .O(N__44939),
            .I(N__44930));
    LocalMux I__6260 (
            .O(N__44936),
            .I(N__44930));
    InMux I__6259 (
            .O(N__44935),
            .I(N__44927));
    Odrv4 I__6258 (
            .O(N__44930),
            .I(\quad_counter0.n3305 ));
    LocalMux I__6257 (
            .O(N__44927),
            .I(\quad_counter0.n3305 ));
    InMux I__6256 (
            .O(N__44922),
            .I(\quad_counter0.n30418 ));
    InMux I__6255 (
            .O(N__44919),
            .I(N__44915));
    InMux I__6254 (
            .O(N__44918),
            .I(N__44912));
    LocalMux I__6253 (
            .O(N__44915),
            .I(N__44907));
    LocalMux I__6252 (
            .O(N__44912),
            .I(N__44907));
    Span4Mux_h I__6251 (
            .O(N__44907),
            .I(N__44903));
    InMux I__6250 (
            .O(N__44906),
            .I(N__44900));
    Odrv4 I__6249 (
            .O(N__44903),
            .I(\quad_counter0.n3304 ));
    LocalMux I__6248 (
            .O(N__44900),
            .I(\quad_counter0.n3304 ));
    InMux I__6247 (
            .O(N__44895),
            .I(bfn_12_11_0_));
    InMux I__6246 (
            .O(N__44892),
            .I(N__44888));
    InMux I__6245 (
            .O(N__44891),
            .I(N__44885));
    LocalMux I__6244 (
            .O(N__44888),
            .I(N__44879));
    LocalMux I__6243 (
            .O(N__44885),
            .I(N__44879));
    InMux I__6242 (
            .O(N__44884),
            .I(N__44876));
    Odrv12 I__6241 (
            .O(N__44879),
            .I(\quad_counter0.n3303 ));
    LocalMux I__6240 (
            .O(N__44876),
            .I(\quad_counter0.n3303 ));
    InMux I__6239 (
            .O(N__44871),
            .I(\quad_counter0.n30420 ));
    InMux I__6238 (
            .O(N__44868),
            .I(N__44863));
    InMux I__6237 (
            .O(N__44867),
            .I(N__44860));
    CascadeMux I__6236 (
            .O(N__44866),
            .I(N__44857));
    LocalMux I__6235 (
            .O(N__44863),
            .I(N__44852));
    LocalMux I__6234 (
            .O(N__44860),
            .I(N__44852));
    InMux I__6233 (
            .O(N__44857),
            .I(N__44849));
    Odrv4 I__6232 (
            .O(N__44852),
            .I(\quad_counter0.n3302 ));
    LocalMux I__6231 (
            .O(N__44849),
            .I(\quad_counter0.n3302 ));
    InMux I__6230 (
            .O(N__44844),
            .I(\quad_counter0.n30421 ));
    InMux I__6229 (
            .O(N__44841),
            .I(\quad_counter0.n30405 ));
    InMux I__6228 (
            .O(N__44838),
            .I(\quad_counter0.n30406 ));
    InMux I__6227 (
            .O(N__44835),
            .I(\quad_counter0.n30407 ));
    InMux I__6226 (
            .O(N__44832),
            .I(\quad_counter0.n30408 ));
    CascadeMux I__6225 (
            .O(N__44829),
            .I(N__44821));
    CascadeMux I__6224 (
            .O(N__44828),
            .I(N__44818));
    CascadeMux I__6223 (
            .O(N__44827),
            .I(N__44815));
    CascadeMux I__6222 (
            .O(N__44826),
            .I(N__44812));
    CascadeMux I__6221 (
            .O(N__44825),
            .I(N__44809));
    CascadeMux I__6220 (
            .O(N__44824),
            .I(N__44806));
    InMux I__6219 (
            .O(N__44821),
            .I(N__44801));
    InMux I__6218 (
            .O(N__44818),
            .I(N__44801));
    InMux I__6217 (
            .O(N__44815),
            .I(N__44792));
    InMux I__6216 (
            .O(N__44812),
            .I(N__44792));
    InMux I__6215 (
            .O(N__44809),
            .I(N__44792));
    InMux I__6214 (
            .O(N__44806),
            .I(N__44792));
    LocalMux I__6213 (
            .O(N__44801),
            .I(\quad_counter0.n36140 ));
    LocalMux I__6212 (
            .O(N__44792),
            .I(\quad_counter0.n36140 ));
    InMux I__6211 (
            .O(N__44787),
            .I(\quad_counter0.n30409 ));
    InMux I__6210 (
            .O(N__44784),
            .I(N__44780));
    InMux I__6209 (
            .O(N__44783),
            .I(N__44777));
    LocalMux I__6208 (
            .O(N__44780),
            .I(N__44771));
    LocalMux I__6207 (
            .O(N__44777),
            .I(N__44771));
    CascadeMux I__6206 (
            .O(N__44776),
            .I(N__44768));
    Span4Mux_h I__6205 (
            .O(N__44771),
            .I(N__44765));
    InMux I__6204 (
            .O(N__44768),
            .I(N__44762));
    Odrv4 I__6203 (
            .O(N__44765),
            .I(\quad_counter0.n3313 ));
    LocalMux I__6202 (
            .O(N__44762),
            .I(\quad_counter0.n3313 ));
    InMux I__6201 (
            .O(N__44757),
            .I(\quad_counter0.n30410 ));
    InMux I__6200 (
            .O(N__44754),
            .I(N__44750));
    InMux I__6199 (
            .O(N__44753),
            .I(N__44747));
    LocalMux I__6198 (
            .O(N__44750),
            .I(N__44742));
    LocalMux I__6197 (
            .O(N__44747),
            .I(N__44742));
    Span4Mux_h I__6196 (
            .O(N__44742),
            .I(N__44738));
    InMux I__6195 (
            .O(N__44741),
            .I(N__44735));
    Odrv4 I__6194 (
            .O(N__44738),
            .I(\quad_counter0.n3312 ));
    LocalMux I__6193 (
            .O(N__44735),
            .I(\quad_counter0.n3312 ));
    InMux I__6192 (
            .O(N__44730),
            .I(bfn_12_10_0_));
    InMux I__6191 (
            .O(N__44727),
            .I(N__44723));
    InMux I__6190 (
            .O(N__44726),
            .I(N__44720));
    LocalMux I__6189 (
            .O(N__44723),
            .I(N__44714));
    LocalMux I__6188 (
            .O(N__44720),
            .I(N__44714));
    InMux I__6187 (
            .O(N__44719),
            .I(N__44711));
    Odrv12 I__6186 (
            .O(N__44714),
            .I(\quad_counter0.n3311 ));
    LocalMux I__6185 (
            .O(N__44711),
            .I(\quad_counter0.n3311 ));
    InMux I__6184 (
            .O(N__44706),
            .I(\quad_counter0.n30412 ));
    InMux I__6183 (
            .O(N__44703),
            .I(N__44698));
    InMux I__6182 (
            .O(N__44702),
            .I(N__44695));
    CascadeMux I__6181 (
            .O(N__44701),
            .I(N__44692));
    LocalMux I__6180 (
            .O(N__44698),
            .I(N__44687));
    LocalMux I__6179 (
            .O(N__44695),
            .I(N__44687));
    InMux I__6178 (
            .O(N__44692),
            .I(N__44684));
    Odrv4 I__6177 (
            .O(N__44687),
            .I(\quad_counter0.n3310 ));
    LocalMux I__6176 (
            .O(N__44684),
            .I(\quad_counter0.n3310 ));
    InMux I__6175 (
            .O(N__44679),
            .I(\quad_counter0.n30413 ));
    CascadeMux I__6174 (
            .O(N__44676),
            .I(N__44673));
    InMux I__6173 (
            .O(N__44673),
            .I(N__44670));
    LocalMux I__6172 (
            .O(N__44670),
            .I(N__44667));
    Odrv4 I__6171 (
            .O(N__44667),
            .I(\quad_counter0.n1847 ));
    InMux I__6170 (
            .O(N__44664),
            .I(\quad_counter0.n30209 ));
    InMux I__6169 (
            .O(N__44661),
            .I(\quad_counter0.n30210 ));
    InMux I__6168 (
            .O(N__44658),
            .I(\quad_counter0.n30211 ));
    InMux I__6167 (
            .O(N__44655),
            .I(\quad_counter0.n30212 ));
    InMux I__6166 (
            .O(N__44652),
            .I(\quad_counter0.n30213 ));
    CascadeMux I__6165 (
            .O(N__44649),
            .I(N__44641));
    CascadeMux I__6164 (
            .O(N__44648),
            .I(N__44638));
    CascadeMux I__6163 (
            .O(N__44647),
            .I(N__44635));
    CascadeMux I__6162 (
            .O(N__44646),
            .I(N__44632));
    CascadeMux I__6161 (
            .O(N__44645),
            .I(N__44629));
    CascadeMux I__6160 (
            .O(N__44644),
            .I(N__44626));
    InMux I__6159 (
            .O(N__44641),
            .I(N__44621));
    InMux I__6158 (
            .O(N__44638),
            .I(N__44621));
    InMux I__6157 (
            .O(N__44635),
            .I(N__44612));
    InMux I__6156 (
            .O(N__44632),
            .I(N__44612));
    InMux I__6155 (
            .O(N__44629),
            .I(N__44612));
    InMux I__6154 (
            .O(N__44626),
            .I(N__44612));
    LocalMux I__6153 (
            .O(N__44621),
            .I(N__44607));
    LocalMux I__6152 (
            .O(N__44612),
            .I(N__44607));
    Odrv4 I__6151 (
            .O(N__44607),
            .I(\quad_counter0.n36158 ));
    InMux I__6150 (
            .O(N__44604),
            .I(\quad_counter0.n30214 ));
    InMux I__6149 (
            .O(N__44601),
            .I(N__44598));
    LocalMux I__6148 (
            .O(N__44598),
            .I(N__44593));
    InMux I__6147 (
            .O(N__44597),
            .I(N__44590));
    InMux I__6146 (
            .O(N__44596),
            .I(N__44586));
    Span4Mux_v I__6145 (
            .O(N__44593),
            .I(N__44581));
    LocalMux I__6144 (
            .O(N__44590),
            .I(N__44581));
    InMux I__6143 (
            .O(N__44589),
            .I(N__44578));
    LocalMux I__6142 (
            .O(N__44586),
            .I(N__44575));
    Span4Mux_v I__6141 (
            .O(N__44581),
            .I(N__44570));
    LocalMux I__6140 (
            .O(N__44578),
            .I(N__44570));
    Span4Mux_v I__6139 (
            .O(N__44575),
            .I(N__44567));
    Span4Mux_h I__6138 (
            .O(N__44570),
            .I(N__44564));
    Sp12to4 I__6137 (
            .O(N__44567),
            .I(N__44561));
    Span4Mux_h I__6136 (
            .O(N__44564),
            .I(N__44558));
    Span12Mux_h I__6135 (
            .O(N__44561),
            .I(N__44555));
    Span4Mux_v I__6134 (
            .O(N__44558),
            .I(N__44552));
    Odrv12 I__6133 (
            .O(N__44555),
            .I(PIN_12_c));
    Odrv4 I__6132 (
            .O(N__44552),
            .I(PIN_12_c));
    InMux I__6131 (
            .O(N__44547),
            .I(N__44544));
    LocalMux I__6130 (
            .O(N__44544),
            .I(N__44541));
    Odrv4 I__6129 (
            .O(N__44541),
            .I(n17985));
    CascadeMux I__6128 (
            .O(N__44538),
            .I(N__44535));
    InMux I__6127 (
            .O(N__44535),
            .I(N__44531));
    InMux I__6126 (
            .O(N__44534),
            .I(N__44528));
    LocalMux I__6125 (
            .O(N__44531),
            .I(N__44524));
    LocalMux I__6124 (
            .O(N__44528),
            .I(N__44521));
    InMux I__6123 (
            .O(N__44527),
            .I(N__44518));
    Odrv4 I__6122 (
            .O(N__44524),
            .I(quadA_delayed_adj_4812));
    Odrv4 I__6121 (
            .O(N__44521),
            .I(quadA_delayed_adj_4812));
    LocalMux I__6120 (
            .O(N__44518),
            .I(quadA_delayed_adj_4812));
    InMux I__6119 (
            .O(N__44511),
            .I(bfn_12_9_0_));
    InMux I__6118 (
            .O(N__44508),
            .I(\quad_counter0.n30404 ));
    InMux I__6117 (
            .O(N__44505),
            .I(N__44502));
    LocalMux I__6116 (
            .O(N__44502),
            .I(N__44499));
    Span4Mux_h I__6115 (
            .O(N__44499),
            .I(N__44493));
    InMux I__6114 (
            .O(N__44498),
            .I(N__44486));
    InMux I__6113 (
            .O(N__44497),
            .I(N__44486));
    InMux I__6112 (
            .O(N__44496),
            .I(N__44486));
    Odrv4 I__6111 (
            .O(N__44493),
            .I(\c0.data_in_frame_17_2 ));
    LocalMux I__6110 (
            .O(N__44486),
            .I(\c0.data_in_frame_17_2 ));
    InMux I__6109 (
            .O(N__44481),
            .I(N__44478));
    LocalMux I__6108 (
            .O(N__44478),
            .I(N__44472));
    InMux I__6107 (
            .O(N__44477),
            .I(N__44469));
    InMux I__6106 (
            .O(N__44476),
            .I(N__44464));
    InMux I__6105 (
            .O(N__44475),
            .I(N__44464));
    Odrv4 I__6104 (
            .O(N__44472),
            .I(\c0.data_in_frame_17_4 ));
    LocalMux I__6103 (
            .O(N__44469),
            .I(\c0.data_in_frame_17_4 ));
    LocalMux I__6102 (
            .O(N__44464),
            .I(\c0.data_in_frame_17_4 ));
    InMux I__6101 (
            .O(N__44457),
            .I(N__44453));
    InMux I__6100 (
            .O(N__44456),
            .I(N__44450));
    LocalMux I__6099 (
            .O(N__44453),
            .I(N__44445));
    LocalMux I__6098 (
            .O(N__44450),
            .I(N__44442));
    InMux I__6097 (
            .O(N__44449),
            .I(N__44439));
    InMux I__6096 (
            .O(N__44448),
            .I(N__44436));
    Span4Mux_h I__6095 (
            .O(N__44445),
            .I(N__44433));
    Span4Mux_v I__6094 (
            .O(N__44442),
            .I(N__44430));
    LocalMux I__6093 (
            .O(N__44439),
            .I(N__44427));
    LocalMux I__6092 (
            .O(N__44436),
            .I(\c0.data_in_frame_14_7 ));
    Odrv4 I__6091 (
            .O(N__44433),
            .I(\c0.data_in_frame_14_7 ));
    Odrv4 I__6090 (
            .O(N__44430),
            .I(\c0.data_in_frame_14_7 ));
    Odrv12 I__6089 (
            .O(N__44427),
            .I(\c0.data_in_frame_14_7 ));
    CascadeMux I__6088 (
            .O(N__44418),
            .I(\quad_counter0.n28397_cascade_ ));
    InMux I__6087 (
            .O(N__44415),
            .I(bfn_12_7_0_));
    InMux I__6086 (
            .O(N__44412),
            .I(N__44409));
    LocalMux I__6085 (
            .O(N__44409),
            .I(N__44406));
    Odrv4 I__6084 (
            .O(N__44406),
            .I(\c0.n33554 ));
    CascadeMux I__6083 (
            .O(N__44403),
            .I(\c0.n33824_cascade_ ));
    CascadeMux I__6082 (
            .O(N__44400),
            .I(\c0.n24_adj_4722_cascade_ ));
    CascadeMux I__6081 (
            .O(N__44397),
            .I(\c0.n26_adj_4724_cascade_ ));
    InMux I__6080 (
            .O(N__44394),
            .I(N__44391));
    LocalMux I__6079 (
            .O(N__44391),
            .I(N__44388));
    Odrv4 I__6078 (
            .O(N__44388),
            .I(\c0.n22_adj_4723 ));
    InMux I__6077 (
            .O(N__44385),
            .I(N__44382));
    LocalMux I__6076 (
            .O(N__44382),
            .I(\c0.n33 ));
    CascadeMux I__6075 (
            .O(N__44379),
            .I(N__44376));
    InMux I__6074 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__6073 (
            .O(N__44373),
            .I(N__44370));
    Odrv4 I__6072 (
            .O(N__44370),
            .I(\c0.n34_adj_4738 ));
    InMux I__6071 (
            .O(N__44367),
            .I(N__44364));
    LocalMux I__6070 (
            .O(N__44364),
            .I(N__44361));
    Odrv12 I__6069 (
            .O(N__44361),
            .I(\c0.n32_adj_4739 ));
    InMux I__6068 (
            .O(N__44358),
            .I(N__44354));
    InMux I__6067 (
            .O(N__44357),
            .I(N__44351));
    LocalMux I__6066 (
            .O(N__44354),
            .I(\c0.data_in_frame_15_0 ));
    LocalMux I__6065 (
            .O(N__44351),
            .I(\c0.data_in_frame_15_0 ));
    InMux I__6064 (
            .O(N__44346),
            .I(N__44339));
    InMux I__6063 (
            .O(N__44345),
            .I(N__44339));
    CascadeMux I__6062 (
            .O(N__44344),
            .I(N__44336));
    LocalMux I__6061 (
            .O(N__44339),
            .I(N__44332));
    InMux I__6060 (
            .O(N__44336),
            .I(N__44327));
    InMux I__6059 (
            .O(N__44335),
            .I(N__44327));
    Span4Mux_h I__6058 (
            .O(N__44332),
            .I(N__44324));
    LocalMux I__6057 (
            .O(N__44327),
            .I(\c0.data_in_frame_14_6 ));
    Odrv4 I__6056 (
            .O(N__44324),
            .I(\c0.data_in_frame_14_6 ));
    InMux I__6055 (
            .O(N__44319),
            .I(N__44315));
    InMux I__6054 (
            .O(N__44318),
            .I(N__44312));
    LocalMux I__6053 (
            .O(N__44315),
            .I(N__44308));
    LocalMux I__6052 (
            .O(N__44312),
            .I(N__44305));
    InMux I__6051 (
            .O(N__44311),
            .I(N__44302));
    Span4Mux_v I__6050 (
            .O(N__44308),
            .I(N__44299));
    Span4Mux_v I__6049 (
            .O(N__44305),
            .I(N__44296));
    LocalMux I__6048 (
            .O(N__44302),
            .I(N__44293));
    Odrv4 I__6047 (
            .O(N__44299),
            .I(\c0.n17582 ));
    Odrv4 I__6046 (
            .O(N__44296),
            .I(\c0.n17582 ));
    Odrv4 I__6045 (
            .O(N__44293),
            .I(\c0.n17582 ));
    CascadeMux I__6044 (
            .O(N__44286),
            .I(N__44283));
    InMux I__6043 (
            .O(N__44283),
            .I(N__44280));
    LocalMux I__6042 (
            .O(N__44280),
            .I(N__44277));
    Span4Mux_v I__6041 (
            .O(N__44277),
            .I(N__44274));
    Odrv4 I__6040 (
            .O(N__44274),
            .I(\c0.n18511 ));
    InMux I__6039 (
            .O(N__44271),
            .I(N__44264));
    InMux I__6038 (
            .O(N__44270),
            .I(N__44264));
    CascadeMux I__6037 (
            .O(N__44269),
            .I(N__44261));
    LocalMux I__6036 (
            .O(N__44264),
            .I(N__44257));
    InMux I__6035 (
            .O(N__44261),
            .I(N__44254));
    InMux I__6034 (
            .O(N__44260),
            .I(N__44251));
    Span4Mux_h I__6033 (
            .O(N__44257),
            .I(N__44248));
    LocalMux I__6032 (
            .O(N__44254),
            .I(N__44245));
    LocalMux I__6031 (
            .O(N__44251),
            .I(\c0.data_in_frame_8_7 ));
    Odrv4 I__6030 (
            .O(N__44248),
            .I(\c0.data_in_frame_8_7 ));
    Odrv12 I__6029 (
            .O(N__44245),
            .I(\c0.data_in_frame_8_7 ));
    CascadeMux I__6028 (
            .O(N__44238),
            .I(N__44234));
    InMux I__6027 (
            .O(N__44237),
            .I(N__44229));
    InMux I__6026 (
            .O(N__44234),
            .I(N__44229));
    LocalMux I__6025 (
            .O(N__44229),
            .I(N__44226));
    Odrv4 I__6024 (
            .O(N__44226),
            .I(\c0.n19102 ));
    InMux I__6023 (
            .O(N__44223),
            .I(N__44220));
    LocalMux I__6022 (
            .O(N__44220),
            .I(N__44217));
    Span4Mux_h I__6021 (
            .O(N__44217),
            .I(N__44214));
    Odrv4 I__6020 (
            .O(N__44214),
            .I(\c0.n33729 ));
    CascadeMux I__6019 (
            .O(N__44211),
            .I(\c0.n33729_cascade_ ));
    CascadeMux I__6018 (
            .O(N__44208),
            .I(N__44205));
    InMux I__6017 (
            .O(N__44205),
            .I(N__44202));
    LocalMux I__6016 (
            .O(N__44202),
            .I(\c0.n14_adj_4582 ));
    InMux I__6015 (
            .O(N__44199),
            .I(N__44196));
    LocalMux I__6014 (
            .O(N__44196),
            .I(N__44193));
    Span4Mux_v I__6013 (
            .O(N__44193),
            .I(N__44190));
    Odrv4 I__6012 (
            .O(N__44190),
            .I(\c0.n34000 ));
    InMux I__6011 (
            .O(N__44187),
            .I(N__44181));
    InMux I__6010 (
            .O(N__44186),
            .I(N__44181));
    LocalMux I__6009 (
            .O(N__44181),
            .I(N__44177));
    InMux I__6008 (
            .O(N__44180),
            .I(N__44174));
    Span4Mux_h I__6007 (
            .O(N__44177),
            .I(N__44170));
    LocalMux I__6006 (
            .O(N__44174),
            .I(N__44167));
    InMux I__6005 (
            .O(N__44173),
            .I(N__44164));
    Odrv4 I__6004 (
            .O(N__44170),
            .I(\c0.n19190 ));
    Odrv4 I__6003 (
            .O(N__44167),
            .I(\c0.n19190 ));
    LocalMux I__6002 (
            .O(N__44164),
            .I(\c0.n19190 ));
    InMux I__6001 (
            .O(N__44157),
            .I(N__44154));
    LocalMux I__6000 (
            .O(N__44154),
            .I(N__44150));
    InMux I__5999 (
            .O(N__44153),
            .I(N__44147));
    Odrv4 I__5998 (
            .O(N__44150),
            .I(\c0.n15998 ));
    LocalMux I__5997 (
            .O(N__44147),
            .I(\c0.n15998 ));
    InMux I__5996 (
            .O(N__44142),
            .I(N__44136));
    InMux I__5995 (
            .O(N__44141),
            .I(N__44131));
    InMux I__5994 (
            .O(N__44140),
            .I(N__44131));
    CascadeMux I__5993 (
            .O(N__44139),
            .I(N__44128));
    LocalMux I__5992 (
            .O(N__44136),
            .I(N__44123));
    LocalMux I__5991 (
            .O(N__44131),
            .I(N__44123));
    InMux I__5990 (
            .O(N__44128),
            .I(N__44120));
    Span4Mux_h I__5989 (
            .O(N__44123),
            .I(N__44117));
    LocalMux I__5988 (
            .O(N__44120),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__5987 (
            .O(N__44117),
            .I(\c0.data_in_frame_7_2 ));
    InMux I__5986 (
            .O(N__44112),
            .I(N__44107));
    InMux I__5985 (
            .O(N__44111),
            .I(N__44103));
    CascadeMux I__5984 (
            .O(N__44110),
            .I(N__44100));
    LocalMux I__5983 (
            .O(N__44107),
            .I(N__44097));
    InMux I__5982 (
            .O(N__44106),
            .I(N__44094));
    LocalMux I__5981 (
            .O(N__44103),
            .I(N__44091));
    InMux I__5980 (
            .O(N__44100),
            .I(N__44088));
    Span4Mux_h I__5979 (
            .O(N__44097),
            .I(N__44085));
    LocalMux I__5978 (
            .O(N__44094),
            .I(N__44082));
    Span4Mux_h I__5977 (
            .O(N__44091),
            .I(N__44079));
    LocalMux I__5976 (
            .O(N__44088),
            .I(\c0.data_in_frame_15_4 ));
    Odrv4 I__5975 (
            .O(N__44085),
            .I(\c0.data_in_frame_15_4 ));
    Odrv12 I__5974 (
            .O(N__44082),
            .I(\c0.data_in_frame_15_4 ));
    Odrv4 I__5973 (
            .O(N__44079),
            .I(\c0.data_in_frame_15_4 ));
    CascadeMux I__5972 (
            .O(N__44070),
            .I(\c0.n33908_cascade_ ));
    InMux I__5971 (
            .O(N__44067),
            .I(N__44064));
    LocalMux I__5970 (
            .O(N__44064),
            .I(\c0.n30_adj_4737 ));
    InMux I__5969 (
            .O(N__44061),
            .I(N__44057));
    InMux I__5968 (
            .O(N__44060),
            .I(N__44054));
    LocalMux I__5967 (
            .O(N__44057),
            .I(\c0.n18544 ));
    LocalMux I__5966 (
            .O(N__44054),
            .I(\c0.n18544 ));
    InMux I__5965 (
            .O(N__44049),
            .I(N__44040));
    InMux I__5964 (
            .O(N__44048),
            .I(N__44040));
    InMux I__5963 (
            .O(N__44047),
            .I(N__44040));
    LocalMux I__5962 (
            .O(N__44040),
            .I(\c0.data_in_frame_7_5 ));
    InMux I__5961 (
            .O(N__44037),
            .I(N__44033));
    InMux I__5960 (
            .O(N__44036),
            .I(N__44030));
    LocalMux I__5959 (
            .O(N__44033),
            .I(N__44027));
    LocalMux I__5958 (
            .O(N__44030),
            .I(N__44024));
    Odrv4 I__5957 (
            .O(N__44027),
            .I(\c0.n33954 ));
    Odrv4 I__5956 (
            .O(N__44024),
            .I(\c0.n33954 ));
    CascadeMux I__5955 (
            .O(N__44019),
            .I(\c0.n34003_cascade_ ));
    InMux I__5954 (
            .O(N__44016),
            .I(N__44012));
    InMux I__5953 (
            .O(N__44015),
            .I(N__44008));
    LocalMux I__5952 (
            .O(N__44012),
            .I(N__44005));
    InMux I__5951 (
            .O(N__44011),
            .I(N__44002));
    LocalMux I__5950 (
            .O(N__44008),
            .I(N__43999));
    Span4Mux_h I__5949 (
            .O(N__44005),
            .I(N__43992));
    LocalMux I__5948 (
            .O(N__44002),
            .I(N__43992));
    Span4Mux_v I__5947 (
            .O(N__43999),
            .I(N__43992));
    Odrv4 I__5946 (
            .O(N__43992),
            .I(\c0.n33758 ));
    CascadeMux I__5945 (
            .O(N__43989),
            .I(N__43984));
    InMux I__5944 (
            .O(N__43988),
            .I(N__43981));
    InMux I__5943 (
            .O(N__43987),
            .I(N__43976));
    InMux I__5942 (
            .O(N__43984),
            .I(N__43976));
    LocalMux I__5941 (
            .O(N__43981),
            .I(\c0.data_in_frame_15_5 ));
    LocalMux I__5940 (
            .O(N__43976),
            .I(\c0.data_in_frame_15_5 ));
    CascadeMux I__5939 (
            .O(N__43971),
            .I(N__43966));
    InMux I__5938 (
            .O(N__43970),
            .I(N__43961));
    InMux I__5937 (
            .O(N__43969),
            .I(N__43961));
    InMux I__5936 (
            .O(N__43966),
            .I(N__43958));
    LocalMux I__5935 (
            .O(N__43961),
            .I(N__43953));
    LocalMux I__5934 (
            .O(N__43958),
            .I(N__43953));
    Span4Mux_v I__5933 (
            .O(N__43953),
            .I(N__43950));
    Span4Mux_h I__5932 (
            .O(N__43950),
            .I(N__43947));
    Odrv4 I__5931 (
            .O(N__43947),
            .I(\c0.n33781 ));
    CascadeMux I__5930 (
            .O(N__43944),
            .I(\c0.n18847_cascade_ ));
    InMux I__5929 (
            .O(N__43941),
            .I(N__43938));
    LocalMux I__5928 (
            .O(N__43938),
            .I(\c0.n10_adj_4708 ));
    CascadeMux I__5927 (
            .O(N__43935),
            .I(N__43931));
    CascadeMux I__5926 (
            .O(N__43934),
            .I(N__43927));
    InMux I__5925 (
            .O(N__43931),
            .I(N__43924));
    InMux I__5924 (
            .O(N__43930),
            .I(N__43921));
    InMux I__5923 (
            .O(N__43927),
            .I(N__43918));
    LocalMux I__5922 (
            .O(N__43924),
            .I(N__43915));
    LocalMux I__5921 (
            .O(N__43921),
            .I(N__43912));
    LocalMux I__5920 (
            .O(N__43918),
            .I(N__43905));
    Span4Mux_h I__5919 (
            .O(N__43915),
            .I(N__43905));
    Span4Mux_v I__5918 (
            .O(N__43912),
            .I(N__43905));
    Odrv4 I__5917 (
            .O(N__43905),
            .I(\c0.data_in_frame_11_5 ));
    InMux I__5916 (
            .O(N__43902),
            .I(N__43898));
    InMux I__5915 (
            .O(N__43901),
            .I(N__43895));
    LocalMux I__5914 (
            .O(N__43898),
            .I(N__43892));
    LocalMux I__5913 (
            .O(N__43895),
            .I(\c0.data_out_frame_0__7__N_2744 ));
    Odrv4 I__5912 (
            .O(N__43892),
            .I(\c0.data_out_frame_0__7__N_2744 ));
    InMux I__5911 (
            .O(N__43887),
            .I(N__43884));
    LocalMux I__5910 (
            .O(N__43884),
            .I(\c0.n33650 ));
    InMux I__5909 (
            .O(N__43881),
            .I(N__43878));
    LocalMux I__5908 (
            .O(N__43878),
            .I(N__43873));
    InMux I__5907 (
            .O(N__43877),
            .I(N__43868));
    InMux I__5906 (
            .O(N__43876),
            .I(N__43868));
    Odrv4 I__5905 (
            .O(N__43873),
            .I(\c0.n32325 ));
    LocalMux I__5904 (
            .O(N__43868),
            .I(\c0.n32325 ));
    InMux I__5903 (
            .O(N__43863),
            .I(N__43860));
    LocalMux I__5902 (
            .O(N__43860),
            .I(N__43857));
    Odrv4 I__5901 (
            .O(N__43857),
            .I(\c0.n33311 ));
    CascadeMux I__5900 (
            .O(N__43854),
            .I(\c0.n33311_cascade_ ));
    CascadeMux I__5899 (
            .O(N__43851),
            .I(N__43848));
    InMux I__5898 (
            .O(N__43848),
            .I(N__43838));
    InMux I__5897 (
            .O(N__43847),
            .I(N__43838));
    InMux I__5896 (
            .O(N__43846),
            .I(N__43838));
    InMux I__5895 (
            .O(N__43845),
            .I(N__43833));
    LocalMux I__5894 (
            .O(N__43838),
            .I(N__43827));
    InMux I__5893 (
            .O(N__43837),
            .I(N__43822));
    InMux I__5892 (
            .O(N__43836),
            .I(N__43822));
    LocalMux I__5891 (
            .O(N__43833),
            .I(N__43819));
    InMux I__5890 (
            .O(N__43832),
            .I(N__43814));
    InMux I__5889 (
            .O(N__43831),
            .I(N__43814));
    CascadeMux I__5888 (
            .O(N__43830),
            .I(N__43811));
    Span4Mux_v I__5887 (
            .O(N__43827),
            .I(N__43806));
    LocalMux I__5886 (
            .O(N__43822),
            .I(N__43806));
    Span4Mux_v I__5885 (
            .O(N__43819),
            .I(N__43803));
    LocalMux I__5884 (
            .O(N__43814),
            .I(N__43800));
    InMux I__5883 (
            .O(N__43811),
            .I(N__43797));
    Span4Mux_h I__5882 (
            .O(N__43806),
            .I(N__43792));
    Span4Mux_h I__5881 (
            .O(N__43803),
            .I(N__43792));
    Span4Mux_h I__5880 (
            .O(N__43800),
            .I(N__43789));
    LocalMux I__5879 (
            .O(N__43797),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__5878 (
            .O(N__43792),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__5877 (
            .O(N__43789),
            .I(\c0.data_in_frame_0_4 ));
    InMux I__5876 (
            .O(N__43782),
            .I(N__43779));
    LocalMux I__5875 (
            .O(N__43779),
            .I(N__43773));
    InMux I__5874 (
            .O(N__43778),
            .I(N__43766));
    InMux I__5873 (
            .O(N__43777),
            .I(N__43766));
    InMux I__5872 (
            .O(N__43776),
            .I(N__43766));
    Odrv4 I__5871 (
            .O(N__43773),
            .I(\c0.data_in_frame_11_7 ));
    LocalMux I__5870 (
            .O(N__43766),
            .I(\c0.data_in_frame_11_7 ));
    InMux I__5869 (
            .O(N__43761),
            .I(N__43758));
    LocalMux I__5868 (
            .O(N__43758),
            .I(N__43754));
    InMux I__5867 (
            .O(N__43757),
            .I(N__43751));
    Odrv4 I__5866 (
            .O(N__43754),
            .I(\c0.n33523 ));
    LocalMux I__5865 (
            .O(N__43751),
            .I(\c0.n33523 ));
    InMux I__5864 (
            .O(N__43746),
            .I(N__43743));
    LocalMux I__5863 (
            .O(N__43743),
            .I(\c0.n14_adj_4771 ));
    InMux I__5862 (
            .O(N__43740),
            .I(N__43737));
    LocalMux I__5861 (
            .O(N__43737),
            .I(\c0.n13_adj_4773 ));
    CascadeMux I__5860 (
            .O(N__43734),
            .I(\c0.n14_adj_4772_cascade_ ));
    InMux I__5859 (
            .O(N__43731),
            .I(N__43728));
    LocalMux I__5858 (
            .O(N__43728),
            .I(\c0.n13_adj_4774 ));
    InMux I__5857 (
            .O(N__43725),
            .I(N__43722));
    LocalMux I__5856 (
            .O(N__43722),
            .I(N__43716));
    CascadeMux I__5855 (
            .O(N__43721),
            .I(N__43713));
    CascadeMux I__5854 (
            .O(N__43720),
            .I(N__43709));
    InMux I__5853 (
            .O(N__43719),
            .I(N__43706));
    Span4Mux_h I__5852 (
            .O(N__43716),
            .I(N__43703));
    InMux I__5851 (
            .O(N__43713),
            .I(N__43696));
    InMux I__5850 (
            .O(N__43712),
            .I(N__43696));
    InMux I__5849 (
            .O(N__43709),
            .I(N__43696));
    LocalMux I__5848 (
            .O(N__43706),
            .I(\c0.data_in_frame_8_5 ));
    Odrv4 I__5847 (
            .O(N__43703),
            .I(\c0.data_in_frame_8_5 ));
    LocalMux I__5846 (
            .O(N__43696),
            .I(\c0.data_in_frame_8_5 ));
    InMux I__5845 (
            .O(N__43689),
            .I(N__43686));
    LocalMux I__5844 (
            .O(N__43686),
            .I(N__43683));
    Odrv4 I__5843 (
            .O(N__43683),
            .I(\c0.n49 ));
    CascadeMux I__5842 (
            .O(N__43680),
            .I(N__43677));
    InMux I__5841 (
            .O(N__43677),
            .I(N__43668));
    InMux I__5840 (
            .O(N__43676),
            .I(N__43668));
    InMux I__5839 (
            .O(N__43675),
            .I(N__43668));
    LocalMux I__5838 (
            .O(N__43668),
            .I(\c0.data_in_frame_11_1 ));
    InMux I__5837 (
            .O(N__43665),
            .I(N__43661));
    InMux I__5836 (
            .O(N__43664),
            .I(N__43658));
    LocalMux I__5835 (
            .O(N__43661),
            .I(N__43653));
    LocalMux I__5834 (
            .O(N__43658),
            .I(N__43653));
    Odrv4 I__5833 (
            .O(N__43653),
            .I(\c0.n33476 ));
    CascadeMux I__5832 (
            .O(N__43650),
            .I(\c0.n19102_cascade_ ));
    InMux I__5831 (
            .O(N__43647),
            .I(N__43642));
    InMux I__5830 (
            .O(N__43646),
            .I(N__43639));
    InMux I__5829 (
            .O(N__43645),
            .I(N__43636));
    LocalMux I__5828 (
            .O(N__43642),
            .I(N__43633));
    LocalMux I__5827 (
            .O(N__43639),
            .I(\quad_counter0.n2909 ));
    LocalMux I__5826 (
            .O(N__43636),
            .I(\quad_counter0.n2909 ));
    Odrv4 I__5825 (
            .O(N__43633),
            .I(\quad_counter0.n2909 ));
    InMux I__5824 (
            .O(N__43626),
            .I(N__43621));
    InMux I__5823 (
            .O(N__43625),
            .I(N__43618));
    InMux I__5822 (
            .O(N__43624),
            .I(N__43615));
    LocalMux I__5821 (
            .O(N__43621),
            .I(N__43612));
    LocalMux I__5820 (
            .O(N__43618),
            .I(\quad_counter0.n2911 ));
    LocalMux I__5819 (
            .O(N__43615),
            .I(\quad_counter0.n2911 ));
    Odrv4 I__5818 (
            .O(N__43612),
            .I(\quad_counter0.n2911 ));
    CascadeMux I__5817 (
            .O(N__43605),
            .I(\quad_counter0.n22_cascade_ ));
    InMux I__5816 (
            .O(N__43602),
            .I(N__43599));
    LocalMux I__5815 (
            .O(N__43599),
            .I(\quad_counter0.n18 ));
    CascadeMux I__5814 (
            .O(N__43596),
            .I(N__43582));
    CascadeMux I__5813 (
            .O(N__43595),
            .I(N__43579));
    CascadeMux I__5812 (
            .O(N__43594),
            .I(N__43576));
    CascadeMux I__5811 (
            .O(N__43593),
            .I(N__43573));
    CascadeMux I__5810 (
            .O(N__43592),
            .I(N__43570));
    CascadeMux I__5809 (
            .O(N__43591),
            .I(N__43567));
    CascadeMux I__5808 (
            .O(N__43590),
            .I(N__43564));
    CascadeMux I__5807 (
            .O(N__43589),
            .I(N__43561));
    CascadeMux I__5806 (
            .O(N__43588),
            .I(N__43558));
    CascadeMux I__5805 (
            .O(N__43587),
            .I(N__43555));
    CascadeMux I__5804 (
            .O(N__43586),
            .I(N__43552));
    CascadeMux I__5803 (
            .O(N__43585),
            .I(N__43549));
    InMux I__5802 (
            .O(N__43582),
            .I(N__43544));
    InMux I__5801 (
            .O(N__43579),
            .I(N__43544));
    InMux I__5800 (
            .O(N__43576),
            .I(N__43540));
    InMux I__5799 (
            .O(N__43573),
            .I(N__43537));
    InMux I__5798 (
            .O(N__43570),
            .I(N__43528));
    InMux I__5797 (
            .O(N__43567),
            .I(N__43528));
    InMux I__5796 (
            .O(N__43564),
            .I(N__43528));
    InMux I__5795 (
            .O(N__43561),
            .I(N__43528));
    InMux I__5794 (
            .O(N__43558),
            .I(N__43519));
    InMux I__5793 (
            .O(N__43555),
            .I(N__43519));
    InMux I__5792 (
            .O(N__43552),
            .I(N__43519));
    InMux I__5791 (
            .O(N__43549),
            .I(N__43519));
    LocalMux I__5790 (
            .O(N__43544),
            .I(N__43516));
    InMux I__5789 (
            .O(N__43543),
            .I(N__43513));
    LocalMux I__5788 (
            .O(N__43540),
            .I(\quad_counter0.n2936 ));
    LocalMux I__5787 (
            .O(N__43537),
            .I(\quad_counter0.n2936 ));
    LocalMux I__5786 (
            .O(N__43528),
            .I(\quad_counter0.n2936 ));
    LocalMux I__5785 (
            .O(N__43519),
            .I(\quad_counter0.n2936 ));
    Odrv4 I__5784 (
            .O(N__43516),
            .I(\quad_counter0.n2936 ));
    LocalMux I__5783 (
            .O(N__43513),
            .I(\quad_counter0.n2936 ));
    InMux I__5782 (
            .O(N__43500),
            .I(N__43495));
    InMux I__5781 (
            .O(N__43499),
            .I(N__43492));
    InMux I__5780 (
            .O(N__43498),
            .I(N__43489));
    LocalMux I__5779 (
            .O(N__43495),
            .I(N__43486));
    LocalMux I__5778 (
            .O(N__43492),
            .I(\quad_counter0.n2917 ));
    LocalMux I__5777 (
            .O(N__43489),
            .I(\quad_counter0.n2917 ));
    Odrv4 I__5776 (
            .O(N__43486),
            .I(\quad_counter0.n2917 ));
    InMux I__5775 (
            .O(N__43479),
            .I(N__43474));
    InMux I__5774 (
            .O(N__43478),
            .I(N__43471));
    InMux I__5773 (
            .O(N__43477),
            .I(N__43468));
    LocalMux I__5772 (
            .O(N__43474),
            .I(N__43465));
    LocalMux I__5771 (
            .O(N__43471),
            .I(\quad_counter0.n2918 ));
    LocalMux I__5770 (
            .O(N__43468),
            .I(\quad_counter0.n2918 ));
    Odrv12 I__5769 (
            .O(N__43465),
            .I(\quad_counter0.n2918 ));
    CascadeMux I__5768 (
            .O(N__43458),
            .I(N__43455));
    InMux I__5767 (
            .O(N__43455),
            .I(N__43450));
    InMux I__5766 (
            .O(N__43454),
            .I(N__43447));
    InMux I__5765 (
            .O(N__43453),
            .I(N__43444));
    LocalMux I__5764 (
            .O(N__43450),
            .I(N__43441));
    LocalMux I__5763 (
            .O(N__43447),
            .I(\quad_counter0.n2914 ));
    LocalMux I__5762 (
            .O(N__43444),
            .I(\quad_counter0.n2914 ));
    Odrv4 I__5761 (
            .O(N__43441),
            .I(\quad_counter0.n2914 ));
    InMux I__5760 (
            .O(N__43434),
            .I(N__43431));
    LocalMux I__5759 (
            .O(N__43431),
            .I(\quad_counter0.n28315 ));
    InMux I__5758 (
            .O(N__43428),
            .I(N__43423));
    InMux I__5757 (
            .O(N__43427),
            .I(N__43420));
    InMux I__5756 (
            .O(N__43426),
            .I(N__43417));
    LocalMux I__5755 (
            .O(N__43423),
            .I(N__43414));
    LocalMux I__5754 (
            .O(N__43420),
            .I(\quad_counter0.n2916 ));
    LocalMux I__5753 (
            .O(N__43417),
            .I(\quad_counter0.n2916 ));
    Odrv4 I__5752 (
            .O(N__43414),
            .I(\quad_counter0.n2916 ));
    InMux I__5751 (
            .O(N__43407),
            .I(N__43402));
    InMux I__5750 (
            .O(N__43406),
            .I(N__43399));
    InMux I__5749 (
            .O(N__43405),
            .I(N__43396));
    LocalMux I__5748 (
            .O(N__43402),
            .I(N__43393));
    LocalMux I__5747 (
            .O(N__43399),
            .I(\quad_counter0.n2915 ));
    LocalMux I__5746 (
            .O(N__43396),
            .I(\quad_counter0.n2915 ));
    Odrv4 I__5745 (
            .O(N__43393),
            .I(\quad_counter0.n2915 ));
    CascadeMux I__5744 (
            .O(N__43386),
            .I(\quad_counter0.n10_adj_4348_cascade_ ));
    InMux I__5743 (
            .O(N__43383),
            .I(N__43378));
    InMux I__5742 (
            .O(N__43382),
            .I(N__43375));
    InMux I__5741 (
            .O(N__43381),
            .I(N__43372));
    LocalMux I__5740 (
            .O(N__43378),
            .I(N__43369));
    LocalMux I__5739 (
            .O(N__43375),
            .I(\quad_counter0.n2906 ));
    LocalMux I__5738 (
            .O(N__43372),
            .I(\quad_counter0.n2906 ));
    Odrv4 I__5737 (
            .O(N__43369),
            .I(\quad_counter0.n2906 ));
    InMux I__5736 (
            .O(N__43362),
            .I(N__43359));
    LocalMux I__5735 (
            .O(N__43359),
            .I(\quad_counter0.n13 ));
    InMux I__5734 (
            .O(N__43356),
            .I(N__43353));
    LocalMux I__5733 (
            .O(N__43353),
            .I(N__43347));
    InMux I__5732 (
            .O(N__43352),
            .I(N__43344));
    InMux I__5731 (
            .O(N__43351),
            .I(N__43339));
    InMux I__5730 (
            .O(N__43350),
            .I(N__43339));
    Span4Mux_v I__5729 (
            .O(N__43347),
            .I(N__43334));
    LocalMux I__5728 (
            .O(N__43344),
            .I(N__43334));
    LocalMux I__5727 (
            .O(N__43339),
            .I(\c0.n33454 ));
    Odrv4 I__5726 (
            .O(N__43334),
            .I(\c0.n33454 ));
    InMux I__5725 (
            .O(N__43329),
            .I(N__43326));
    LocalMux I__5724 (
            .O(N__43326),
            .I(N__43323));
    Odrv4 I__5723 (
            .O(N__43323),
            .I(\c0.n33720 ));
    InMux I__5722 (
            .O(N__43320),
            .I(N__43317));
    LocalMux I__5721 (
            .O(N__43317),
            .I(N__43312));
    InMux I__5720 (
            .O(N__43316),
            .I(N__43309));
    InMux I__5719 (
            .O(N__43315),
            .I(N__43306));
    Span4Mux_h I__5718 (
            .O(N__43312),
            .I(N__43303));
    LocalMux I__5717 (
            .O(N__43309),
            .I(N__43298));
    LocalMux I__5716 (
            .O(N__43306),
            .I(N__43298));
    Odrv4 I__5715 (
            .O(N__43303),
            .I(\c0.n33341 ));
    Odrv12 I__5714 (
            .O(N__43298),
            .I(\c0.n33341 ));
    InMux I__5713 (
            .O(N__43293),
            .I(\quad_counter0.n30327 ));
    InMux I__5712 (
            .O(N__43290),
            .I(\quad_counter0.n30328 ));
    InMux I__5711 (
            .O(N__43287),
            .I(bfn_11_16_0_));
    CascadeMux I__5710 (
            .O(N__43284),
            .I(N__43276));
    CascadeMux I__5709 (
            .O(N__43283),
            .I(N__43273));
    CascadeMux I__5708 (
            .O(N__43282),
            .I(N__43270));
    CascadeMux I__5707 (
            .O(N__43281),
            .I(N__43267));
    CascadeMux I__5706 (
            .O(N__43280),
            .I(N__43264));
    CascadeMux I__5705 (
            .O(N__43279),
            .I(N__43261));
    InMux I__5704 (
            .O(N__43276),
            .I(N__43256));
    InMux I__5703 (
            .O(N__43273),
            .I(N__43256));
    InMux I__5702 (
            .O(N__43270),
            .I(N__43247));
    InMux I__5701 (
            .O(N__43267),
            .I(N__43247));
    InMux I__5700 (
            .O(N__43264),
            .I(N__43247));
    InMux I__5699 (
            .O(N__43261),
            .I(N__43247));
    LocalMux I__5698 (
            .O(N__43256),
            .I(N__43242));
    LocalMux I__5697 (
            .O(N__43247),
            .I(N__43242));
    Odrv4 I__5696 (
            .O(N__43242),
            .I(\quad_counter0.n36147 ));
    CascadeMux I__5695 (
            .O(N__43239),
            .I(N__43234));
    InMux I__5694 (
            .O(N__43238),
            .I(N__43231));
    InMux I__5693 (
            .O(N__43237),
            .I(N__43228));
    InMux I__5692 (
            .O(N__43234),
            .I(N__43225));
    LocalMux I__5691 (
            .O(N__43231),
            .I(\quad_counter0.n2908 ));
    LocalMux I__5690 (
            .O(N__43228),
            .I(\quad_counter0.n2908 ));
    LocalMux I__5689 (
            .O(N__43225),
            .I(\quad_counter0.n2908 ));
    InMux I__5688 (
            .O(N__43218),
            .I(N__43215));
    LocalMux I__5687 (
            .O(N__43215),
            .I(N__43211));
    InMux I__5686 (
            .O(N__43214),
            .I(N__43208));
    Span4Mux_h I__5685 (
            .O(N__43211),
            .I(N__43204));
    LocalMux I__5684 (
            .O(N__43208),
            .I(N__43201));
    InMux I__5683 (
            .O(N__43207),
            .I(N__43198));
    Odrv4 I__5682 (
            .O(N__43204),
            .I(\quad_counter0.n2904 ));
    Odrv4 I__5681 (
            .O(N__43201),
            .I(\quad_counter0.n2904 ));
    LocalMux I__5680 (
            .O(N__43198),
            .I(\quad_counter0.n2904 ));
    InMux I__5679 (
            .O(N__43191),
            .I(N__43186));
    InMux I__5678 (
            .O(N__43190),
            .I(N__43183));
    InMux I__5677 (
            .O(N__43189),
            .I(N__43180));
    LocalMux I__5676 (
            .O(N__43186),
            .I(\quad_counter0.n2910 ));
    LocalMux I__5675 (
            .O(N__43183),
            .I(\quad_counter0.n2910 ));
    LocalMux I__5674 (
            .O(N__43180),
            .I(\quad_counter0.n2910 ));
    InMux I__5673 (
            .O(N__43173),
            .I(N__43168));
    InMux I__5672 (
            .O(N__43172),
            .I(N__43165));
    InMux I__5671 (
            .O(N__43171),
            .I(N__43162));
    LocalMux I__5670 (
            .O(N__43168),
            .I(N__43159));
    LocalMux I__5669 (
            .O(N__43165),
            .I(\quad_counter0.n2913 ));
    LocalMux I__5668 (
            .O(N__43162),
            .I(\quad_counter0.n2913 ));
    Odrv4 I__5667 (
            .O(N__43159),
            .I(\quad_counter0.n2913 ));
    CascadeMux I__5666 (
            .O(N__43152),
            .I(N__43147));
    InMux I__5665 (
            .O(N__43151),
            .I(N__43144));
    InMux I__5664 (
            .O(N__43150),
            .I(N__43141));
    InMux I__5663 (
            .O(N__43147),
            .I(N__43138));
    LocalMux I__5662 (
            .O(N__43144),
            .I(\quad_counter0.n2907 ));
    LocalMux I__5661 (
            .O(N__43141),
            .I(\quad_counter0.n2907 ));
    LocalMux I__5660 (
            .O(N__43138),
            .I(\quad_counter0.n2907 ));
    InMux I__5659 (
            .O(N__43131),
            .I(N__43126));
    InMux I__5658 (
            .O(N__43130),
            .I(N__43123));
    InMux I__5657 (
            .O(N__43129),
            .I(N__43120));
    LocalMux I__5656 (
            .O(N__43126),
            .I(\quad_counter0.n2905 ));
    LocalMux I__5655 (
            .O(N__43123),
            .I(\quad_counter0.n2905 ));
    LocalMux I__5654 (
            .O(N__43120),
            .I(\quad_counter0.n2905 ));
    InMux I__5653 (
            .O(N__43113),
            .I(N__43108));
    InMux I__5652 (
            .O(N__43112),
            .I(N__43105));
    InMux I__5651 (
            .O(N__43111),
            .I(N__43102));
    LocalMux I__5650 (
            .O(N__43108),
            .I(N__43099));
    LocalMux I__5649 (
            .O(N__43105),
            .I(\quad_counter0.n2919 ));
    LocalMux I__5648 (
            .O(N__43102),
            .I(\quad_counter0.n2919 ));
    Odrv4 I__5647 (
            .O(N__43099),
            .I(\quad_counter0.n2919 ));
    CascadeMux I__5646 (
            .O(N__43092),
            .I(N__43084));
    CascadeMux I__5645 (
            .O(N__43091),
            .I(N__43081));
    CascadeMux I__5644 (
            .O(N__43090),
            .I(N__43078));
    CascadeMux I__5643 (
            .O(N__43089),
            .I(N__43075));
    CascadeMux I__5642 (
            .O(N__43088),
            .I(N__43072));
    CascadeMux I__5641 (
            .O(N__43087),
            .I(N__43069));
    InMux I__5640 (
            .O(N__43084),
            .I(N__43064));
    InMux I__5639 (
            .O(N__43081),
            .I(N__43064));
    InMux I__5638 (
            .O(N__43078),
            .I(N__43055));
    InMux I__5637 (
            .O(N__43075),
            .I(N__43055));
    InMux I__5636 (
            .O(N__43072),
            .I(N__43055));
    InMux I__5635 (
            .O(N__43069),
            .I(N__43055));
    LocalMux I__5634 (
            .O(N__43064),
            .I(\quad_counter0.n36145 ));
    LocalMux I__5633 (
            .O(N__43055),
            .I(\quad_counter0.n36145 ));
    InMux I__5632 (
            .O(N__43050),
            .I(N__43047));
    LocalMux I__5631 (
            .O(N__43047),
            .I(N__43042));
    InMux I__5630 (
            .O(N__43046),
            .I(N__43039));
    InMux I__5629 (
            .O(N__43045),
            .I(N__43036));
    Span4Mux_h I__5628 (
            .O(N__43042),
            .I(N__43033));
    LocalMux I__5627 (
            .O(N__43039),
            .I(N__43030));
    LocalMux I__5626 (
            .O(N__43036),
            .I(N__43027));
    Odrv4 I__5625 (
            .O(N__43033),
            .I(\quad_counter0.n2912 ));
    Odrv4 I__5624 (
            .O(N__43030),
            .I(\quad_counter0.n2912 ));
    Odrv4 I__5623 (
            .O(N__43027),
            .I(\quad_counter0.n2912 ));
    InMux I__5622 (
            .O(N__43020),
            .I(N__43015));
    InMux I__5621 (
            .O(N__43019),
            .I(N__43012));
    InMux I__5620 (
            .O(N__43018),
            .I(N__43009));
    LocalMux I__5619 (
            .O(N__43015),
            .I(\quad_counter0.n2903 ));
    LocalMux I__5618 (
            .O(N__43012),
            .I(\quad_counter0.n2903 ));
    LocalMux I__5617 (
            .O(N__43009),
            .I(\quad_counter0.n2903 ));
    CascadeMux I__5616 (
            .O(N__43002),
            .I(N__42999));
    InMux I__5615 (
            .O(N__42999),
            .I(N__42996));
    LocalMux I__5614 (
            .O(N__42996),
            .I(\quad_counter0.n20 ));
    InMux I__5613 (
            .O(N__42993),
            .I(\quad_counter0.n30318 ));
    InMux I__5612 (
            .O(N__42990),
            .I(\quad_counter0.n30319 ));
    InMux I__5611 (
            .O(N__42987),
            .I(\quad_counter0.n30320 ));
    InMux I__5610 (
            .O(N__42984),
            .I(bfn_11_15_0_));
    InMux I__5609 (
            .O(N__42981),
            .I(\quad_counter0.n30322 ));
    InMux I__5608 (
            .O(N__42978),
            .I(\quad_counter0.n30323 ));
    InMux I__5607 (
            .O(N__42975),
            .I(\quad_counter0.n30324 ));
    InMux I__5606 (
            .O(N__42972),
            .I(\quad_counter0.n30325 ));
    InMux I__5605 (
            .O(N__42969),
            .I(\quad_counter0.n30326 ));
    InMux I__5604 (
            .O(N__42966),
            .I(N__42962));
    CascadeMux I__5603 (
            .O(N__42965),
            .I(N__42959));
    LocalMux I__5602 (
            .O(N__42962),
            .I(N__42956));
    InMux I__5601 (
            .O(N__42959),
            .I(N__42953));
    Span4Mux_h I__5600 (
            .O(N__42956),
            .I(N__42950));
    LocalMux I__5599 (
            .O(N__42953),
            .I(r_Tx_Data_2));
    Odrv4 I__5598 (
            .O(N__42950),
            .I(r_Tx_Data_2));
    InMux I__5597 (
            .O(N__42945),
            .I(N__42940));
    InMux I__5596 (
            .O(N__42944),
            .I(N__42937));
    InMux I__5595 (
            .O(N__42943),
            .I(N__42934));
    LocalMux I__5594 (
            .O(N__42940),
            .I(N__42930));
    LocalMux I__5593 (
            .O(N__42937),
            .I(N__42927));
    LocalMux I__5592 (
            .O(N__42934),
            .I(N__42924));
    InMux I__5591 (
            .O(N__42933),
            .I(N__42921));
    Span4Mux_v I__5590 (
            .O(N__42930),
            .I(N__42918));
    Span4Mux_v I__5589 (
            .O(N__42927),
            .I(N__42915));
    Span4Mux_v I__5588 (
            .O(N__42924),
            .I(N__42908));
    LocalMux I__5587 (
            .O(N__42921),
            .I(N__42908));
    Span4Mux_h I__5586 (
            .O(N__42918),
            .I(N__42908));
    Span4Mux_h I__5585 (
            .O(N__42915),
            .I(N__42905));
    Odrv4 I__5584 (
            .O(N__42908),
            .I(data_in_3_5));
    Odrv4 I__5583 (
            .O(N__42905),
            .I(data_in_3_5));
    InMux I__5582 (
            .O(N__42900),
            .I(N__42896));
    InMux I__5581 (
            .O(N__42899),
            .I(N__42893));
    LocalMux I__5580 (
            .O(N__42896),
            .I(N__42890));
    LocalMux I__5579 (
            .O(N__42893),
            .I(r_Tx_Data_1));
    Odrv12 I__5578 (
            .O(N__42890),
            .I(r_Tx_Data_1));
    CascadeMux I__5577 (
            .O(N__42885),
            .I(N__42882));
    InMux I__5576 (
            .O(N__42882),
            .I(N__42878));
    InMux I__5575 (
            .O(N__42881),
            .I(N__42875));
    LocalMux I__5574 (
            .O(N__42878),
            .I(N__42872));
    LocalMux I__5573 (
            .O(N__42875),
            .I(N__42869));
    Span4Mux_v I__5572 (
            .O(N__42872),
            .I(N__42866));
    Span4Mux_v I__5571 (
            .O(N__42869),
            .I(N__42863));
    Odrv4 I__5570 (
            .O(N__42866),
            .I(\c0.n11057 ));
    Odrv4 I__5569 (
            .O(N__42863),
            .I(\c0.n11057 ));
    InMux I__5568 (
            .O(N__42858),
            .I(bfn_11_14_0_));
    InMux I__5567 (
            .O(N__42855),
            .I(\quad_counter0.n30314 ));
    InMux I__5566 (
            .O(N__42852),
            .I(\quad_counter0.n30315 ));
    InMux I__5565 (
            .O(N__42849),
            .I(\quad_counter0.n30316 ));
    InMux I__5564 (
            .O(N__42846),
            .I(\quad_counter0.n30317 ));
    InMux I__5563 (
            .O(N__42843),
            .I(N__42838));
    InMux I__5562 (
            .O(N__42842),
            .I(N__42835));
    InMux I__5561 (
            .O(N__42841),
            .I(N__42832));
    LocalMux I__5560 (
            .O(N__42838),
            .I(N__42829));
    LocalMux I__5559 (
            .O(N__42835),
            .I(N__42824));
    LocalMux I__5558 (
            .O(N__42832),
            .I(N__42824));
    Span4Mux_v I__5557 (
            .O(N__42829),
            .I(N__42821));
    Odrv4 I__5556 (
            .O(N__42824),
            .I(\quad_counter0.n3019 ));
    Odrv4 I__5555 (
            .O(N__42821),
            .I(\quad_counter0.n3019 ));
    CascadeMux I__5554 (
            .O(N__42816),
            .I(\quad_counter0.n10_adj_4376_cascade_ ));
    CascadeMux I__5553 (
            .O(N__42813),
            .I(\quad_counter0.n1847_cascade_ ));
    CascadeMux I__5552 (
            .O(N__42810),
            .I(N__42804));
    InMux I__5551 (
            .O(N__42809),
            .I(N__42797));
    InMux I__5550 (
            .O(N__42808),
            .I(N__42797));
    InMux I__5549 (
            .O(N__42807),
            .I(N__42794));
    InMux I__5548 (
            .O(N__42804),
            .I(N__42791));
    InMux I__5547 (
            .O(N__42803),
            .I(N__42786));
    InMux I__5546 (
            .O(N__42802),
            .I(N__42786));
    LocalMux I__5545 (
            .O(N__42797),
            .I(N__42783));
    LocalMux I__5544 (
            .O(N__42794),
            .I(N__42780));
    LocalMux I__5543 (
            .O(N__42791),
            .I(r_Bit_Index_1));
    LocalMux I__5542 (
            .O(N__42786),
            .I(r_Bit_Index_1));
    Odrv4 I__5541 (
            .O(N__42783),
            .I(r_Bit_Index_1));
    Odrv12 I__5540 (
            .O(N__42780),
            .I(r_Bit_Index_1));
    InMux I__5539 (
            .O(N__42771),
            .I(N__42768));
    LocalMux I__5538 (
            .O(N__42768),
            .I(N__42765));
    Span4Mux_h I__5537 (
            .O(N__42765),
            .I(N__42762));
    Span4Mux_v I__5536 (
            .O(N__42762),
            .I(N__42758));
    InMux I__5535 (
            .O(N__42761),
            .I(N__42755));
    Span4Mux_v I__5534 (
            .O(N__42758),
            .I(N__42752));
    LocalMux I__5533 (
            .O(N__42755),
            .I(r_Tx_Data_4));
    Odrv4 I__5532 (
            .O(N__42752),
            .I(r_Tx_Data_4));
    CascadeMux I__5531 (
            .O(N__42747),
            .I(N__42743));
    CascadeMux I__5530 (
            .O(N__42746),
            .I(N__42739));
    InMux I__5529 (
            .O(N__42743),
            .I(N__42736));
    InMux I__5528 (
            .O(N__42742),
            .I(N__42733));
    InMux I__5527 (
            .O(N__42739),
            .I(N__42730));
    LocalMux I__5526 (
            .O(N__42736),
            .I(N__42725));
    LocalMux I__5525 (
            .O(N__42733),
            .I(N__42722));
    LocalMux I__5524 (
            .O(N__42730),
            .I(N__42717));
    InMux I__5523 (
            .O(N__42729),
            .I(N__42712));
    InMux I__5522 (
            .O(N__42728),
            .I(N__42712));
    Span4Mux_h I__5521 (
            .O(N__42725),
            .I(N__42709));
    Span4Mux_h I__5520 (
            .O(N__42722),
            .I(N__42706));
    InMux I__5519 (
            .O(N__42721),
            .I(N__42703));
    InMux I__5518 (
            .O(N__42720),
            .I(N__42700));
    Span4Mux_v I__5517 (
            .O(N__42717),
            .I(N__42697));
    LocalMux I__5516 (
            .O(N__42712),
            .I(N__42692));
    Span4Mux_h I__5515 (
            .O(N__42709),
            .I(N__42692));
    Span4Mux_h I__5514 (
            .O(N__42706),
            .I(N__42689));
    LocalMux I__5513 (
            .O(N__42703),
            .I(r_Bit_Index_0));
    LocalMux I__5512 (
            .O(N__42700),
            .I(r_Bit_Index_0));
    Odrv4 I__5511 (
            .O(N__42697),
            .I(r_Bit_Index_0));
    Odrv4 I__5510 (
            .O(N__42692),
            .I(r_Bit_Index_0));
    Odrv4 I__5509 (
            .O(N__42689),
            .I(r_Bit_Index_0));
    InMux I__5508 (
            .O(N__42678),
            .I(N__42675));
    LocalMux I__5507 (
            .O(N__42675),
            .I(\c0.n36167 ));
    InMux I__5506 (
            .O(N__42672),
            .I(N__42669));
    LocalMux I__5505 (
            .O(N__42669),
            .I(N__42666));
    Span4Mux_h I__5504 (
            .O(N__42666),
            .I(N__42663));
    Odrv4 I__5503 (
            .O(N__42663),
            .I(\c0.n36170 ));
    InMux I__5502 (
            .O(N__42660),
            .I(N__42653));
    InMux I__5501 (
            .O(N__42659),
            .I(N__42653));
    InMux I__5500 (
            .O(N__42658),
            .I(N__42650));
    LocalMux I__5499 (
            .O(N__42653),
            .I(N__42647));
    LocalMux I__5498 (
            .O(N__42650),
            .I(N__42644));
    Odrv12 I__5497 (
            .O(N__42647),
            .I(\c0.n10_adj_4629 ));
    Odrv4 I__5496 (
            .O(N__42644),
            .I(\c0.n10_adj_4629 ));
    InMux I__5495 (
            .O(N__42639),
            .I(N__42634));
    InMux I__5494 (
            .O(N__42638),
            .I(N__42631));
    InMux I__5493 (
            .O(N__42637),
            .I(N__42628));
    LocalMux I__5492 (
            .O(N__42634),
            .I(N__42623));
    LocalMux I__5491 (
            .O(N__42631),
            .I(N__42623));
    LocalMux I__5490 (
            .O(N__42628),
            .I(N__42620));
    Odrv4 I__5489 (
            .O(N__42623),
            .I(\quad_counter0.n3018 ));
    Odrv4 I__5488 (
            .O(N__42620),
            .I(\quad_counter0.n3018 ));
    InMux I__5487 (
            .O(N__42615),
            .I(N__42610));
    InMux I__5486 (
            .O(N__42614),
            .I(N__42607));
    InMux I__5485 (
            .O(N__42613),
            .I(N__42604));
    LocalMux I__5484 (
            .O(N__42610),
            .I(N__42599));
    LocalMux I__5483 (
            .O(N__42607),
            .I(N__42599));
    LocalMux I__5482 (
            .O(N__42604),
            .I(N__42596));
    Odrv4 I__5481 (
            .O(N__42599),
            .I(\quad_counter0.n3014 ));
    Odrv4 I__5480 (
            .O(N__42596),
            .I(\quad_counter0.n3014 ));
    CascadeMux I__5479 (
            .O(N__42591),
            .I(N__42586));
    InMux I__5478 (
            .O(N__42590),
            .I(N__42583));
    InMux I__5477 (
            .O(N__42589),
            .I(N__42580));
    InMux I__5476 (
            .O(N__42586),
            .I(N__42577));
    LocalMux I__5475 (
            .O(N__42583),
            .I(N__42572));
    LocalMux I__5474 (
            .O(N__42580),
            .I(N__42572));
    LocalMux I__5473 (
            .O(N__42577),
            .I(N__42569));
    Odrv4 I__5472 (
            .O(N__42572),
            .I(\quad_counter0.n3017 ));
    Odrv4 I__5471 (
            .O(N__42569),
            .I(\quad_counter0.n3017 ));
    InMux I__5470 (
            .O(N__42564),
            .I(N__42561));
    LocalMux I__5469 (
            .O(N__42561),
            .I(N__42558));
    Odrv4 I__5468 (
            .O(N__42558),
            .I(\quad_counter0.n28307 ));
    InMux I__5467 (
            .O(N__42555),
            .I(N__42552));
    LocalMux I__5466 (
            .O(N__42552),
            .I(N__42549));
    Span4Mux_h I__5465 (
            .O(N__42549),
            .I(N__42546));
    Odrv4 I__5464 (
            .O(N__42546),
            .I(\quad_counter0.n10_adj_4349 ));
    InMux I__5463 (
            .O(N__42543),
            .I(N__42539));
    InMux I__5462 (
            .O(N__42542),
            .I(N__42536));
    LocalMux I__5461 (
            .O(N__42539),
            .I(N__42533));
    LocalMux I__5460 (
            .O(N__42536),
            .I(\quad_counter1.b_delay_counter_10 ));
    Odrv4 I__5459 (
            .O(N__42533),
            .I(\quad_counter1.b_delay_counter_10 ));
    InMux I__5458 (
            .O(N__42528),
            .I(\quad_counter1.n30040 ));
    InMux I__5457 (
            .O(N__42525),
            .I(N__42521));
    InMux I__5456 (
            .O(N__42524),
            .I(N__42518));
    LocalMux I__5455 (
            .O(N__42521),
            .I(N__42515));
    LocalMux I__5454 (
            .O(N__42518),
            .I(\quad_counter1.b_delay_counter_11 ));
    Odrv4 I__5453 (
            .O(N__42515),
            .I(\quad_counter1.b_delay_counter_11 ));
    InMux I__5452 (
            .O(N__42510),
            .I(\quad_counter1.n30041 ));
    InMux I__5451 (
            .O(N__42507),
            .I(N__42503));
    InMux I__5450 (
            .O(N__42506),
            .I(N__42500));
    LocalMux I__5449 (
            .O(N__42503),
            .I(N__42497));
    LocalMux I__5448 (
            .O(N__42500),
            .I(\quad_counter1.b_delay_counter_12 ));
    Odrv4 I__5447 (
            .O(N__42497),
            .I(\quad_counter1.b_delay_counter_12 ));
    InMux I__5446 (
            .O(N__42492),
            .I(\quad_counter1.n30042 ));
    InMux I__5445 (
            .O(N__42489),
            .I(N__42485));
    InMux I__5444 (
            .O(N__42488),
            .I(N__42482));
    LocalMux I__5443 (
            .O(N__42485),
            .I(N__42479));
    LocalMux I__5442 (
            .O(N__42482),
            .I(\quad_counter1.b_delay_counter_13 ));
    Odrv4 I__5441 (
            .O(N__42479),
            .I(\quad_counter1.b_delay_counter_13 ));
    InMux I__5440 (
            .O(N__42474),
            .I(\quad_counter1.n30043 ));
    InMux I__5439 (
            .O(N__42471),
            .I(N__42467));
    InMux I__5438 (
            .O(N__42470),
            .I(N__42464));
    LocalMux I__5437 (
            .O(N__42467),
            .I(N__42461));
    LocalMux I__5436 (
            .O(N__42464),
            .I(\quad_counter1.b_delay_counter_14 ));
    Odrv4 I__5435 (
            .O(N__42461),
            .I(\quad_counter1.b_delay_counter_14 ));
    InMux I__5434 (
            .O(N__42456),
            .I(\quad_counter1.n30044 ));
    InMux I__5433 (
            .O(N__42453),
            .I(\quad_counter1.n30045 ));
    InMux I__5432 (
            .O(N__42450),
            .I(N__42446));
    InMux I__5431 (
            .O(N__42449),
            .I(N__42443));
    LocalMux I__5430 (
            .O(N__42446),
            .I(N__42440));
    LocalMux I__5429 (
            .O(N__42443),
            .I(\quad_counter1.b_delay_counter_15 ));
    Odrv4 I__5428 (
            .O(N__42440),
            .I(\quad_counter1.b_delay_counter_15 ));
    CEMux I__5427 (
            .O(N__42435),
            .I(N__42432));
    LocalMux I__5426 (
            .O(N__42432),
            .I(N__42428));
    CEMux I__5425 (
            .O(N__42431),
            .I(N__42425));
    Span4Mux_h I__5424 (
            .O(N__42428),
            .I(N__42422));
    LocalMux I__5423 (
            .O(N__42425),
            .I(N__42419));
    Odrv4 I__5422 (
            .O(N__42422),
            .I(n19463));
    Odrv4 I__5421 (
            .O(N__42419),
            .I(n19463));
    SRMux I__5420 (
            .O(N__42414),
            .I(N__42411));
    LocalMux I__5419 (
            .O(N__42411),
            .I(N__42407));
    SRMux I__5418 (
            .O(N__42410),
            .I(N__42404));
    Span4Mux_v I__5417 (
            .O(N__42407),
            .I(N__42401));
    LocalMux I__5416 (
            .O(N__42404),
            .I(N__42398));
    Odrv4 I__5415 (
            .O(N__42401),
            .I(\quad_counter1.b_delay_counter_15__N_4237 ));
    Odrv12 I__5414 (
            .O(N__42398),
            .I(\quad_counter1.b_delay_counter_15__N_4237 ));
    InMux I__5413 (
            .O(N__42393),
            .I(N__42390));
    LocalMux I__5412 (
            .O(N__42390),
            .I(N__42385));
    InMux I__5411 (
            .O(N__42389),
            .I(N__42382));
    InMux I__5410 (
            .O(N__42388),
            .I(N__42379));
    Span4Mux_v I__5409 (
            .O(N__42385),
            .I(N__42376));
    LocalMux I__5408 (
            .O(N__42382),
            .I(N__42371));
    LocalMux I__5407 (
            .O(N__42379),
            .I(N__42371));
    Odrv4 I__5406 (
            .O(N__42376),
            .I(\quad_counter0.n3219 ));
    Odrv4 I__5405 (
            .O(N__42371),
            .I(\quad_counter0.n3219 ));
    InMux I__5404 (
            .O(N__42366),
            .I(N__42361));
    InMux I__5403 (
            .O(N__42365),
            .I(N__42358));
    InMux I__5402 (
            .O(N__42364),
            .I(N__42355));
    LocalMux I__5401 (
            .O(N__42361),
            .I(N__42352));
    LocalMux I__5400 (
            .O(N__42358),
            .I(N__42347));
    LocalMux I__5399 (
            .O(N__42355),
            .I(N__42347));
    Odrv4 I__5398 (
            .O(N__42352),
            .I(\quad_counter0.n3218 ));
    Odrv4 I__5397 (
            .O(N__42347),
            .I(\quad_counter0.n3218 ));
    InMux I__5396 (
            .O(N__42342),
            .I(N__42337));
    InMux I__5395 (
            .O(N__42341),
            .I(N__42334));
    InMux I__5394 (
            .O(N__42340),
            .I(N__42331));
    LocalMux I__5393 (
            .O(N__42337),
            .I(N__42326));
    LocalMux I__5392 (
            .O(N__42334),
            .I(N__42326));
    LocalMux I__5391 (
            .O(N__42331),
            .I(N__42323));
    Odrv4 I__5390 (
            .O(N__42326),
            .I(\quad_counter0.n3217 ));
    Odrv4 I__5389 (
            .O(N__42323),
            .I(\quad_counter0.n3217 ));
    CascadeMux I__5388 (
            .O(N__42318),
            .I(\quad_counter0.n28297_cascade_ ));
    InMux I__5387 (
            .O(N__42315),
            .I(N__42310));
    InMux I__5386 (
            .O(N__42314),
            .I(N__42307));
    InMux I__5385 (
            .O(N__42313),
            .I(N__42304));
    LocalMux I__5384 (
            .O(N__42310),
            .I(N__42301));
    LocalMux I__5383 (
            .O(N__42307),
            .I(N__42296));
    LocalMux I__5382 (
            .O(N__42304),
            .I(N__42296));
    Odrv4 I__5381 (
            .O(N__42301),
            .I(\quad_counter0.n3214 ));
    Odrv4 I__5380 (
            .O(N__42296),
            .I(\quad_counter0.n3214 ));
    CascadeMux I__5379 (
            .O(N__42291),
            .I(N__42288));
    InMux I__5378 (
            .O(N__42288),
            .I(N__42285));
    LocalMux I__5377 (
            .O(N__42285),
            .I(N__42282));
    Odrv4 I__5376 (
            .O(N__42282),
            .I(\quad_counter0.n10_adj_4357 ));
    InMux I__5375 (
            .O(N__42279),
            .I(N__42275));
    InMux I__5374 (
            .O(N__42278),
            .I(N__42272));
    LocalMux I__5373 (
            .O(N__42275),
            .I(\quad_counter1.b_delay_counter_2 ));
    LocalMux I__5372 (
            .O(N__42272),
            .I(\quad_counter1.b_delay_counter_2 ));
    InMux I__5371 (
            .O(N__42267),
            .I(\quad_counter1.n30032 ));
    InMux I__5370 (
            .O(N__42264),
            .I(N__42260));
    InMux I__5369 (
            .O(N__42263),
            .I(N__42257));
    LocalMux I__5368 (
            .O(N__42260),
            .I(\quad_counter1.b_delay_counter_3 ));
    LocalMux I__5367 (
            .O(N__42257),
            .I(\quad_counter1.b_delay_counter_3 ));
    InMux I__5366 (
            .O(N__42252),
            .I(\quad_counter1.n30033 ));
    InMux I__5365 (
            .O(N__42249),
            .I(N__42245));
    InMux I__5364 (
            .O(N__42248),
            .I(N__42242));
    LocalMux I__5363 (
            .O(N__42245),
            .I(\quad_counter1.b_delay_counter_4 ));
    LocalMux I__5362 (
            .O(N__42242),
            .I(\quad_counter1.b_delay_counter_4 ));
    InMux I__5361 (
            .O(N__42237),
            .I(\quad_counter1.n30034 ));
    InMux I__5360 (
            .O(N__42234),
            .I(N__42230));
    InMux I__5359 (
            .O(N__42233),
            .I(N__42227));
    LocalMux I__5358 (
            .O(N__42230),
            .I(\quad_counter1.b_delay_counter_5 ));
    LocalMux I__5357 (
            .O(N__42227),
            .I(\quad_counter1.b_delay_counter_5 ));
    InMux I__5356 (
            .O(N__42222),
            .I(\quad_counter1.n30035 ));
    InMux I__5355 (
            .O(N__42219),
            .I(N__42215));
    InMux I__5354 (
            .O(N__42218),
            .I(N__42212));
    LocalMux I__5353 (
            .O(N__42215),
            .I(\quad_counter1.b_delay_counter_6 ));
    LocalMux I__5352 (
            .O(N__42212),
            .I(\quad_counter1.b_delay_counter_6 ));
    InMux I__5351 (
            .O(N__42207),
            .I(\quad_counter1.n30036 ));
    CascadeMux I__5350 (
            .O(N__42204),
            .I(N__42200));
    InMux I__5349 (
            .O(N__42203),
            .I(N__42197));
    InMux I__5348 (
            .O(N__42200),
            .I(N__42194));
    LocalMux I__5347 (
            .O(N__42197),
            .I(\quad_counter1.b_delay_counter_7 ));
    LocalMux I__5346 (
            .O(N__42194),
            .I(\quad_counter1.b_delay_counter_7 ));
    InMux I__5345 (
            .O(N__42189),
            .I(\quad_counter1.n30037 ));
    CascadeMux I__5344 (
            .O(N__42186),
            .I(N__42183));
    InMux I__5343 (
            .O(N__42183),
            .I(N__42179));
    InMux I__5342 (
            .O(N__42182),
            .I(N__42176));
    LocalMux I__5341 (
            .O(N__42179),
            .I(N__42173));
    LocalMux I__5340 (
            .O(N__42176),
            .I(\quad_counter1.b_delay_counter_8 ));
    Odrv4 I__5339 (
            .O(N__42173),
            .I(\quad_counter1.b_delay_counter_8 ));
    InMux I__5338 (
            .O(N__42168),
            .I(bfn_11_8_0_));
    InMux I__5337 (
            .O(N__42165),
            .I(N__42161));
    InMux I__5336 (
            .O(N__42164),
            .I(N__42158));
    LocalMux I__5335 (
            .O(N__42161),
            .I(N__42155));
    LocalMux I__5334 (
            .O(N__42158),
            .I(\quad_counter1.b_delay_counter_9 ));
    Odrv4 I__5333 (
            .O(N__42155),
            .I(\quad_counter1.b_delay_counter_9 ));
    InMux I__5332 (
            .O(N__42150),
            .I(\quad_counter1.n30039 ));
    InMux I__5331 (
            .O(N__42147),
            .I(N__42137));
    InMux I__5330 (
            .O(N__42146),
            .I(N__42137));
    InMux I__5329 (
            .O(N__42145),
            .I(N__42137));
    InMux I__5328 (
            .O(N__42144),
            .I(N__42134));
    LocalMux I__5327 (
            .O(N__42137),
            .I(N__42129));
    LocalMux I__5326 (
            .O(N__42134),
            .I(N__42129));
    Span4Mux_v I__5325 (
            .O(N__42129),
            .I(N__42126));
    Sp12to4 I__5324 (
            .O(N__42126),
            .I(N__42123));
    Odrv12 I__5323 (
            .O(N__42123),
            .I(PIN_13_c));
    InMux I__5322 (
            .O(N__42120),
            .I(N__42111));
    InMux I__5321 (
            .O(N__42119),
            .I(N__42111));
    InMux I__5320 (
            .O(N__42118),
            .I(N__42111));
    LocalMux I__5319 (
            .O(N__42111),
            .I(quadB_delayed_adj_4813));
    CascadeMux I__5318 (
            .O(N__42108),
            .I(\quad_counter1.n26_adj_4447_cascade_ ));
    CascadeMux I__5317 (
            .O(N__42105),
            .I(N__42102));
    InMux I__5316 (
            .O(N__42102),
            .I(N__42096));
    InMux I__5315 (
            .O(N__42101),
            .I(N__42096));
    LocalMux I__5314 (
            .O(N__42096),
            .I(n17983));
    InMux I__5313 (
            .O(N__42093),
            .I(N__42090));
    LocalMux I__5312 (
            .O(N__42090),
            .I(\quad_counter1.n27_adj_4448 ));
    InMux I__5311 (
            .O(N__42087),
            .I(N__42084));
    LocalMux I__5310 (
            .O(N__42084),
            .I(\quad_counter1.n25_adj_4449 ));
    InMux I__5309 (
            .O(N__42081),
            .I(N__42078));
    LocalMux I__5308 (
            .O(N__42078),
            .I(\quad_counter1.n28_adj_4446 ));
    CascadeMux I__5307 (
            .O(N__42075),
            .I(N__42071));
    InMux I__5306 (
            .O(N__42074),
            .I(N__42068));
    InMux I__5305 (
            .O(N__42071),
            .I(N__42065));
    LocalMux I__5304 (
            .O(N__42068),
            .I(\quad_counter1.b_delay_counter_0 ));
    LocalMux I__5303 (
            .O(N__42065),
            .I(\quad_counter1.b_delay_counter_0 ));
    InMux I__5302 (
            .O(N__42060),
            .I(bfn_11_7_0_));
    CascadeMux I__5301 (
            .O(N__42057),
            .I(N__42053));
    InMux I__5300 (
            .O(N__42056),
            .I(N__42050));
    InMux I__5299 (
            .O(N__42053),
            .I(N__42047));
    LocalMux I__5298 (
            .O(N__42050),
            .I(\quad_counter1.b_delay_counter_1 ));
    LocalMux I__5297 (
            .O(N__42047),
            .I(\quad_counter1.b_delay_counter_1 ));
    InMux I__5296 (
            .O(N__42042),
            .I(\quad_counter1.n30031 ));
    CascadeMux I__5295 (
            .O(N__42039),
            .I(N__42034));
    InMux I__5294 (
            .O(N__42038),
            .I(N__42028));
    InMux I__5293 (
            .O(N__42037),
            .I(N__42028));
    InMux I__5292 (
            .O(N__42034),
            .I(N__42025));
    InMux I__5291 (
            .O(N__42033),
            .I(N__42022));
    LocalMux I__5290 (
            .O(N__42028),
            .I(N__42019));
    LocalMux I__5289 (
            .O(N__42025),
            .I(\c0.data_in_frame_10_6 ));
    LocalMux I__5288 (
            .O(N__42022),
            .I(\c0.data_in_frame_10_6 ));
    Odrv4 I__5287 (
            .O(N__42019),
            .I(\c0.data_in_frame_10_6 ));
    CascadeMux I__5286 (
            .O(N__42012),
            .I(\c0.n6_adj_4539_cascade_ ));
    CascadeMux I__5285 (
            .O(N__42009),
            .I(\c0.n19199_cascade_ ));
    InMux I__5284 (
            .O(N__42006),
            .I(N__42002));
    CascadeMux I__5283 (
            .O(N__42005),
            .I(N__41998));
    LocalMux I__5282 (
            .O(N__42002),
            .I(N__41995));
    InMux I__5281 (
            .O(N__42001),
            .I(N__41992));
    InMux I__5280 (
            .O(N__41998),
            .I(N__41989));
    Span4Mux_h I__5279 (
            .O(N__41995),
            .I(N__41986));
    LocalMux I__5278 (
            .O(N__41992),
            .I(N__41983));
    LocalMux I__5277 (
            .O(N__41989),
            .I(\c0.data_in_frame_11_4 ));
    Odrv4 I__5276 (
            .O(N__41986),
            .I(\c0.data_in_frame_11_4 ));
    Odrv4 I__5275 (
            .O(N__41983),
            .I(\c0.data_in_frame_11_4 ));
    CascadeMux I__5274 (
            .O(N__41976),
            .I(N__41973));
    InMux I__5273 (
            .O(N__41973),
            .I(N__41970));
    LocalMux I__5272 (
            .O(N__41970),
            .I(N__41967));
    Span4Mux_v I__5271 (
            .O(N__41967),
            .I(N__41962));
    InMux I__5270 (
            .O(N__41966),
            .I(N__41957));
    InMux I__5269 (
            .O(N__41965),
            .I(N__41957));
    Odrv4 I__5268 (
            .O(N__41962),
            .I(\c0.data_in_frame_11_3 ));
    LocalMux I__5267 (
            .O(N__41957),
            .I(\c0.data_in_frame_11_3 ));
    CascadeMux I__5266 (
            .O(N__41952),
            .I(N__41948));
    InMux I__5265 (
            .O(N__41951),
            .I(N__41945));
    InMux I__5264 (
            .O(N__41948),
            .I(N__41942));
    LocalMux I__5263 (
            .O(N__41945),
            .I(N__41939));
    LocalMux I__5262 (
            .O(N__41942),
            .I(\c0.data_in_frame_11_6 ));
    Odrv4 I__5261 (
            .O(N__41939),
            .I(\c0.data_in_frame_11_6 ));
    CascadeMux I__5260 (
            .O(N__41934),
            .I(N__41931));
    InMux I__5259 (
            .O(N__41931),
            .I(N__41926));
    InMux I__5258 (
            .O(N__41930),
            .I(N__41921));
    InMux I__5257 (
            .O(N__41929),
            .I(N__41921));
    LocalMux I__5256 (
            .O(N__41926),
            .I(\c0.data_in_frame_9_4 ));
    LocalMux I__5255 (
            .O(N__41921),
            .I(\c0.data_in_frame_9_4 ));
    CascadeMux I__5254 (
            .O(N__41916),
            .I(N__41913));
    InMux I__5253 (
            .O(N__41913),
            .I(N__41910));
    LocalMux I__5252 (
            .O(N__41910),
            .I(N__41907));
    Odrv4 I__5251 (
            .O(N__41907),
            .I(\c0.n33641 ));
    InMux I__5250 (
            .O(N__41904),
            .I(N__41901));
    LocalMux I__5249 (
            .O(N__41901),
            .I(N__41896));
    InMux I__5248 (
            .O(N__41900),
            .I(N__41893));
    CascadeMux I__5247 (
            .O(N__41899),
            .I(N__41890));
    Span4Mux_v I__5246 (
            .O(N__41896),
            .I(N__41885));
    LocalMux I__5245 (
            .O(N__41893),
            .I(N__41885));
    InMux I__5244 (
            .O(N__41890),
            .I(N__41882));
    Span4Mux_h I__5243 (
            .O(N__41885),
            .I(N__41879));
    LocalMux I__5242 (
            .O(N__41882),
            .I(\c0.data_in_frame_7_3 ));
    Odrv4 I__5241 (
            .O(N__41879),
            .I(\c0.data_in_frame_7_3 ));
    InMux I__5240 (
            .O(N__41874),
            .I(N__41871));
    LocalMux I__5239 (
            .O(N__41871),
            .I(N__41868));
    Odrv4 I__5238 (
            .O(N__41868),
            .I(\c0.n31505 ));
    CascadeMux I__5237 (
            .O(N__41865),
            .I(\c0.n33641_cascade_ ));
    InMux I__5236 (
            .O(N__41862),
            .I(N__41858));
    InMux I__5235 (
            .O(N__41861),
            .I(N__41855));
    LocalMux I__5234 (
            .O(N__41858),
            .I(N__41852));
    LocalMux I__5233 (
            .O(N__41855),
            .I(N__41849));
    Odrv12 I__5232 (
            .O(N__41852),
            .I(\c0.n33836 ));
    Odrv4 I__5231 (
            .O(N__41849),
            .I(\c0.n33836 ));
    InMux I__5230 (
            .O(N__41844),
            .I(N__41841));
    LocalMux I__5229 (
            .O(N__41841),
            .I(N__41838));
    Span4Mux_h I__5228 (
            .O(N__41838),
            .I(N__41835));
    Odrv4 I__5227 (
            .O(N__41835),
            .I(\c0.n6_adj_4557 ));
    InMux I__5226 (
            .O(N__41832),
            .I(N__41829));
    LocalMux I__5225 (
            .O(N__41829),
            .I(\c0.n33982 ));
    CascadeMux I__5224 (
            .O(N__41826),
            .I(\c0.n18_adj_4725_cascade_ ));
    InMux I__5223 (
            .O(N__41823),
            .I(N__41819));
    InMux I__5222 (
            .O(N__41822),
            .I(N__41816));
    LocalMux I__5221 (
            .O(N__41819),
            .I(N__41813));
    LocalMux I__5220 (
            .O(N__41816),
            .I(\c0.n33951 ));
    Odrv4 I__5219 (
            .O(N__41813),
            .I(\c0.n33951 ));
    InMux I__5218 (
            .O(N__41808),
            .I(N__41805));
    LocalMux I__5217 (
            .O(N__41805),
            .I(N__41802));
    Span4Mux_h I__5216 (
            .O(N__41802),
            .I(N__41799));
    Odrv4 I__5215 (
            .O(N__41799),
            .I(\c0.n16_adj_4726 ));
    CascadeMux I__5214 (
            .O(N__41796),
            .I(\c0.n20_adj_4727_cascade_ ));
    InMux I__5213 (
            .O(N__41793),
            .I(N__41788));
    InMux I__5212 (
            .O(N__41792),
            .I(N__41785));
    CascadeMux I__5211 (
            .O(N__41791),
            .I(N__41782));
    LocalMux I__5210 (
            .O(N__41788),
            .I(N__41778));
    LocalMux I__5209 (
            .O(N__41785),
            .I(N__41775));
    InMux I__5208 (
            .O(N__41782),
            .I(N__41770));
    InMux I__5207 (
            .O(N__41781),
            .I(N__41770));
    Odrv4 I__5206 (
            .O(N__41778),
            .I(\c0.data_in_frame_8_6 ));
    Odrv4 I__5205 (
            .O(N__41775),
            .I(\c0.data_in_frame_8_6 ));
    LocalMux I__5204 (
            .O(N__41770),
            .I(\c0.data_in_frame_8_6 ));
    InMux I__5203 (
            .O(N__41763),
            .I(N__41759));
    InMux I__5202 (
            .O(N__41762),
            .I(N__41755));
    LocalMux I__5201 (
            .O(N__41759),
            .I(N__41752));
    InMux I__5200 (
            .O(N__41758),
            .I(N__41749));
    LocalMux I__5199 (
            .O(N__41755),
            .I(\c0.data_in_frame_8_4 ));
    Odrv4 I__5198 (
            .O(N__41752),
            .I(\c0.data_in_frame_8_4 ));
    LocalMux I__5197 (
            .O(N__41749),
            .I(\c0.data_in_frame_8_4 ));
    InMux I__5196 (
            .O(N__41742),
            .I(N__41739));
    LocalMux I__5195 (
            .O(N__41739),
            .I(\c0.n33723 ));
    CascadeMux I__5194 (
            .O(N__41736),
            .I(\c0.n33723_cascade_ ));
    InMux I__5193 (
            .O(N__41733),
            .I(N__41730));
    LocalMux I__5192 (
            .O(N__41730),
            .I(N__41725));
    InMux I__5191 (
            .O(N__41729),
            .I(N__41720));
    InMux I__5190 (
            .O(N__41728),
            .I(N__41720));
    Span4Mux_h I__5189 (
            .O(N__41725),
            .I(N__41714));
    LocalMux I__5188 (
            .O(N__41720),
            .I(N__41714));
    InMux I__5187 (
            .O(N__41719),
            .I(N__41710));
    Span4Mux_h I__5186 (
            .O(N__41714),
            .I(N__41707));
    InMux I__5185 (
            .O(N__41713),
            .I(N__41704));
    LocalMux I__5184 (
            .O(N__41710),
            .I(\c0.data_in_frame_12_7 ));
    Odrv4 I__5183 (
            .O(N__41707),
            .I(\c0.data_in_frame_12_7 ));
    LocalMux I__5182 (
            .O(N__41704),
            .I(\c0.data_in_frame_12_7 ));
    InMux I__5181 (
            .O(N__41697),
            .I(N__41694));
    LocalMux I__5180 (
            .O(N__41694),
            .I(\c0.n48 ));
    CascadeMux I__5179 (
            .O(N__41691),
            .I(\c0.n6_adj_4556_cascade_ ));
    InMux I__5178 (
            .O(N__41688),
            .I(N__41684));
    InMux I__5177 (
            .O(N__41687),
            .I(N__41681));
    LocalMux I__5176 (
            .O(N__41684),
            .I(\c0.n33404 ));
    LocalMux I__5175 (
            .O(N__41681),
            .I(\c0.n33404 ));
    CascadeMux I__5174 (
            .O(N__41676),
            .I(\c0.n12_adj_4735_cascade_ ));
    CascadeMux I__5173 (
            .O(N__41673),
            .I(\c0.n31526_cascade_ ));
    InMux I__5172 (
            .O(N__41670),
            .I(N__41667));
    LocalMux I__5171 (
            .O(N__41667),
            .I(\c0.n33624 ));
    InMux I__5170 (
            .O(N__41664),
            .I(N__41661));
    LocalMux I__5169 (
            .O(N__41661),
            .I(N__41658));
    Span4Mux_h I__5168 (
            .O(N__41658),
            .I(N__41655));
    Odrv4 I__5167 (
            .O(N__41655),
            .I(\c0.n5860 ));
    InMux I__5166 (
            .O(N__41652),
            .I(N__41649));
    LocalMux I__5165 (
            .O(N__41649),
            .I(N__41645));
    InMux I__5164 (
            .O(N__41648),
            .I(N__41642));
    Odrv4 I__5163 (
            .O(N__41645),
            .I(\c0.n33883 ));
    LocalMux I__5162 (
            .O(N__41642),
            .I(\c0.n33883 ));
    InMux I__5161 (
            .O(N__41637),
            .I(N__41634));
    LocalMux I__5160 (
            .O(N__41634),
            .I(\c0.n44_adj_4731 ));
    InMux I__5159 (
            .O(N__41631),
            .I(N__41627));
    CascadeMux I__5158 (
            .O(N__41630),
            .I(N__41624));
    LocalMux I__5157 (
            .O(N__41627),
            .I(N__41621));
    InMux I__5156 (
            .O(N__41624),
            .I(N__41618));
    Span4Mux_v I__5155 (
            .O(N__41621),
            .I(N__41615));
    LocalMux I__5154 (
            .O(N__41618),
            .I(N__41612));
    Odrv4 I__5153 (
            .O(N__41615),
            .I(\c0.n33800 ));
    Odrv12 I__5152 (
            .O(N__41612),
            .I(\c0.n33800 ));
    CascadeMux I__5151 (
            .O(N__41607),
            .I(\c0.n33720_cascade_ ));
    CascadeMux I__5150 (
            .O(N__41604),
            .I(\c0.n17559_cascade_ ));
    InMux I__5149 (
            .O(N__41601),
            .I(N__41597));
    InMux I__5148 (
            .O(N__41600),
            .I(N__41594));
    LocalMux I__5147 (
            .O(N__41597),
            .I(N__41591));
    LocalMux I__5146 (
            .O(N__41594),
            .I(\c0.data_in_frame_9_5 ));
    Odrv12 I__5145 (
            .O(N__41591),
            .I(\c0.data_in_frame_9_5 ));
    CascadeMux I__5144 (
            .O(N__41586),
            .I(\c0.n18544_cascade_ ));
    CascadeMux I__5143 (
            .O(N__41583),
            .I(\c0.n31505_cascade_ ));
    CascadeMux I__5142 (
            .O(N__41580),
            .I(N__41577));
    InMux I__5141 (
            .O(N__41577),
            .I(N__41571));
    InMux I__5140 (
            .O(N__41576),
            .I(N__41571));
    LocalMux I__5139 (
            .O(N__41571),
            .I(N__41568));
    Span4Mux_h I__5138 (
            .O(N__41568),
            .I(N__41565));
    Odrv4 I__5137 (
            .O(N__41565),
            .I(\c0.n4_adj_4548 ));
    CascadeMux I__5136 (
            .O(N__41562),
            .I(\c0.n43_adj_4732_cascade_ ));
    InMux I__5135 (
            .O(N__41559),
            .I(N__41555));
    InMux I__5134 (
            .O(N__41558),
            .I(N__41552));
    LocalMux I__5133 (
            .O(N__41555),
            .I(N__41549));
    LocalMux I__5132 (
            .O(N__41552),
            .I(\c0.n33778 ));
    Odrv12 I__5131 (
            .O(N__41549),
            .I(\c0.n33778 ));
    InMux I__5130 (
            .O(N__41544),
            .I(N__41541));
    LocalMux I__5129 (
            .O(N__41541),
            .I(\c0.n46_adj_4728 ));
    InMux I__5128 (
            .O(N__41538),
            .I(N__41535));
    LocalMux I__5127 (
            .O(N__41535),
            .I(\c0.n47_adj_4729 ));
    CascadeMux I__5126 (
            .O(N__41532),
            .I(\c0.n45_adj_4730_cascade_ ));
    InMux I__5125 (
            .O(N__41529),
            .I(N__41526));
    LocalMux I__5124 (
            .O(N__41526),
            .I(\c0.n54 ));
    InMux I__5123 (
            .O(N__41523),
            .I(N__41519));
    InMux I__5122 (
            .O(N__41522),
            .I(N__41516));
    LocalMux I__5121 (
            .O(N__41519),
            .I(N__41513));
    LocalMux I__5120 (
            .O(N__41516),
            .I(N__41510));
    Odrv4 I__5119 (
            .O(N__41513),
            .I(\c0.n17559 ));
    Odrv4 I__5118 (
            .O(N__41510),
            .I(\c0.n17559 ));
    InMux I__5117 (
            .O(N__41505),
            .I(N__41501));
    InMux I__5116 (
            .O(N__41504),
            .I(N__41498));
    LocalMux I__5115 (
            .O(N__41501),
            .I(\c0.n19030 ));
    LocalMux I__5114 (
            .O(N__41498),
            .I(\c0.n19030 ));
    InMux I__5113 (
            .O(N__41493),
            .I(N__41487));
    InMux I__5112 (
            .O(N__41492),
            .I(N__41480));
    InMux I__5111 (
            .O(N__41491),
            .I(N__41480));
    InMux I__5110 (
            .O(N__41490),
            .I(N__41480));
    LocalMux I__5109 (
            .O(N__41487),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__5108 (
            .O(N__41480),
            .I(\c0.data_in_frame_2_5 ));
    InMux I__5107 (
            .O(N__41475),
            .I(N__41472));
    LocalMux I__5106 (
            .O(N__41472),
            .I(\c0.n33386 ));
    CascadeMux I__5105 (
            .O(N__41469),
            .I(\c0.n33386_cascade_ ));
    InMux I__5104 (
            .O(N__41466),
            .I(N__41461));
    CascadeMux I__5103 (
            .O(N__41465),
            .I(N__41458));
    InMux I__5102 (
            .O(N__41464),
            .I(N__41455));
    LocalMux I__5101 (
            .O(N__41461),
            .I(N__41452));
    InMux I__5100 (
            .O(N__41458),
            .I(N__41448));
    LocalMux I__5099 (
            .O(N__41455),
            .I(N__41445));
    Span4Mux_h I__5098 (
            .O(N__41452),
            .I(N__41442));
    InMux I__5097 (
            .O(N__41451),
            .I(N__41439));
    LocalMux I__5096 (
            .O(N__41448),
            .I(\c0.data_in_frame_4_7 ));
    Odrv4 I__5095 (
            .O(N__41445),
            .I(\c0.data_in_frame_4_7 ));
    Odrv4 I__5094 (
            .O(N__41442),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__5093 (
            .O(N__41439),
            .I(\c0.data_in_frame_4_7 ));
    CascadeMux I__5092 (
            .O(N__41430),
            .I(N__41427));
    InMux I__5091 (
            .O(N__41427),
            .I(N__41421));
    InMux I__5090 (
            .O(N__41426),
            .I(N__41421));
    LocalMux I__5089 (
            .O(N__41421),
            .I(\c0.data_in_frame_3_0 ));
    CascadeMux I__5088 (
            .O(N__41418),
            .I(N__41414));
    InMux I__5087 (
            .O(N__41417),
            .I(N__41411));
    InMux I__5086 (
            .O(N__41414),
            .I(N__41407));
    LocalMux I__5085 (
            .O(N__41411),
            .I(N__41404));
    InMux I__5084 (
            .O(N__41410),
            .I(N__41401));
    LocalMux I__5083 (
            .O(N__41407),
            .I(\c0.data_in_frame_3_1 ));
    Odrv4 I__5082 (
            .O(N__41404),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__5081 (
            .O(N__41401),
            .I(\c0.data_in_frame_3_1 ));
    InMux I__5080 (
            .O(N__41394),
            .I(N__41391));
    LocalMux I__5079 (
            .O(N__41391),
            .I(N__41388));
    Span4Mux_h I__5078 (
            .O(N__41388),
            .I(N__41385));
    Odrv4 I__5077 (
            .O(N__41385),
            .I(\c0.n33473 ));
    InMux I__5076 (
            .O(N__41382),
            .I(N__41379));
    LocalMux I__5075 (
            .O(N__41379),
            .I(N__41376));
    Span4Mux_h I__5074 (
            .O(N__41376),
            .I(N__41372));
    InMux I__5073 (
            .O(N__41375),
            .I(N__41369));
    Odrv4 I__5072 (
            .O(N__41372),
            .I(\c0.n33451 ));
    LocalMux I__5071 (
            .O(N__41369),
            .I(\c0.n33451 ));
    CascadeMux I__5070 (
            .O(N__41364),
            .I(\c0.n6_adj_4503_cascade_ ));
    CascadeMux I__5069 (
            .O(N__41361),
            .I(N__41358));
    InMux I__5068 (
            .O(N__41358),
            .I(N__41353));
    InMux I__5067 (
            .O(N__41357),
            .I(N__41348));
    InMux I__5066 (
            .O(N__41356),
            .I(N__41348));
    LocalMux I__5065 (
            .O(N__41353),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__5064 (
            .O(N__41348),
            .I(\c0.data_in_frame_2_4 ));
    InMux I__5063 (
            .O(N__41343),
            .I(N__41339));
    InMux I__5062 (
            .O(N__41342),
            .I(N__41336));
    LocalMux I__5061 (
            .O(N__41339),
            .I(N__41332));
    LocalMux I__5060 (
            .O(N__41336),
            .I(N__41329));
    InMux I__5059 (
            .O(N__41335),
            .I(N__41326));
    Odrv4 I__5058 (
            .O(N__41332),
            .I(\quad_counter0.n3008 ));
    Odrv4 I__5057 (
            .O(N__41329),
            .I(\quad_counter0.n3008 ));
    LocalMux I__5056 (
            .O(N__41326),
            .I(\quad_counter0.n3008 ));
    InMux I__5055 (
            .O(N__41319),
            .I(\quad_counter0.n30340 ));
    InMux I__5054 (
            .O(N__41316),
            .I(N__41311));
    InMux I__5053 (
            .O(N__41315),
            .I(N__41308));
    CascadeMux I__5052 (
            .O(N__41314),
            .I(N__41305));
    LocalMux I__5051 (
            .O(N__41311),
            .I(N__41300));
    LocalMux I__5050 (
            .O(N__41308),
            .I(N__41300));
    InMux I__5049 (
            .O(N__41305),
            .I(N__41297));
    Odrv4 I__5048 (
            .O(N__41300),
            .I(\quad_counter0.n3007 ));
    LocalMux I__5047 (
            .O(N__41297),
            .I(\quad_counter0.n3007 ));
    InMux I__5046 (
            .O(N__41292),
            .I(\quad_counter0.n30341 ));
    InMux I__5045 (
            .O(N__41289),
            .I(N__41285));
    InMux I__5044 (
            .O(N__41288),
            .I(N__41282));
    LocalMux I__5043 (
            .O(N__41285),
            .I(N__41276));
    LocalMux I__5042 (
            .O(N__41282),
            .I(N__41276));
    InMux I__5041 (
            .O(N__41281),
            .I(N__41273));
    Odrv4 I__5040 (
            .O(N__41276),
            .I(\quad_counter0.n3006 ));
    LocalMux I__5039 (
            .O(N__41273),
            .I(\quad_counter0.n3006 ));
    InMux I__5038 (
            .O(N__41268),
            .I(\quad_counter0.n30342 ));
    InMux I__5037 (
            .O(N__41265),
            .I(N__41262));
    LocalMux I__5036 (
            .O(N__41262),
            .I(N__41257));
    InMux I__5035 (
            .O(N__41261),
            .I(N__41254));
    CascadeMux I__5034 (
            .O(N__41260),
            .I(N__41251));
    Span4Mux_h I__5033 (
            .O(N__41257),
            .I(N__41248));
    LocalMux I__5032 (
            .O(N__41254),
            .I(N__41245));
    InMux I__5031 (
            .O(N__41251),
            .I(N__41242));
    Odrv4 I__5030 (
            .O(N__41248),
            .I(\quad_counter0.n3005 ));
    Odrv4 I__5029 (
            .O(N__41245),
            .I(\quad_counter0.n3005 ));
    LocalMux I__5028 (
            .O(N__41242),
            .I(\quad_counter0.n3005 ));
    InMux I__5027 (
            .O(N__41235),
            .I(\quad_counter0.n30343 ));
    InMux I__5026 (
            .O(N__41232),
            .I(N__41229));
    LocalMux I__5025 (
            .O(N__41229),
            .I(N__41225));
    InMux I__5024 (
            .O(N__41228),
            .I(N__41221));
    Span4Mux_h I__5023 (
            .O(N__41225),
            .I(N__41218));
    InMux I__5022 (
            .O(N__41224),
            .I(N__41215));
    LocalMux I__5021 (
            .O(N__41221),
            .I(\quad_counter0.n3004 ));
    Odrv4 I__5020 (
            .O(N__41218),
            .I(\quad_counter0.n3004 ));
    LocalMux I__5019 (
            .O(N__41215),
            .I(\quad_counter0.n3004 ));
    InMux I__5018 (
            .O(N__41208),
            .I(\quad_counter0.n30344 ));
    InMux I__5017 (
            .O(N__41205),
            .I(N__41201));
    InMux I__5016 (
            .O(N__41204),
            .I(N__41198));
    LocalMux I__5015 (
            .O(N__41201),
            .I(N__41194));
    LocalMux I__5014 (
            .O(N__41198),
            .I(N__41191));
    InMux I__5013 (
            .O(N__41197),
            .I(N__41188));
    Odrv4 I__5012 (
            .O(N__41194),
            .I(\quad_counter0.n3003 ));
    Odrv4 I__5011 (
            .O(N__41191),
            .I(\quad_counter0.n3003 ));
    LocalMux I__5010 (
            .O(N__41188),
            .I(\quad_counter0.n3003 ));
    InMux I__5009 (
            .O(N__41181),
            .I(bfn_10_17_0_));
    InMux I__5008 (
            .O(N__41178),
            .I(\quad_counter0.n30346 ));
    InMux I__5007 (
            .O(N__41175),
            .I(N__41171));
    InMux I__5006 (
            .O(N__41174),
            .I(N__41168));
    LocalMux I__5005 (
            .O(N__41171),
            .I(N__41164));
    LocalMux I__5004 (
            .O(N__41168),
            .I(N__41161));
    InMux I__5003 (
            .O(N__41167),
            .I(N__41158));
    Odrv4 I__5002 (
            .O(N__41164),
            .I(\quad_counter0.n3002 ));
    Odrv4 I__5001 (
            .O(N__41161),
            .I(\quad_counter0.n3002 ));
    LocalMux I__5000 (
            .O(N__41158),
            .I(\quad_counter0.n3002 ));
    InMux I__4999 (
            .O(N__41151),
            .I(N__41146));
    InMux I__4998 (
            .O(N__41150),
            .I(N__41143));
    InMux I__4997 (
            .O(N__41149),
            .I(N__41139));
    LocalMux I__4996 (
            .O(N__41146),
            .I(N__41134));
    LocalMux I__4995 (
            .O(N__41143),
            .I(N__41134));
    InMux I__4994 (
            .O(N__41142),
            .I(N__41131));
    LocalMux I__4993 (
            .O(N__41139),
            .I(N__41128));
    Span4Mux_v I__4992 (
            .O(N__41134),
            .I(N__41125));
    LocalMux I__4991 (
            .O(N__41131),
            .I(data_in_2_5));
    Odrv12 I__4990 (
            .O(N__41128),
            .I(data_in_2_5));
    Odrv4 I__4989 (
            .O(N__41125),
            .I(data_in_2_5));
    InMux I__4988 (
            .O(N__41118),
            .I(N__41114));
    InMux I__4987 (
            .O(N__41117),
            .I(N__41111));
    LocalMux I__4986 (
            .O(N__41114),
            .I(N__41105));
    LocalMux I__4985 (
            .O(N__41111),
            .I(N__41105));
    CascadeMux I__4984 (
            .O(N__41110),
            .I(N__41102));
    Span4Mux_v I__4983 (
            .O(N__41105),
            .I(N__41099));
    InMux I__4982 (
            .O(N__41102),
            .I(N__41096));
    Odrv4 I__4981 (
            .O(N__41099),
            .I(\quad_counter0.n3016 ));
    LocalMux I__4980 (
            .O(N__41096),
            .I(\quad_counter0.n3016 ));
    InMux I__4979 (
            .O(N__41091),
            .I(\quad_counter0.n30332 ));
    InMux I__4978 (
            .O(N__41088),
            .I(N__41084));
    InMux I__4977 (
            .O(N__41087),
            .I(N__41081));
    LocalMux I__4976 (
            .O(N__41084),
            .I(N__41075));
    LocalMux I__4975 (
            .O(N__41081),
            .I(N__41075));
    InMux I__4974 (
            .O(N__41080),
            .I(N__41072));
    Odrv4 I__4973 (
            .O(N__41075),
            .I(\quad_counter0.n3015 ));
    LocalMux I__4972 (
            .O(N__41072),
            .I(\quad_counter0.n3015 ));
    InMux I__4971 (
            .O(N__41067),
            .I(\quad_counter0.n30333 ));
    InMux I__4970 (
            .O(N__41064),
            .I(\quad_counter0.n30334 ));
    InMux I__4969 (
            .O(N__41061),
            .I(N__41058));
    LocalMux I__4968 (
            .O(N__41058),
            .I(N__41054));
    InMux I__4967 (
            .O(N__41057),
            .I(N__41051));
    Span4Mux_h I__4966 (
            .O(N__41054),
            .I(N__41047));
    LocalMux I__4965 (
            .O(N__41051),
            .I(N__41044));
    InMux I__4964 (
            .O(N__41050),
            .I(N__41041));
    Odrv4 I__4963 (
            .O(N__41047),
            .I(\quad_counter0.n3013 ));
    Odrv4 I__4962 (
            .O(N__41044),
            .I(\quad_counter0.n3013 ));
    LocalMux I__4961 (
            .O(N__41041),
            .I(\quad_counter0.n3013 ));
    InMux I__4960 (
            .O(N__41034),
            .I(\quad_counter0.n30335 ));
    InMux I__4959 (
            .O(N__41031),
            .I(N__41026));
    InMux I__4958 (
            .O(N__41030),
            .I(N__41023));
    InMux I__4957 (
            .O(N__41029),
            .I(N__41020));
    LocalMux I__4956 (
            .O(N__41026),
            .I(\quad_counter0.n3012 ));
    LocalMux I__4955 (
            .O(N__41023),
            .I(\quad_counter0.n3012 ));
    LocalMux I__4954 (
            .O(N__41020),
            .I(\quad_counter0.n3012 ));
    InMux I__4953 (
            .O(N__41013),
            .I(\quad_counter0.n30336 ));
    InMux I__4952 (
            .O(N__41010),
            .I(N__41006));
    InMux I__4951 (
            .O(N__41009),
            .I(N__41003));
    LocalMux I__4950 (
            .O(N__41006),
            .I(N__40997));
    LocalMux I__4949 (
            .O(N__41003),
            .I(N__40997));
    InMux I__4948 (
            .O(N__41002),
            .I(N__40994));
    Odrv4 I__4947 (
            .O(N__40997),
            .I(\quad_counter0.n3011 ));
    LocalMux I__4946 (
            .O(N__40994),
            .I(\quad_counter0.n3011 ));
    InMux I__4945 (
            .O(N__40989),
            .I(bfn_10_16_0_));
    InMux I__4944 (
            .O(N__40986),
            .I(N__40982));
    InMux I__4943 (
            .O(N__40985),
            .I(N__40979));
    LocalMux I__4942 (
            .O(N__40982),
            .I(N__40975));
    LocalMux I__4941 (
            .O(N__40979),
            .I(N__40972));
    InMux I__4940 (
            .O(N__40978),
            .I(N__40969));
    Odrv4 I__4939 (
            .O(N__40975),
            .I(\quad_counter0.n3010 ));
    Odrv4 I__4938 (
            .O(N__40972),
            .I(\quad_counter0.n3010 ));
    LocalMux I__4937 (
            .O(N__40969),
            .I(\quad_counter0.n3010 ));
    InMux I__4936 (
            .O(N__40962),
            .I(\quad_counter0.n30338 ));
    InMux I__4935 (
            .O(N__40959),
            .I(N__40955));
    InMux I__4934 (
            .O(N__40958),
            .I(N__40952));
    LocalMux I__4933 (
            .O(N__40955),
            .I(N__40946));
    LocalMux I__4932 (
            .O(N__40952),
            .I(N__40946));
    InMux I__4931 (
            .O(N__40951),
            .I(N__40943));
    Odrv4 I__4930 (
            .O(N__40946),
            .I(\quad_counter0.n3009 ));
    LocalMux I__4929 (
            .O(N__40943),
            .I(\quad_counter0.n3009 ));
    InMux I__4928 (
            .O(N__40938),
            .I(\quad_counter0.n30339 ));
    InMux I__4927 (
            .O(N__40935),
            .I(N__40930));
    InMux I__4926 (
            .O(N__40934),
            .I(N__40927));
    InMux I__4925 (
            .O(N__40933),
            .I(N__40924));
    LocalMux I__4924 (
            .O(N__40930),
            .I(\quad_counter0.n3103 ));
    LocalMux I__4923 (
            .O(N__40927),
            .I(\quad_counter0.n3103 ));
    LocalMux I__4922 (
            .O(N__40924),
            .I(\quad_counter0.n3103 ));
    InMux I__4921 (
            .O(N__40917),
            .I(N__40912));
    InMux I__4920 (
            .O(N__40916),
            .I(N__40909));
    InMux I__4919 (
            .O(N__40915),
            .I(N__40906));
    LocalMux I__4918 (
            .O(N__40912),
            .I(N__40903));
    LocalMux I__4917 (
            .O(N__40909),
            .I(N__40898));
    LocalMux I__4916 (
            .O(N__40906),
            .I(N__40898));
    Span4Mux_h I__4915 (
            .O(N__40903),
            .I(N__40895));
    Odrv4 I__4914 (
            .O(N__40898),
            .I(\quad_counter0.n3202 ));
    Odrv4 I__4913 (
            .O(N__40895),
            .I(\quad_counter0.n3202 ));
    InMux I__4912 (
            .O(N__40890),
            .I(\quad_counter0.n30381 ));
    InMux I__4911 (
            .O(N__40887),
            .I(N__40882));
    InMux I__4910 (
            .O(N__40886),
            .I(N__40879));
    InMux I__4909 (
            .O(N__40885),
            .I(N__40876));
    LocalMux I__4908 (
            .O(N__40882),
            .I(N__40873));
    LocalMux I__4907 (
            .O(N__40879),
            .I(\quad_counter0.n3102 ));
    LocalMux I__4906 (
            .O(N__40876),
            .I(\quad_counter0.n3102 ));
    Odrv4 I__4905 (
            .O(N__40873),
            .I(\quad_counter0.n3102 ));
    InMux I__4904 (
            .O(N__40866),
            .I(N__40861));
    InMux I__4903 (
            .O(N__40865),
            .I(N__40856));
    InMux I__4902 (
            .O(N__40864),
            .I(N__40856));
    LocalMux I__4901 (
            .O(N__40861),
            .I(N__40851));
    LocalMux I__4900 (
            .O(N__40856),
            .I(N__40851));
    Odrv4 I__4899 (
            .O(N__40851),
            .I(\quad_counter0.n3201 ));
    InMux I__4898 (
            .O(N__40848),
            .I(\quad_counter0.n30382 ));
    InMux I__4897 (
            .O(N__40845),
            .I(N__40840));
    InMux I__4896 (
            .O(N__40844),
            .I(N__40837));
    InMux I__4895 (
            .O(N__40843),
            .I(N__40834));
    LocalMux I__4894 (
            .O(N__40840),
            .I(N__40831));
    LocalMux I__4893 (
            .O(N__40837),
            .I(\quad_counter0.n3101 ));
    LocalMux I__4892 (
            .O(N__40834),
            .I(\quad_counter0.n3101 ));
    Odrv4 I__4891 (
            .O(N__40831),
            .I(\quad_counter0.n3101 ));
    CascadeMux I__4890 (
            .O(N__40824),
            .I(N__40818));
    CascadeMux I__4889 (
            .O(N__40823),
            .I(N__40815));
    CascadeMux I__4888 (
            .O(N__40822),
            .I(N__40812));
    CascadeMux I__4887 (
            .O(N__40821),
            .I(N__40809));
    InMux I__4886 (
            .O(N__40818),
            .I(N__40794));
    InMux I__4885 (
            .O(N__40815),
            .I(N__40794));
    InMux I__4884 (
            .O(N__40812),
            .I(N__40789));
    InMux I__4883 (
            .O(N__40809),
            .I(N__40789));
    CascadeMux I__4882 (
            .O(N__40808),
            .I(N__40786));
    CascadeMux I__4881 (
            .O(N__40807),
            .I(N__40783));
    CascadeMux I__4880 (
            .O(N__40806),
            .I(N__40780));
    CascadeMux I__4879 (
            .O(N__40805),
            .I(N__40777));
    CascadeMux I__4878 (
            .O(N__40804),
            .I(N__40774));
    CascadeMux I__4877 (
            .O(N__40803),
            .I(N__40771));
    CascadeMux I__4876 (
            .O(N__40802),
            .I(N__40768));
    CascadeMux I__4875 (
            .O(N__40801),
            .I(N__40765));
    CascadeMux I__4874 (
            .O(N__40800),
            .I(N__40762));
    CascadeMux I__4873 (
            .O(N__40799),
            .I(N__40759));
    LocalMux I__4872 (
            .O(N__40794),
            .I(N__40753));
    LocalMux I__4871 (
            .O(N__40789),
            .I(N__40753));
    InMux I__4870 (
            .O(N__40786),
            .I(N__40744));
    InMux I__4869 (
            .O(N__40783),
            .I(N__40744));
    InMux I__4868 (
            .O(N__40780),
            .I(N__40744));
    InMux I__4867 (
            .O(N__40777),
            .I(N__40744));
    InMux I__4866 (
            .O(N__40774),
            .I(N__40735));
    InMux I__4865 (
            .O(N__40771),
            .I(N__40735));
    InMux I__4864 (
            .O(N__40768),
            .I(N__40735));
    InMux I__4863 (
            .O(N__40765),
            .I(N__40735));
    InMux I__4862 (
            .O(N__40762),
            .I(N__40730));
    InMux I__4861 (
            .O(N__40759),
            .I(N__40730));
    InMux I__4860 (
            .O(N__40758),
            .I(N__40727));
    Odrv4 I__4859 (
            .O(N__40753),
            .I(\quad_counter0.n3134 ));
    LocalMux I__4858 (
            .O(N__40744),
            .I(\quad_counter0.n3134 ));
    LocalMux I__4857 (
            .O(N__40735),
            .I(\quad_counter0.n3134 ));
    LocalMux I__4856 (
            .O(N__40730),
            .I(\quad_counter0.n3134 ));
    LocalMux I__4855 (
            .O(N__40727),
            .I(\quad_counter0.n3134 ));
    InMux I__4854 (
            .O(N__40716),
            .I(\quad_counter0.n30383 ));
    CascadeMux I__4853 (
            .O(N__40713),
            .I(N__40708));
    InMux I__4852 (
            .O(N__40712),
            .I(N__40705));
    InMux I__4851 (
            .O(N__40711),
            .I(N__40702));
    InMux I__4850 (
            .O(N__40708),
            .I(N__40699));
    LocalMux I__4849 (
            .O(N__40705),
            .I(N__40692));
    LocalMux I__4848 (
            .O(N__40702),
            .I(N__40692));
    LocalMux I__4847 (
            .O(N__40699),
            .I(N__40692));
    Odrv4 I__4846 (
            .O(N__40692),
            .I(\quad_counter0.n3200 ));
    InMux I__4845 (
            .O(N__40689),
            .I(N__40686));
    LocalMux I__4844 (
            .O(N__40686),
            .I(N__40683));
    Span4Mux_h I__4843 (
            .O(N__40683),
            .I(N__40680));
    Odrv4 I__4842 (
            .O(N__40680),
            .I(\c0.n93_adj_4634 ));
    InMux I__4841 (
            .O(N__40677),
            .I(bfn_10_15_0_));
    InMux I__4840 (
            .O(N__40674),
            .I(\quad_counter0.n30330 ));
    InMux I__4839 (
            .O(N__40671),
            .I(\quad_counter0.n30331 ));
    InMux I__4838 (
            .O(N__40668),
            .I(N__40663));
    InMux I__4837 (
            .O(N__40667),
            .I(N__40660));
    InMux I__4836 (
            .O(N__40666),
            .I(N__40657));
    LocalMux I__4835 (
            .O(N__40663),
            .I(N__40654));
    LocalMux I__4834 (
            .O(N__40660),
            .I(\quad_counter0.n3111 ));
    LocalMux I__4833 (
            .O(N__40657),
            .I(\quad_counter0.n3111 ));
    Odrv4 I__4832 (
            .O(N__40654),
            .I(\quad_counter0.n3111 ));
    InMux I__4831 (
            .O(N__40647),
            .I(N__40643));
    InMux I__4830 (
            .O(N__40646),
            .I(N__40640));
    LocalMux I__4829 (
            .O(N__40643),
            .I(N__40634));
    LocalMux I__4828 (
            .O(N__40640),
            .I(N__40634));
    InMux I__4827 (
            .O(N__40639),
            .I(N__40631));
    Span4Mux_h I__4826 (
            .O(N__40634),
            .I(N__40626));
    LocalMux I__4825 (
            .O(N__40631),
            .I(N__40626));
    Odrv4 I__4824 (
            .O(N__40626),
            .I(\quad_counter0.n3210 ));
    InMux I__4823 (
            .O(N__40623),
            .I(\quad_counter0.n30373 ));
    InMux I__4822 (
            .O(N__40620),
            .I(N__40615));
    InMux I__4821 (
            .O(N__40619),
            .I(N__40612));
    InMux I__4820 (
            .O(N__40618),
            .I(N__40609));
    LocalMux I__4819 (
            .O(N__40615),
            .I(N__40606));
    LocalMux I__4818 (
            .O(N__40612),
            .I(\quad_counter0.n3110 ));
    LocalMux I__4817 (
            .O(N__40609),
            .I(\quad_counter0.n3110 ));
    Odrv4 I__4816 (
            .O(N__40606),
            .I(\quad_counter0.n3110 ));
    InMux I__4815 (
            .O(N__40599),
            .I(N__40594));
    InMux I__4814 (
            .O(N__40598),
            .I(N__40591));
    InMux I__4813 (
            .O(N__40597),
            .I(N__40588));
    LocalMux I__4812 (
            .O(N__40594),
            .I(N__40581));
    LocalMux I__4811 (
            .O(N__40591),
            .I(N__40581));
    LocalMux I__4810 (
            .O(N__40588),
            .I(N__40581));
    Odrv4 I__4809 (
            .O(N__40581),
            .I(\quad_counter0.n3209 ));
    InMux I__4808 (
            .O(N__40578),
            .I(\quad_counter0.n30374 ));
    InMux I__4807 (
            .O(N__40575),
            .I(N__40570));
    InMux I__4806 (
            .O(N__40574),
            .I(N__40567));
    InMux I__4805 (
            .O(N__40573),
            .I(N__40564));
    LocalMux I__4804 (
            .O(N__40570),
            .I(N__40561));
    LocalMux I__4803 (
            .O(N__40567),
            .I(\quad_counter0.n3109 ));
    LocalMux I__4802 (
            .O(N__40564),
            .I(\quad_counter0.n3109 ));
    Odrv4 I__4801 (
            .O(N__40561),
            .I(\quad_counter0.n3109 ));
    InMux I__4800 (
            .O(N__40554),
            .I(N__40549));
    InMux I__4799 (
            .O(N__40553),
            .I(N__40546));
    InMux I__4798 (
            .O(N__40552),
            .I(N__40543));
    LocalMux I__4797 (
            .O(N__40549),
            .I(N__40538));
    LocalMux I__4796 (
            .O(N__40546),
            .I(N__40538));
    LocalMux I__4795 (
            .O(N__40543),
            .I(N__40535));
    Odrv4 I__4794 (
            .O(N__40538),
            .I(\quad_counter0.n3208 ));
    Odrv4 I__4793 (
            .O(N__40535),
            .I(\quad_counter0.n3208 ));
    InMux I__4792 (
            .O(N__40530),
            .I(\quad_counter0.n30375 ));
    InMux I__4791 (
            .O(N__40527),
            .I(N__40522));
    InMux I__4790 (
            .O(N__40526),
            .I(N__40519));
    InMux I__4789 (
            .O(N__40525),
            .I(N__40516));
    LocalMux I__4788 (
            .O(N__40522),
            .I(\quad_counter0.n3108 ));
    LocalMux I__4787 (
            .O(N__40519),
            .I(\quad_counter0.n3108 ));
    LocalMux I__4786 (
            .O(N__40516),
            .I(\quad_counter0.n3108 ));
    CascadeMux I__4785 (
            .O(N__40509),
            .I(N__40504));
    InMux I__4784 (
            .O(N__40508),
            .I(N__40501));
    InMux I__4783 (
            .O(N__40507),
            .I(N__40498));
    InMux I__4782 (
            .O(N__40504),
            .I(N__40495));
    LocalMux I__4781 (
            .O(N__40501),
            .I(N__40488));
    LocalMux I__4780 (
            .O(N__40498),
            .I(N__40488));
    LocalMux I__4779 (
            .O(N__40495),
            .I(N__40488));
    Odrv4 I__4778 (
            .O(N__40488),
            .I(\quad_counter0.n3207 ));
    InMux I__4777 (
            .O(N__40485),
            .I(\quad_counter0.n30376 ));
    CascadeMux I__4776 (
            .O(N__40482),
            .I(N__40477));
    InMux I__4775 (
            .O(N__40481),
            .I(N__40474));
    InMux I__4774 (
            .O(N__40480),
            .I(N__40471));
    InMux I__4773 (
            .O(N__40477),
            .I(N__40468));
    LocalMux I__4772 (
            .O(N__40474),
            .I(\quad_counter0.n3107 ));
    LocalMux I__4771 (
            .O(N__40471),
            .I(\quad_counter0.n3107 ));
    LocalMux I__4770 (
            .O(N__40468),
            .I(\quad_counter0.n3107 ));
    InMux I__4769 (
            .O(N__40461),
            .I(N__40456));
    InMux I__4768 (
            .O(N__40460),
            .I(N__40453));
    InMux I__4767 (
            .O(N__40459),
            .I(N__40450));
    LocalMux I__4766 (
            .O(N__40456),
            .I(N__40447));
    LocalMux I__4765 (
            .O(N__40453),
            .I(N__40440));
    LocalMux I__4764 (
            .O(N__40450),
            .I(N__40440));
    Span4Mux_h I__4763 (
            .O(N__40447),
            .I(N__40440));
    Odrv4 I__4762 (
            .O(N__40440),
            .I(\quad_counter0.n3206 ));
    InMux I__4761 (
            .O(N__40437),
            .I(\quad_counter0.n30377 ));
    InMux I__4760 (
            .O(N__40434),
            .I(N__40430));
    InMux I__4759 (
            .O(N__40433),
            .I(N__40427));
    LocalMux I__4758 (
            .O(N__40430),
            .I(N__40421));
    LocalMux I__4757 (
            .O(N__40427),
            .I(N__40421));
    InMux I__4756 (
            .O(N__40426),
            .I(N__40418));
    Odrv4 I__4755 (
            .O(N__40421),
            .I(\quad_counter0.n3106 ));
    LocalMux I__4754 (
            .O(N__40418),
            .I(\quad_counter0.n3106 ));
    InMux I__4753 (
            .O(N__40413),
            .I(N__40409));
    InMux I__4752 (
            .O(N__40412),
            .I(N__40406));
    LocalMux I__4751 (
            .O(N__40409),
            .I(N__40400));
    LocalMux I__4750 (
            .O(N__40406),
            .I(N__40400));
    InMux I__4749 (
            .O(N__40405),
            .I(N__40397));
    Span4Mux_h I__4748 (
            .O(N__40400),
            .I(N__40392));
    LocalMux I__4747 (
            .O(N__40397),
            .I(N__40392));
    Odrv4 I__4746 (
            .O(N__40392),
            .I(\quad_counter0.n3205 ));
    InMux I__4745 (
            .O(N__40389),
            .I(\quad_counter0.n30378 ));
    InMux I__4744 (
            .O(N__40386),
            .I(N__40381));
    InMux I__4743 (
            .O(N__40385),
            .I(N__40378));
    InMux I__4742 (
            .O(N__40384),
            .I(N__40375));
    LocalMux I__4741 (
            .O(N__40381),
            .I(N__40372));
    LocalMux I__4740 (
            .O(N__40378),
            .I(\quad_counter0.n3105 ));
    LocalMux I__4739 (
            .O(N__40375),
            .I(\quad_counter0.n3105 ));
    Odrv4 I__4738 (
            .O(N__40372),
            .I(\quad_counter0.n3105 ));
    InMux I__4737 (
            .O(N__40365),
            .I(N__40360));
    InMux I__4736 (
            .O(N__40364),
            .I(N__40355));
    InMux I__4735 (
            .O(N__40363),
            .I(N__40355));
    LocalMux I__4734 (
            .O(N__40360),
            .I(N__40350));
    LocalMux I__4733 (
            .O(N__40355),
            .I(N__40350));
    Odrv4 I__4732 (
            .O(N__40350),
            .I(\quad_counter0.n3204 ));
    InMux I__4731 (
            .O(N__40347),
            .I(\quad_counter0.n30379 ));
    InMux I__4730 (
            .O(N__40344),
            .I(N__40339));
    InMux I__4729 (
            .O(N__40343),
            .I(N__40336));
    InMux I__4728 (
            .O(N__40342),
            .I(N__40333));
    LocalMux I__4727 (
            .O(N__40339),
            .I(N__40330));
    LocalMux I__4726 (
            .O(N__40336),
            .I(\quad_counter0.n3104 ));
    LocalMux I__4725 (
            .O(N__40333),
            .I(\quad_counter0.n3104 ));
    Odrv4 I__4724 (
            .O(N__40330),
            .I(\quad_counter0.n3104 ));
    InMux I__4723 (
            .O(N__40323),
            .I(N__40318));
    InMux I__4722 (
            .O(N__40322),
            .I(N__40313));
    InMux I__4721 (
            .O(N__40321),
            .I(N__40313));
    LocalMux I__4720 (
            .O(N__40318),
            .I(N__40308));
    LocalMux I__4719 (
            .O(N__40313),
            .I(N__40308));
    Odrv4 I__4718 (
            .O(N__40308),
            .I(\quad_counter0.n3203 ));
    InMux I__4717 (
            .O(N__40305),
            .I(bfn_10_14_0_));
    InMux I__4716 (
            .O(N__40302),
            .I(N__40297));
    InMux I__4715 (
            .O(N__40301),
            .I(N__40294));
    InMux I__4714 (
            .O(N__40300),
            .I(N__40291));
    LocalMux I__4713 (
            .O(N__40297),
            .I(\quad_counter0.n3119 ));
    LocalMux I__4712 (
            .O(N__40294),
            .I(\quad_counter0.n3119 ));
    LocalMux I__4711 (
            .O(N__40291),
            .I(\quad_counter0.n3119 ));
    InMux I__4710 (
            .O(N__40284),
            .I(\quad_counter0.n30365 ));
    CascadeMux I__4709 (
            .O(N__40281),
            .I(N__40276));
    InMux I__4708 (
            .O(N__40280),
            .I(N__40273));
    InMux I__4707 (
            .O(N__40279),
            .I(N__40270));
    InMux I__4706 (
            .O(N__40276),
            .I(N__40267));
    LocalMux I__4705 (
            .O(N__40273),
            .I(\quad_counter0.n3118 ));
    LocalMux I__4704 (
            .O(N__40270),
            .I(\quad_counter0.n3118 ));
    LocalMux I__4703 (
            .O(N__40267),
            .I(\quad_counter0.n3118 ));
    InMux I__4702 (
            .O(N__40260),
            .I(\quad_counter0.n30366 ));
    InMux I__4701 (
            .O(N__40257),
            .I(N__40252));
    InMux I__4700 (
            .O(N__40256),
            .I(N__40249));
    InMux I__4699 (
            .O(N__40255),
            .I(N__40246));
    LocalMux I__4698 (
            .O(N__40252),
            .I(N__40243));
    LocalMux I__4697 (
            .O(N__40249),
            .I(N__40240));
    LocalMux I__4696 (
            .O(N__40246),
            .I(N__40237));
    Span4Mux_h I__4695 (
            .O(N__40243),
            .I(N__40234));
    Odrv4 I__4694 (
            .O(N__40240),
            .I(\quad_counter0.n3216 ));
    Odrv4 I__4693 (
            .O(N__40237),
            .I(\quad_counter0.n3216 ));
    Odrv4 I__4692 (
            .O(N__40234),
            .I(\quad_counter0.n3216 ));
    InMux I__4691 (
            .O(N__40227),
            .I(\quad_counter0.n30367 ));
    InMux I__4690 (
            .O(N__40224),
            .I(N__40220));
    InMux I__4689 (
            .O(N__40223),
            .I(N__40217));
    LocalMux I__4688 (
            .O(N__40220),
            .I(N__40211));
    LocalMux I__4687 (
            .O(N__40217),
            .I(N__40211));
    InMux I__4686 (
            .O(N__40216),
            .I(N__40208));
    Odrv4 I__4685 (
            .O(N__40211),
            .I(\quad_counter0.n3116 ));
    LocalMux I__4684 (
            .O(N__40208),
            .I(\quad_counter0.n3116 ));
    InMux I__4683 (
            .O(N__40203),
            .I(N__40198));
    InMux I__4682 (
            .O(N__40202),
            .I(N__40195));
    InMux I__4681 (
            .O(N__40201),
            .I(N__40192));
    LocalMux I__4680 (
            .O(N__40198),
            .I(N__40189));
    LocalMux I__4679 (
            .O(N__40195),
            .I(N__40184));
    LocalMux I__4678 (
            .O(N__40192),
            .I(N__40184));
    Odrv4 I__4677 (
            .O(N__40189),
            .I(\quad_counter0.n3215 ));
    Odrv4 I__4676 (
            .O(N__40184),
            .I(\quad_counter0.n3215 ));
    InMux I__4675 (
            .O(N__40179),
            .I(\quad_counter0.n30368 ));
    InMux I__4674 (
            .O(N__40176),
            .I(N__40171));
    InMux I__4673 (
            .O(N__40175),
            .I(N__40168));
    InMux I__4672 (
            .O(N__40174),
            .I(N__40165));
    LocalMux I__4671 (
            .O(N__40171),
            .I(\quad_counter0.n3115 ));
    LocalMux I__4670 (
            .O(N__40168),
            .I(\quad_counter0.n3115 ));
    LocalMux I__4669 (
            .O(N__40165),
            .I(\quad_counter0.n3115 ));
    InMux I__4668 (
            .O(N__40158),
            .I(\quad_counter0.n30369 ));
    CascadeMux I__4667 (
            .O(N__40155),
            .I(N__40147));
    CascadeMux I__4666 (
            .O(N__40154),
            .I(N__40144));
    CascadeMux I__4665 (
            .O(N__40153),
            .I(N__40141));
    CascadeMux I__4664 (
            .O(N__40152),
            .I(N__40138));
    CascadeMux I__4663 (
            .O(N__40151),
            .I(N__40135));
    CascadeMux I__4662 (
            .O(N__40150),
            .I(N__40132));
    InMux I__4661 (
            .O(N__40147),
            .I(N__40127));
    InMux I__4660 (
            .O(N__40144),
            .I(N__40127));
    InMux I__4659 (
            .O(N__40141),
            .I(N__40118));
    InMux I__4658 (
            .O(N__40138),
            .I(N__40118));
    InMux I__4657 (
            .O(N__40135),
            .I(N__40118));
    InMux I__4656 (
            .O(N__40132),
            .I(N__40118));
    LocalMux I__4655 (
            .O(N__40127),
            .I(\quad_counter0.n36143 ));
    LocalMux I__4654 (
            .O(N__40118),
            .I(\quad_counter0.n36143 ));
    InMux I__4653 (
            .O(N__40113),
            .I(N__40109));
    InMux I__4652 (
            .O(N__40112),
            .I(N__40106));
    LocalMux I__4651 (
            .O(N__40109),
            .I(N__40100));
    LocalMux I__4650 (
            .O(N__40106),
            .I(N__40100));
    InMux I__4649 (
            .O(N__40105),
            .I(N__40097));
    Span4Mux_v I__4648 (
            .O(N__40100),
            .I(N__40094));
    LocalMux I__4647 (
            .O(N__40097),
            .I(N__40091));
    Odrv4 I__4646 (
            .O(N__40094),
            .I(\quad_counter0.n3213 ));
    Odrv4 I__4645 (
            .O(N__40091),
            .I(\quad_counter0.n3213 ));
    InMux I__4644 (
            .O(N__40086),
            .I(\quad_counter0.n30370 ));
    InMux I__4643 (
            .O(N__40083),
            .I(N__40078));
    InMux I__4642 (
            .O(N__40082),
            .I(N__40075));
    InMux I__4641 (
            .O(N__40081),
            .I(N__40072));
    LocalMux I__4640 (
            .O(N__40078),
            .I(\quad_counter0.n3113 ));
    LocalMux I__4639 (
            .O(N__40075),
            .I(\quad_counter0.n3113 ));
    LocalMux I__4638 (
            .O(N__40072),
            .I(\quad_counter0.n3113 ));
    InMux I__4637 (
            .O(N__40065),
            .I(N__40060));
    InMux I__4636 (
            .O(N__40064),
            .I(N__40057));
    CascadeMux I__4635 (
            .O(N__40063),
            .I(N__40054));
    LocalMux I__4634 (
            .O(N__40060),
            .I(N__40049));
    LocalMux I__4633 (
            .O(N__40057),
            .I(N__40049));
    InMux I__4632 (
            .O(N__40054),
            .I(N__40046));
    Odrv4 I__4631 (
            .O(N__40049),
            .I(\quad_counter0.n3212 ));
    LocalMux I__4630 (
            .O(N__40046),
            .I(\quad_counter0.n3212 ));
    InMux I__4629 (
            .O(N__40041),
            .I(\quad_counter0.n30371 ));
    InMux I__4628 (
            .O(N__40038),
            .I(N__40033));
    InMux I__4627 (
            .O(N__40037),
            .I(N__40030));
    InMux I__4626 (
            .O(N__40036),
            .I(N__40027));
    LocalMux I__4625 (
            .O(N__40033),
            .I(\quad_counter0.n3112 ));
    LocalMux I__4624 (
            .O(N__40030),
            .I(\quad_counter0.n3112 ));
    LocalMux I__4623 (
            .O(N__40027),
            .I(\quad_counter0.n3112 ));
    InMux I__4622 (
            .O(N__40020),
            .I(N__40016));
    InMux I__4621 (
            .O(N__40019),
            .I(N__40012));
    LocalMux I__4620 (
            .O(N__40016),
            .I(N__40009));
    InMux I__4619 (
            .O(N__40015),
            .I(N__40006));
    LocalMux I__4618 (
            .O(N__40012),
            .I(N__40003));
    Span4Mux_h I__4617 (
            .O(N__40009),
            .I(N__39998));
    LocalMux I__4616 (
            .O(N__40006),
            .I(N__39998));
    Odrv4 I__4615 (
            .O(N__40003),
            .I(\quad_counter0.n3211 ));
    Odrv4 I__4614 (
            .O(N__39998),
            .I(\quad_counter0.n3211 ));
    InMux I__4613 (
            .O(N__39993),
            .I(bfn_10_13_0_));
    InMux I__4612 (
            .O(N__39990),
            .I(bfn_10_11_0_));
    InMux I__4611 (
            .O(N__39987),
            .I(\quad_counter0.n30400 ));
    InMux I__4610 (
            .O(N__39984),
            .I(\quad_counter0.n30401 ));
    InMux I__4609 (
            .O(N__39981),
            .I(\quad_counter0.n30402 ));
    InMux I__4608 (
            .O(N__39978),
            .I(\quad_counter0.n30403 ));
    CascadeMux I__4607 (
            .O(N__39975),
            .I(N__39961));
    CascadeMux I__4606 (
            .O(N__39974),
            .I(N__39958));
    CascadeMux I__4605 (
            .O(N__39973),
            .I(N__39952));
    CascadeMux I__4604 (
            .O(N__39972),
            .I(N__39949));
    CascadeMux I__4603 (
            .O(N__39971),
            .I(N__39946));
    CascadeMux I__4602 (
            .O(N__39970),
            .I(N__39943));
    CascadeMux I__4601 (
            .O(N__39969),
            .I(N__39940));
    CascadeMux I__4600 (
            .O(N__39968),
            .I(N__39937));
    CascadeMux I__4599 (
            .O(N__39967),
            .I(N__39934));
    CascadeMux I__4598 (
            .O(N__39966),
            .I(N__39931));
    CascadeMux I__4597 (
            .O(N__39965),
            .I(N__39928));
    CascadeMux I__4596 (
            .O(N__39964),
            .I(N__39925));
    InMux I__4595 (
            .O(N__39961),
            .I(N__39920));
    InMux I__4594 (
            .O(N__39958),
            .I(N__39920));
    CascadeMux I__4593 (
            .O(N__39957),
            .I(N__39917));
    CascadeMux I__4592 (
            .O(N__39956),
            .I(N__39914));
    CascadeMux I__4591 (
            .O(N__39955),
            .I(N__39911));
    InMux I__4590 (
            .O(N__39952),
            .I(N__39905));
    InMux I__4589 (
            .O(N__39949),
            .I(N__39905));
    InMux I__4588 (
            .O(N__39946),
            .I(N__39896));
    InMux I__4587 (
            .O(N__39943),
            .I(N__39896));
    InMux I__4586 (
            .O(N__39940),
            .I(N__39896));
    InMux I__4585 (
            .O(N__39937),
            .I(N__39896));
    InMux I__4584 (
            .O(N__39934),
            .I(N__39887));
    InMux I__4583 (
            .O(N__39931),
            .I(N__39887));
    InMux I__4582 (
            .O(N__39928),
            .I(N__39887));
    InMux I__4581 (
            .O(N__39925),
            .I(N__39887));
    LocalMux I__4580 (
            .O(N__39920),
            .I(N__39884));
    InMux I__4579 (
            .O(N__39917),
            .I(N__39875));
    InMux I__4578 (
            .O(N__39914),
            .I(N__39875));
    InMux I__4577 (
            .O(N__39911),
            .I(N__39875));
    InMux I__4576 (
            .O(N__39910),
            .I(N__39875));
    LocalMux I__4575 (
            .O(N__39905),
            .I(\quad_counter0.n3233 ));
    LocalMux I__4574 (
            .O(N__39896),
            .I(\quad_counter0.n3233 ));
    LocalMux I__4573 (
            .O(N__39887),
            .I(\quad_counter0.n3233 ));
    Odrv4 I__4572 (
            .O(N__39884),
            .I(\quad_counter0.n3233 ));
    LocalMux I__4571 (
            .O(N__39875),
            .I(\quad_counter0.n3233 ));
    CascadeMux I__4570 (
            .O(N__39864),
            .I(N__39856));
    CascadeMux I__4569 (
            .O(N__39863),
            .I(N__39853));
    CascadeMux I__4568 (
            .O(N__39862),
            .I(N__39850));
    CascadeMux I__4567 (
            .O(N__39861),
            .I(N__39847));
    CascadeMux I__4566 (
            .O(N__39860),
            .I(N__39844));
    CascadeMux I__4565 (
            .O(N__39859),
            .I(N__39841));
    InMux I__4564 (
            .O(N__39856),
            .I(N__39836));
    InMux I__4563 (
            .O(N__39853),
            .I(N__39836));
    InMux I__4562 (
            .O(N__39850),
            .I(N__39827));
    InMux I__4561 (
            .O(N__39847),
            .I(N__39827));
    InMux I__4560 (
            .O(N__39844),
            .I(N__39827));
    InMux I__4559 (
            .O(N__39841),
            .I(N__39827));
    LocalMux I__4558 (
            .O(N__39836),
            .I(N__39824));
    LocalMux I__4557 (
            .O(N__39827),
            .I(N__39821));
    Odrv4 I__4556 (
            .O(N__39824),
            .I(\quad_counter0.n36141 ));
    Odrv4 I__4555 (
            .O(N__39821),
            .I(\quad_counter0.n36141 ));
    CascadeMux I__4554 (
            .O(N__39816),
            .I(N__39813));
    InMux I__4553 (
            .O(N__39813),
            .I(N__39810));
    LocalMux I__4552 (
            .O(N__39810),
            .I(\quad_counter0.n26_adj_4358 ));
    InMux I__4551 (
            .O(N__39807),
            .I(N__39804));
    LocalMux I__4550 (
            .O(N__39804),
            .I(\quad_counter0.n16_adj_4359 ));
    InMux I__4549 (
            .O(N__39801),
            .I(bfn_10_12_0_));
    InMux I__4548 (
            .O(N__39798),
            .I(\quad_counter0.n30390 ));
    InMux I__4547 (
            .O(N__39795),
            .I(bfn_10_10_0_));
    InMux I__4546 (
            .O(N__39792),
            .I(\quad_counter0.n30392 ));
    InMux I__4545 (
            .O(N__39789),
            .I(\quad_counter0.n30393 ));
    InMux I__4544 (
            .O(N__39786),
            .I(\quad_counter0.n30394 ));
    InMux I__4543 (
            .O(N__39783),
            .I(\quad_counter0.n30395 ));
    InMux I__4542 (
            .O(N__39780),
            .I(\quad_counter0.n30396 ));
    InMux I__4541 (
            .O(N__39777),
            .I(\quad_counter0.n30397 ));
    InMux I__4540 (
            .O(N__39774),
            .I(\quad_counter0.n30398 ));
    CascadeMux I__4539 (
            .O(N__39771),
            .I(n17985_cascade_));
    CEMux I__4538 (
            .O(N__39768),
            .I(N__39763));
    CEMux I__4537 (
            .O(N__39767),
            .I(N__39760));
    InMux I__4536 (
            .O(N__39766),
            .I(N__39757));
    LocalMux I__4535 (
            .O(N__39763),
            .I(n19433));
    LocalMux I__4534 (
            .O(N__39760),
            .I(n19433));
    LocalMux I__4533 (
            .O(N__39757),
            .I(n19433));
    InMux I__4532 (
            .O(N__39750),
            .I(N__39746));
    InMux I__4531 (
            .O(N__39749),
            .I(N__39743));
    LocalMux I__4530 (
            .O(N__39746),
            .I(\quad_counter1.a_delay_counter_11 ));
    LocalMux I__4529 (
            .O(N__39743),
            .I(\quad_counter1.a_delay_counter_11 ));
    InMux I__4528 (
            .O(N__39738),
            .I(N__39734));
    InMux I__4527 (
            .O(N__39737),
            .I(N__39731));
    LocalMux I__4526 (
            .O(N__39734),
            .I(\quad_counter1.a_delay_counter_6 ));
    LocalMux I__4525 (
            .O(N__39731),
            .I(\quad_counter1.a_delay_counter_6 ));
    CascadeMux I__4524 (
            .O(N__39726),
            .I(N__39723));
    InMux I__4523 (
            .O(N__39723),
            .I(N__39719));
    InMux I__4522 (
            .O(N__39722),
            .I(N__39716));
    LocalMux I__4521 (
            .O(N__39719),
            .I(N__39713));
    LocalMux I__4520 (
            .O(N__39716),
            .I(\quad_counter1.a_delay_counter_10 ));
    Odrv4 I__4519 (
            .O(N__39713),
            .I(\quad_counter1.a_delay_counter_10 ));
    InMux I__4518 (
            .O(N__39708),
            .I(N__39704));
    InMux I__4517 (
            .O(N__39707),
            .I(N__39701));
    LocalMux I__4516 (
            .O(N__39704),
            .I(\quad_counter1.a_delay_counter_8 ));
    LocalMux I__4515 (
            .O(N__39701),
            .I(\quad_counter1.a_delay_counter_8 ));
    InMux I__4514 (
            .O(N__39696),
            .I(N__39693));
    LocalMux I__4513 (
            .O(N__39693),
            .I(\quad_counter1.n26_adj_4441 ));
    InMux I__4512 (
            .O(N__39690),
            .I(bfn_10_9_0_));
    InMux I__4511 (
            .O(N__39687),
            .I(\quad_counter0.n30384 ));
    InMux I__4510 (
            .O(N__39684),
            .I(\quad_counter0.n30385 ));
    InMux I__4509 (
            .O(N__39681),
            .I(\quad_counter0.n30386 ));
    InMux I__4508 (
            .O(N__39678),
            .I(\quad_counter0.n30387 ));
    InMux I__4507 (
            .O(N__39675),
            .I(\quad_counter0.n30388 ));
    InMux I__4506 (
            .O(N__39672),
            .I(\quad_counter0.n30389 ));
    SRMux I__4505 (
            .O(N__39669),
            .I(N__39665));
    SRMux I__4504 (
            .O(N__39668),
            .I(N__39662));
    LocalMux I__4503 (
            .O(N__39665),
            .I(N__39658));
    LocalMux I__4502 (
            .O(N__39662),
            .I(N__39655));
    InMux I__4501 (
            .O(N__39661),
            .I(N__39652));
    Span4Mux_v I__4500 (
            .O(N__39658),
            .I(N__39645));
    Span4Mux_h I__4499 (
            .O(N__39655),
            .I(N__39645));
    LocalMux I__4498 (
            .O(N__39652),
            .I(N__39645));
    Odrv4 I__4497 (
            .O(N__39645),
            .I(a_delay_counter_15__N_4220_adj_4817));
    InMux I__4496 (
            .O(N__39642),
            .I(N__39639));
    LocalMux I__4495 (
            .O(N__39639),
            .I(n39_adj_4816));
    InMux I__4494 (
            .O(N__39636),
            .I(N__39632));
    InMux I__4493 (
            .O(N__39635),
            .I(N__39629));
    LocalMux I__4492 (
            .O(N__39632),
            .I(\quad_counter1.a_delay_counter_13 ));
    LocalMux I__4491 (
            .O(N__39629),
            .I(\quad_counter1.a_delay_counter_13 ));
    InMux I__4490 (
            .O(N__39624),
            .I(N__39620));
    InMux I__4489 (
            .O(N__39623),
            .I(N__39617));
    LocalMux I__4488 (
            .O(N__39620),
            .I(\quad_counter1.a_delay_counter_2 ));
    LocalMux I__4487 (
            .O(N__39617),
            .I(\quad_counter1.a_delay_counter_2 ));
    CascadeMux I__4486 (
            .O(N__39612),
            .I(N__39608));
    InMux I__4485 (
            .O(N__39611),
            .I(N__39605));
    InMux I__4484 (
            .O(N__39608),
            .I(N__39602));
    LocalMux I__4483 (
            .O(N__39605),
            .I(\quad_counter1.a_delay_counter_1 ));
    LocalMux I__4482 (
            .O(N__39602),
            .I(\quad_counter1.a_delay_counter_1 ));
    InMux I__4481 (
            .O(N__39597),
            .I(N__39593));
    InMux I__4480 (
            .O(N__39596),
            .I(N__39590));
    LocalMux I__4479 (
            .O(N__39593),
            .I(\quad_counter1.a_delay_counter_5 ));
    LocalMux I__4478 (
            .O(N__39590),
            .I(\quad_counter1.a_delay_counter_5 ));
    InMux I__4477 (
            .O(N__39585),
            .I(N__39581));
    InMux I__4476 (
            .O(N__39584),
            .I(N__39578));
    LocalMux I__4475 (
            .O(N__39581),
            .I(\quad_counter1.a_delay_counter_9 ));
    LocalMux I__4474 (
            .O(N__39578),
            .I(\quad_counter1.a_delay_counter_9 ));
    CascadeMux I__4473 (
            .O(N__39573),
            .I(N__39570));
    InMux I__4472 (
            .O(N__39570),
            .I(N__39567));
    LocalMux I__4471 (
            .O(N__39567),
            .I(N__39562));
    InMux I__4470 (
            .O(N__39566),
            .I(N__39559));
    InMux I__4469 (
            .O(N__39565),
            .I(N__39556));
    Odrv4 I__4468 (
            .O(N__39562),
            .I(a_delay_counter_0_adj_4811));
    LocalMux I__4467 (
            .O(N__39559),
            .I(a_delay_counter_0_adj_4811));
    LocalMux I__4466 (
            .O(N__39556),
            .I(a_delay_counter_0_adj_4811));
    CascadeMux I__4465 (
            .O(N__39549),
            .I(N__39545));
    InMux I__4464 (
            .O(N__39548),
            .I(N__39542));
    InMux I__4463 (
            .O(N__39545),
            .I(N__39539));
    LocalMux I__4462 (
            .O(N__39542),
            .I(\quad_counter1.a_delay_counter_3 ));
    LocalMux I__4461 (
            .O(N__39539),
            .I(\quad_counter1.a_delay_counter_3 ));
    InMux I__4460 (
            .O(N__39534),
            .I(N__39530));
    InMux I__4459 (
            .O(N__39533),
            .I(N__39527));
    LocalMux I__4458 (
            .O(N__39530),
            .I(\quad_counter1.a_delay_counter_4 ));
    LocalMux I__4457 (
            .O(N__39527),
            .I(\quad_counter1.a_delay_counter_4 ));
    InMux I__4456 (
            .O(N__39522),
            .I(N__39518));
    InMux I__4455 (
            .O(N__39521),
            .I(N__39515));
    LocalMux I__4454 (
            .O(N__39518),
            .I(\quad_counter1.a_delay_counter_14 ));
    LocalMux I__4453 (
            .O(N__39515),
            .I(\quad_counter1.a_delay_counter_14 ));
    InMux I__4452 (
            .O(N__39510),
            .I(N__39506));
    InMux I__4451 (
            .O(N__39509),
            .I(N__39503));
    LocalMux I__4450 (
            .O(N__39506),
            .I(\quad_counter1.a_delay_counter_7 ));
    LocalMux I__4449 (
            .O(N__39503),
            .I(\quad_counter1.a_delay_counter_7 ));
    CascadeMux I__4448 (
            .O(N__39498),
            .I(N__39494));
    InMux I__4447 (
            .O(N__39497),
            .I(N__39491));
    InMux I__4446 (
            .O(N__39494),
            .I(N__39488));
    LocalMux I__4445 (
            .O(N__39491),
            .I(\quad_counter1.a_delay_counter_12 ));
    LocalMux I__4444 (
            .O(N__39488),
            .I(\quad_counter1.a_delay_counter_12 ));
    InMux I__4443 (
            .O(N__39483),
            .I(N__39479));
    InMux I__4442 (
            .O(N__39482),
            .I(N__39476));
    LocalMux I__4441 (
            .O(N__39479),
            .I(\quad_counter1.a_delay_counter_15 ));
    LocalMux I__4440 (
            .O(N__39476),
            .I(\quad_counter1.a_delay_counter_15 ));
    InMux I__4439 (
            .O(N__39471),
            .I(N__39468));
    LocalMux I__4438 (
            .O(N__39468),
            .I(\quad_counter1.n25_adj_4443 ));
    CascadeMux I__4437 (
            .O(N__39465),
            .I(\quad_counter1.n27_adj_4442_cascade_ ));
    InMux I__4436 (
            .O(N__39462),
            .I(N__39459));
    LocalMux I__4435 (
            .O(N__39459),
            .I(\quad_counter1.n28_adj_4440 ));
    InMux I__4434 (
            .O(N__39456),
            .I(N__39452));
    CascadeMux I__4433 (
            .O(N__39455),
            .I(N__39448));
    LocalMux I__4432 (
            .O(N__39452),
            .I(N__39445));
    InMux I__4431 (
            .O(N__39451),
            .I(N__39440));
    InMux I__4430 (
            .O(N__39448),
            .I(N__39440));
    Odrv12 I__4429 (
            .O(N__39445),
            .I(\c0.data_in_frame_11_0 ));
    LocalMux I__4428 (
            .O(N__39440),
            .I(\c0.data_in_frame_11_0 ));
    InMux I__4427 (
            .O(N__39435),
            .I(N__39432));
    LocalMux I__4426 (
            .O(N__39432),
            .I(\c0.n6_adj_4713 ));
    InMux I__4425 (
            .O(N__39429),
            .I(N__39423));
    InMux I__4424 (
            .O(N__39428),
            .I(N__39423));
    LocalMux I__4423 (
            .O(N__39423),
            .I(N__39420));
    Span4Mux_h I__4422 (
            .O(N__39420),
            .I(N__39417));
    Sp12to4 I__4421 (
            .O(N__39417),
            .I(N__39413));
    InMux I__4420 (
            .O(N__39416),
            .I(N__39410));
    Span12Mux_v I__4419 (
            .O(N__39413),
            .I(N__39407));
    LocalMux I__4418 (
            .O(N__39410),
            .I(B_filtered));
    Odrv12 I__4417 (
            .O(N__39407),
            .I(B_filtered));
    InMux I__4416 (
            .O(N__39402),
            .I(N__39395));
    InMux I__4415 (
            .O(N__39401),
            .I(N__39395));
    InMux I__4414 (
            .O(N__39400),
            .I(N__39392));
    LocalMux I__4413 (
            .O(N__39395),
            .I(N__39389));
    LocalMux I__4412 (
            .O(N__39392),
            .I(\quad_counter0.B_delayed ));
    Odrv4 I__4411 (
            .O(N__39389),
            .I(\quad_counter0.B_delayed ));
    InMux I__4410 (
            .O(N__39384),
            .I(N__39381));
    LocalMux I__4409 (
            .O(N__39381),
            .I(N__39378));
    Odrv4 I__4408 (
            .O(N__39378),
            .I(\c0.n33714 ));
    InMux I__4407 (
            .O(N__39375),
            .I(N__39372));
    LocalMux I__4406 (
            .O(N__39372),
            .I(N__39369));
    Odrv4 I__4405 (
            .O(N__39369),
            .I(\c0.n33923 ));
    CascadeMux I__4404 (
            .O(N__39366),
            .I(\c0.n33982_cascade_ ));
    CascadeMux I__4403 (
            .O(N__39363),
            .I(N__39358));
    InMux I__4402 (
            .O(N__39362),
            .I(N__39353));
    InMux I__4401 (
            .O(N__39361),
            .I(N__39353));
    InMux I__4400 (
            .O(N__39358),
            .I(N__39350));
    LocalMux I__4399 (
            .O(N__39353),
            .I(N__39347));
    LocalMux I__4398 (
            .O(N__39350),
            .I(\c0.data_in_frame_10_5 ));
    Odrv4 I__4397 (
            .O(N__39347),
            .I(\c0.data_in_frame_10_5 ));
    InMux I__4396 (
            .O(N__39342),
            .I(N__39339));
    LocalMux I__4395 (
            .O(N__39339),
            .I(N__39336));
    Odrv4 I__4394 (
            .O(N__39336),
            .I(\c0.n33997 ));
    CascadeMux I__4393 (
            .O(N__39333),
            .I(\c0.n33997_cascade_ ));
    InMux I__4392 (
            .O(N__39330),
            .I(N__39322));
    InMux I__4391 (
            .O(N__39329),
            .I(N__39322));
    InMux I__4390 (
            .O(N__39328),
            .I(N__39319));
    InMux I__4389 (
            .O(N__39327),
            .I(N__39316));
    LocalMux I__4388 (
            .O(N__39322),
            .I(N__39311));
    LocalMux I__4387 (
            .O(N__39319),
            .I(N__39311));
    LocalMux I__4386 (
            .O(N__39316),
            .I(\c0.data_in_frame_10_7 ));
    Odrv4 I__4385 (
            .O(N__39311),
            .I(\c0.data_in_frame_10_7 ));
    InMux I__4384 (
            .O(N__39306),
            .I(N__39303));
    LocalMux I__4383 (
            .O(N__39303),
            .I(\quad_counter0.A_delayed ));
    CascadeMux I__4382 (
            .O(N__39300),
            .I(N__39296));
    InMux I__4381 (
            .O(N__39299),
            .I(N__39290));
    InMux I__4380 (
            .O(N__39296),
            .I(N__39290));
    CascadeMux I__4379 (
            .O(N__39295),
            .I(N__39285));
    LocalMux I__4378 (
            .O(N__39290),
            .I(N__39282));
    InMux I__4377 (
            .O(N__39289),
            .I(N__39277));
    InMux I__4376 (
            .O(N__39288),
            .I(N__39277));
    InMux I__4375 (
            .O(N__39285),
            .I(N__39274));
    Span12Mux_h I__4374 (
            .O(N__39282),
            .I(N__39269));
    LocalMux I__4373 (
            .O(N__39277),
            .I(N__39269));
    LocalMux I__4372 (
            .O(N__39274),
            .I(N__39264));
    Span12Mux_v I__4371 (
            .O(N__39269),
            .I(N__39264));
    Odrv12 I__4370 (
            .O(N__39264),
            .I(A_filtered));
    InMux I__4369 (
            .O(N__39261),
            .I(N__39257));
    InMux I__4368 (
            .O(N__39260),
            .I(N__39254));
    LocalMux I__4367 (
            .O(N__39257),
            .I(N__39249));
    LocalMux I__4366 (
            .O(N__39254),
            .I(N__39249));
    Odrv12 I__4365 (
            .O(N__39249),
            .I(\c0.n33695 ));
    InMux I__4364 (
            .O(N__39246),
            .I(N__39242));
    InMux I__4363 (
            .O(N__39245),
            .I(N__39238));
    LocalMux I__4362 (
            .O(N__39242),
            .I(N__39235));
    InMux I__4361 (
            .O(N__39241),
            .I(N__39232));
    LocalMux I__4360 (
            .O(N__39238),
            .I(N__39229));
    Span4Mux_v I__4359 (
            .O(N__39235),
            .I(N__39224));
    LocalMux I__4358 (
            .O(N__39232),
            .I(N__39224));
    Odrv12 I__4357 (
            .O(N__39229),
            .I(\c0.n18671 ));
    Odrv4 I__4356 (
            .O(N__39224),
            .I(\c0.n18671 ));
    CascadeMux I__4355 (
            .O(N__39219),
            .I(\c0.n10_adj_4769_cascade_ ));
    InMux I__4354 (
            .O(N__39216),
            .I(N__39211));
    InMux I__4353 (
            .O(N__39215),
            .I(N__39208));
    CascadeMux I__4352 (
            .O(N__39214),
            .I(N__39205));
    LocalMux I__4351 (
            .O(N__39211),
            .I(N__39202));
    LocalMux I__4350 (
            .O(N__39208),
            .I(N__39199));
    InMux I__4349 (
            .O(N__39205),
            .I(N__39196));
    Span4Mux_h I__4348 (
            .O(N__39202),
            .I(N__39191));
    Span4Mux_h I__4347 (
            .O(N__39199),
            .I(N__39191));
    LocalMux I__4346 (
            .O(N__39196),
            .I(\c0.data_in_frame_4_4 ));
    Odrv4 I__4345 (
            .O(N__39191),
            .I(\c0.data_in_frame_4_4 ));
    CascadeMux I__4344 (
            .O(N__39186),
            .I(\c0.n18330_cascade_ ));
    InMux I__4343 (
            .O(N__39183),
            .I(N__39177));
    InMux I__4342 (
            .O(N__39182),
            .I(N__39177));
    LocalMux I__4341 (
            .O(N__39177),
            .I(\c0.data_in_frame_6_5 ));
    InMux I__4340 (
            .O(N__39174),
            .I(N__39171));
    LocalMux I__4339 (
            .O(N__39171),
            .I(N__39167));
    InMux I__4338 (
            .O(N__39170),
            .I(N__39164));
    Span4Mux_v I__4337 (
            .O(N__39167),
            .I(N__39159));
    LocalMux I__4336 (
            .O(N__39164),
            .I(N__39159));
    Odrv4 I__4335 (
            .O(N__39159),
            .I(n4));
    CascadeMux I__4334 (
            .O(N__39156),
            .I(N__39152));
    CascadeMux I__4333 (
            .O(N__39155),
            .I(N__39149));
    InMux I__4332 (
            .O(N__39152),
            .I(N__39145));
    InMux I__4331 (
            .O(N__39149),
            .I(N__39142));
    InMux I__4330 (
            .O(N__39148),
            .I(N__39139));
    LocalMux I__4329 (
            .O(N__39145),
            .I(N__39134));
    LocalMux I__4328 (
            .O(N__39142),
            .I(N__39134));
    LocalMux I__4327 (
            .O(N__39139),
            .I(\c0.data_in_frame_11_2 ));
    Odrv4 I__4326 (
            .O(N__39134),
            .I(\c0.data_in_frame_11_2 ));
    InMux I__4325 (
            .O(N__39129),
            .I(N__39126));
    LocalMux I__4324 (
            .O(N__39126),
            .I(N__39123));
    Odrv4 I__4323 (
            .O(N__39123),
            .I(\c0.n33985 ));
    CascadeMux I__4322 (
            .O(N__39120),
            .I(\c0.n33714_cascade_ ));
    CascadeMux I__4321 (
            .O(N__39117),
            .I(N__39113));
    InMux I__4320 (
            .O(N__39116),
            .I(N__39109));
    InMux I__4319 (
            .O(N__39113),
            .I(N__39104));
    InMux I__4318 (
            .O(N__39112),
            .I(N__39104));
    LocalMux I__4317 (
            .O(N__39109),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__4316 (
            .O(N__39104),
            .I(\c0.data_in_frame_2_3 ));
    InMux I__4315 (
            .O(N__39099),
            .I(N__39096));
    LocalMux I__4314 (
            .O(N__39096),
            .I(\c0.n6_adj_4564 ));
    CascadeMux I__4313 (
            .O(N__39093),
            .I(\c0.n5452_cascade_ ));
    CascadeMux I__4312 (
            .O(N__39090),
            .I(N__39085));
    InMux I__4311 (
            .O(N__39089),
            .I(N__39080));
    InMux I__4310 (
            .O(N__39088),
            .I(N__39080));
    InMux I__4309 (
            .O(N__39085),
            .I(N__39076));
    LocalMux I__4308 (
            .O(N__39080),
            .I(N__39073));
    InMux I__4307 (
            .O(N__39079),
            .I(N__39070));
    LocalMux I__4306 (
            .O(N__39076),
            .I(\c0.data_in_frame_4_5 ));
    Odrv4 I__4305 (
            .O(N__39073),
            .I(\c0.data_in_frame_4_5 ));
    LocalMux I__4304 (
            .O(N__39070),
            .I(\c0.data_in_frame_4_5 ));
    CascadeMux I__4303 (
            .O(N__39063),
            .I(\c0.n19030_cascade_ ));
    CascadeMux I__4302 (
            .O(N__39060),
            .I(\c0.n33215_cascade_ ));
    CascadeMux I__4301 (
            .O(N__39057),
            .I(N__39054));
    InMux I__4300 (
            .O(N__39054),
            .I(N__39051));
    LocalMux I__4299 (
            .O(N__39051),
            .I(\c0.n6_adj_4616 ));
    InMux I__4298 (
            .O(N__39048),
            .I(N__39042));
    InMux I__4297 (
            .O(N__39047),
            .I(N__39042));
    LocalMux I__4296 (
            .O(N__39042),
            .I(N__39037));
    InMux I__4295 (
            .O(N__39041),
            .I(N__39032));
    InMux I__4294 (
            .O(N__39040),
            .I(N__39032));
    Odrv4 I__4293 (
            .O(N__39037),
            .I(\c0.n33263 ));
    LocalMux I__4292 (
            .O(N__39032),
            .I(\c0.n33263 ));
    CascadeMux I__4291 (
            .O(N__39027),
            .I(N__39023));
    InMux I__4290 (
            .O(N__39026),
            .I(N__39019));
    InMux I__4289 (
            .O(N__39023),
            .I(N__39014));
    InMux I__4288 (
            .O(N__39022),
            .I(N__39014));
    LocalMux I__4287 (
            .O(N__39019),
            .I(N__39011));
    LocalMux I__4286 (
            .O(N__39014),
            .I(N__39008));
    Span4Mux_h I__4285 (
            .O(N__39011),
            .I(N__39005));
    Odrv4 I__4284 (
            .O(N__39008),
            .I(\c0.n29676 ));
    Odrv4 I__4283 (
            .O(N__39005),
            .I(\c0.n29676 ));
    InMux I__4282 (
            .O(N__39000),
            .I(N__38997));
    LocalMux I__4281 (
            .O(N__38997),
            .I(\c0.n10800 ));
    InMux I__4280 (
            .O(N__38994),
            .I(N__38988));
    InMux I__4279 (
            .O(N__38993),
            .I(N__38988));
    LocalMux I__4278 (
            .O(N__38988),
            .I(N__38985));
    Span4Mux_v I__4277 (
            .O(N__38985),
            .I(N__38981));
    InMux I__4276 (
            .O(N__38984),
            .I(N__38978));
    Odrv4 I__4275 (
            .O(N__38981),
            .I(\c0.data_out_frame_0__7__N_2568 ));
    LocalMux I__4274 (
            .O(N__38978),
            .I(\c0.data_out_frame_0__7__N_2568 ));
    InMux I__4273 (
            .O(N__38973),
            .I(N__38969));
    InMux I__4272 (
            .O(N__38972),
            .I(N__38966));
    LocalMux I__4271 (
            .O(N__38969),
            .I(N__38963));
    LocalMux I__4270 (
            .O(N__38966),
            .I(N__38959));
    Span4Mux_h I__4269 (
            .O(N__38963),
            .I(N__38956));
    InMux I__4268 (
            .O(N__38962),
            .I(N__38953));
    Odrv4 I__4267 (
            .O(N__38959),
            .I(\c0.n22387 ));
    Odrv4 I__4266 (
            .O(N__38956),
            .I(\c0.n22387 ));
    LocalMux I__4265 (
            .O(N__38953),
            .I(\c0.n22387 ));
    CascadeMux I__4264 (
            .O(N__38946),
            .I(\c0.n10800_cascade_ ));
    InMux I__4263 (
            .O(N__38943),
            .I(N__38940));
    LocalMux I__4262 (
            .O(N__38940),
            .I(\c0.n4_adj_4615 ));
    CascadeMux I__4261 (
            .O(N__38937),
            .I(N__38934));
    InMux I__4260 (
            .O(N__38934),
            .I(N__38931));
    LocalMux I__4259 (
            .O(N__38931),
            .I(N__38928));
    Odrv4 I__4258 (
            .O(N__38928),
            .I(\c0.FRAME_MATCHER_state_1 ));
    CascadeMux I__4257 (
            .O(N__38925),
            .I(N__38921));
    InMux I__4256 (
            .O(N__38924),
            .I(N__38918));
    InMux I__4255 (
            .O(N__38921),
            .I(N__38913));
    LocalMux I__4254 (
            .O(N__38918),
            .I(N__38910));
    InMux I__4253 (
            .O(N__38917),
            .I(N__38907));
    InMux I__4252 (
            .O(N__38916),
            .I(N__38904));
    LocalMux I__4251 (
            .O(N__38913),
            .I(N__38899));
    Span4Mux_v I__4250 (
            .O(N__38910),
            .I(N__38899));
    LocalMux I__4249 (
            .O(N__38907),
            .I(N__38896));
    LocalMux I__4248 (
            .O(N__38904),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__4247 (
            .O(N__38899),
            .I(\c0.data_in_frame_7_0 ));
    Odrv4 I__4246 (
            .O(N__38896),
            .I(\c0.data_in_frame_7_0 ));
    CascadeMux I__4245 (
            .O(N__38889),
            .I(N__38886));
    InMux I__4244 (
            .O(N__38886),
            .I(N__38882));
    CascadeMux I__4243 (
            .O(N__38885),
            .I(N__38878));
    LocalMux I__4242 (
            .O(N__38882),
            .I(N__38874));
    CascadeMux I__4241 (
            .O(N__38881),
            .I(N__38871));
    InMux I__4240 (
            .O(N__38878),
            .I(N__38866));
    InMux I__4239 (
            .O(N__38877),
            .I(N__38866));
    Span4Mux_h I__4238 (
            .O(N__38874),
            .I(N__38863));
    InMux I__4237 (
            .O(N__38871),
            .I(N__38860));
    LocalMux I__4236 (
            .O(N__38866),
            .I(\c0.data_in_frame_9_1 ));
    Odrv4 I__4235 (
            .O(N__38863),
            .I(\c0.data_in_frame_9_1 ));
    LocalMux I__4234 (
            .O(N__38860),
            .I(\c0.data_in_frame_9_1 ));
    InMux I__4233 (
            .O(N__38853),
            .I(N__38850));
    LocalMux I__4232 (
            .O(N__38850),
            .I(N__38847));
    Odrv4 I__4231 (
            .O(N__38847),
            .I(\c0.n93 ));
    CascadeMux I__4230 (
            .O(N__38844),
            .I(N__38841));
    InMux I__4229 (
            .O(N__38841),
            .I(N__38838));
    LocalMux I__4228 (
            .O(N__38838),
            .I(\quad_counter0.n20_adj_4351 ));
    CascadeMux I__4227 (
            .O(N__38835),
            .I(\quad_counter0.n22_adj_4350_cascade_ ));
    InMux I__4226 (
            .O(N__38832),
            .I(N__38829));
    LocalMux I__4225 (
            .O(N__38829),
            .I(\quad_counter0.n16 ));
    InMux I__4224 (
            .O(N__38826),
            .I(N__38823));
    LocalMux I__4223 (
            .O(N__38823),
            .I(\quad_counter0.n24_adj_4352 ));
    InMux I__4222 (
            .O(N__38820),
            .I(N__38817));
    LocalMux I__4221 (
            .O(N__38817),
            .I(N__38814));
    Span4Mux_v I__4220 (
            .O(N__38814),
            .I(N__38811));
    Odrv4 I__4219 (
            .O(N__38811),
            .I(\c0.n11_adj_4614 ));
    CascadeMux I__4218 (
            .O(N__38808),
            .I(N__38805));
    InMux I__4217 (
            .O(N__38805),
            .I(N__38802));
    LocalMux I__4216 (
            .O(N__38802),
            .I(N__38799));
    Odrv4 I__4215 (
            .O(N__38799),
            .I(\c0.FRAME_MATCHER_state_2 ));
    CascadeMux I__4214 (
            .O(N__38796),
            .I(N__38793));
    InMux I__4213 (
            .O(N__38793),
            .I(N__38790));
    LocalMux I__4212 (
            .O(N__38790),
            .I(\c0.n3844 ));
    InMux I__4211 (
            .O(N__38787),
            .I(N__38784));
    LocalMux I__4210 (
            .O(N__38784),
            .I(\c0.n6_adj_4618 ));
    InMux I__4209 (
            .O(N__38781),
            .I(\quad_counter0.n30359 ));
    InMux I__4208 (
            .O(N__38778),
            .I(\quad_counter0.n30360 ));
    InMux I__4207 (
            .O(N__38775),
            .I(\quad_counter0.n30361 ));
    InMux I__4206 (
            .O(N__38772),
            .I(bfn_9_15_0_));
    InMux I__4205 (
            .O(N__38769),
            .I(\quad_counter0.n30363 ));
    InMux I__4204 (
            .O(N__38766),
            .I(\quad_counter0.n30364 ));
    CascadeMux I__4203 (
            .O(N__38763),
            .I(N__38755));
    CascadeMux I__4202 (
            .O(N__38762),
            .I(N__38752));
    CascadeMux I__4201 (
            .O(N__38761),
            .I(N__38749));
    CascadeMux I__4200 (
            .O(N__38760),
            .I(N__38746));
    CascadeMux I__4199 (
            .O(N__38759),
            .I(N__38743));
    CascadeMux I__4198 (
            .O(N__38758),
            .I(N__38740));
    InMux I__4197 (
            .O(N__38755),
            .I(N__38735));
    InMux I__4196 (
            .O(N__38752),
            .I(N__38735));
    InMux I__4195 (
            .O(N__38749),
            .I(N__38726));
    InMux I__4194 (
            .O(N__38746),
            .I(N__38726));
    InMux I__4193 (
            .O(N__38743),
            .I(N__38726));
    InMux I__4192 (
            .O(N__38740),
            .I(N__38726));
    LocalMux I__4191 (
            .O(N__38735),
            .I(N__38721));
    LocalMux I__4190 (
            .O(N__38726),
            .I(N__38721));
    Odrv4 I__4189 (
            .O(N__38721),
            .I(\quad_counter0.n36144 ));
    InMux I__4188 (
            .O(N__38718),
            .I(N__38715));
    LocalMux I__4187 (
            .O(N__38715),
            .I(N__38712));
    Odrv4 I__4186 (
            .O(N__38712),
            .I(\quad_counter0.n24_adj_4354 ));
    CascadeMux I__4185 (
            .O(N__38709),
            .I(N__38696));
    CascadeMux I__4184 (
            .O(N__38708),
            .I(N__38693));
    CascadeMux I__4183 (
            .O(N__38707),
            .I(N__38688));
    CascadeMux I__4182 (
            .O(N__38706),
            .I(N__38685));
    CascadeMux I__4181 (
            .O(N__38705),
            .I(N__38682));
    CascadeMux I__4180 (
            .O(N__38704),
            .I(N__38679));
    CascadeMux I__4179 (
            .O(N__38703),
            .I(N__38676));
    CascadeMux I__4178 (
            .O(N__38702),
            .I(N__38673));
    CascadeMux I__4177 (
            .O(N__38701),
            .I(N__38670));
    CascadeMux I__4176 (
            .O(N__38700),
            .I(N__38667));
    CascadeMux I__4175 (
            .O(N__38699),
            .I(N__38664));
    InMux I__4174 (
            .O(N__38696),
            .I(N__38659));
    InMux I__4173 (
            .O(N__38693),
            .I(N__38659));
    CascadeMux I__4172 (
            .O(N__38692),
            .I(N__38656));
    CascadeMux I__4171 (
            .O(N__38691),
            .I(N__38653));
    InMux I__4170 (
            .O(N__38688),
            .I(N__38649));
    InMux I__4169 (
            .O(N__38685),
            .I(N__38640));
    InMux I__4168 (
            .O(N__38682),
            .I(N__38640));
    InMux I__4167 (
            .O(N__38679),
            .I(N__38640));
    InMux I__4166 (
            .O(N__38676),
            .I(N__38640));
    InMux I__4165 (
            .O(N__38673),
            .I(N__38631));
    InMux I__4164 (
            .O(N__38670),
            .I(N__38631));
    InMux I__4163 (
            .O(N__38667),
            .I(N__38631));
    InMux I__4162 (
            .O(N__38664),
            .I(N__38631));
    LocalMux I__4161 (
            .O(N__38659),
            .I(N__38628));
    InMux I__4160 (
            .O(N__38656),
            .I(N__38621));
    InMux I__4159 (
            .O(N__38653),
            .I(N__38621));
    InMux I__4158 (
            .O(N__38652),
            .I(N__38621));
    LocalMux I__4157 (
            .O(N__38649),
            .I(\quad_counter0.n3035 ));
    LocalMux I__4156 (
            .O(N__38640),
            .I(\quad_counter0.n3035 ));
    LocalMux I__4155 (
            .O(N__38631),
            .I(\quad_counter0.n3035 ));
    Odrv4 I__4154 (
            .O(N__38628),
            .I(\quad_counter0.n3035 ));
    LocalMux I__4153 (
            .O(N__38621),
            .I(\quad_counter0.n3035 ));
    InMux I__4152 (
            .O(N__38610),
            .I(\quad_counter0.n30350 ));
    InMux I__4151 (
            .O(N__38607),
            .I(\quad_counter0.n30351 ));
    InMux I__4150 (
            .O(N__38604),
            .I(\quad_counter0.n30352 ));
    InMux I__4149 (
            .O(N__38601),
            .I(\quad_counter0.n30353 ));
    InMux I__4148 (
            .O(N__38598),
            .I(bfn_9_14_0_));
    InMux I__4147 (
            .O(N__38595),
            .I(\quad_counter0.n30355 ));
    InMux I__4146 (
            .O(N__38592),
            .I(\quad_counter0.n30356 ));
    InMux I__4145 (
            .O(N__38589),
            .I(\quad_counter0.n30357 ));
    InMux I__4144 (
            .O(N__38586),
            .I(\quad_counter0.n30358 ));
    CascadeMux I__4143 (
            .O(N__38583),
            .I(\quad_counter0.n18_adj_4353_cascade_ ));
    CascadeMux I__4142 (
            .O(N__38580),
            .I(\quad_counter0.n7_cascade_ ));
    CascadeMux I__4141 (
            .O(N__38577),
            .I(\quad_counter0.n34617_cascade_ ));
    CascadeMux I__4140 (
            .O(N__38574),
            .I(\quad_counter0.n22_adj_4355_cascade_ ));
    InMux I__4139 (
            .O(N__38571),
            .I(N__38568));
    LocalMux I__4138 (
            .O(N__38568),
            .I(\quad_counter0.n26_adj_4356 ));
    InMux I__4137 (
            .O(N__38565),
            .I(bfn_9_13_0_));
    InMux I__4136 (
            .O(N__38562),
            .I(\quad_counter0.n30347 ));
    InMux I__4135 (
            .O(N__38559),
            .I(\quad_counter0.n30348 ));
    InMux I__4134 (
            .O(N__38556),
            .I(\quad_counter0.n30349 ));
    InMux I__4133 (
            .O(N__38553),
            .I(N__38550));
    LocalMux I__4132 (
            .O(N__38550),
            .I(\quad_counter0.n27_adj_4366 ));
    InMux I__4131 (
            .O(N__38547),
            .I(N__38544));
    LocalMux I__4130 (
            .O(N__38544),
            .I(\quad_counter0.n28_adj_4364 ));
    InMux I__4129 (
            .O(N__38541),
            .I(N__38538));
    LocalMux I__4128 (
            .O(N__38538),
            .I(\quad_counter0.n26_adj_4365 ));
    InMux I__4127 (
            .O(N__38535),
            .I(N__38532));
    LocalMux I__4126 (
            .O(N__38532),
            .I(N__38529));
    Odrv4 I__4125 (
            .O(N__38529),
            .I(\quad_counter0.n19 ));
    CascadeMux I__4124 (
            .O(N__38526),
            .I(\quad_counter0.n28_adj_4361_cascade_ ));
    InMux I__4123 (
            .O(N__38523),
            .I(N__38520));
    LocalMux I__4122 (
            .O(N__38520),
            .I(\quad_counter0.n24_adj_4360 ));
    InMux I__4121 (
            .O(N__38517),
            .I(N__38514));
    LocalMux I__4120 (
            .O(N__38514),
            .I(N__38511));
    Odrv4 I__4119 (
            .O(N__38511),
            .I(\c0.rx.r_Rx_Data_R ));
    InMux I__4118 (
            .O(N__38508),
            .I(\quad_counter1.n30056 ));
    InMux I__4117 (
            .O(N__38505),
            .I(\quad_counter1.n30057 ));
    InMux I__4116 (
            .O(N__38502),
            .I(\quad_counter1.n30058 ));
    InMux I__4115 (
            .O(N__38499),
            .I(\quad_counter1.n30059 ));
    InMux I__4114 (
            .O(N__38496),
            .I(\quad_counter1.n30060 ));
    InMux I__4113 (
            .O(N__38493),
            .I(N__38490));
    LocalMux I__4112 (
            .O(N__38490),
            .I(N__38487));
    Span4Mux_v I__4111 (
            .O(N__38487),
            .I(N__38484));
    Sp12to4 I__4110 (
            .O(N__38484),
            .I(N__38480));
    InMux I__4109 (
            .O(N__38483),
            .I(N__38477));
    Span12Mux_h I__4108 (
            .O(N__38480),
            .I(N__38474));
    LocalMux I__4107 (
            .O(N__38477),
            .I(N__38471));
    Span12Mux_v I__4106 (
            .O(N__38474),
            .I(N__38466));
    Span12Mux_h I__4105 (
            .O(N__38471),
            .I(N__38466));
    Odrv12 I__4104 (
            .O(N__38466),
            .I(rx_i));
    CascadeMux I__4103 (
            .O(N__38463),
            .I(\quad_counter0.n25_adj_4367_cascade_ ));
    InMux I__4102 (
            .O(N__38460),
            .I(\quad_counter1.n30047 ));
    InMux I__4101 (
            .O(N__38457),
            .I(\quad_counter1.n30048 ));
    InMux I__4100 (
            .O(N__38454),
            .I(\quad_counter1.n30049 ));
    InMux I__4099 (
            .O(N__38451),
            .I(\quad_counter1.n30050 ));
    InMux I__4098 (
            .O(N__38448),
            .I(\quad_counter1.n30051 ));
    InMux I__4097 (
            .O(N__38445),
            .I(\quad_counter1.n30052 ));
    InMux I__4096 (
            .O(N__38442),
            .I(bfn_9_8_0_));
    InMux I__4095 (
            .O(N__38439),
            .I(\quad_counter1.n30054 ));
    InMux I__4094 (
            .O(N__38436),
            .I(\quad_counter1.n30055 ));
    InMux I__4093 (
            .O(N__38433),
            .I(bfn_9_7_0_));
    InMux I__4092 (
            .O(N__38430),
            .I(\quad_counter1.n30046 ));
    CascadeMux I__4091 (
            .O(N__38427),
            .I(\c0.n33985_cascade_ ));
    InMux I__4090 (
            .O(N__38424),
            .I(N__38419));
    InMux I__4089 (
            .O(N__38423),
            .I(N__38414));
    InMux I__4088 (
            .O(N__38422),
            .I(N__38414));
    LocalMux I__4087 (
            .O(N__38419),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__4086 (
            .O(N__38414),
            .I(\c0.data_in_frame_7_1 ));
    InMux I__4085 (
            .O(N__38409),
            .I(N__38403));
    InMux I__4084 (
            .O(N__38408),
            .I(N__38403));
    LocalMux I__4083 (
            .O(N__38403),
            .I(\c0.n33444 ));
    CascadeMux I__4082 (
            .O(N__38400),
            .I(N__38395));
    CascadeMux I__4081 (
            .O(N__38399),
            .I(N__38392));
    CascadeMux I__4080 (
            .O(N__38398),
            .I(N__38389));
    InMux I__4079 (
            .O(N__38395),
            .I(N__38386));
    InMux I__4078 (
            .O(N__38392),
            .I(N__38383));
    InMux I__4077 (
            .O(N__38389),
            .I(N__38380));
    LocalMux I__4076 (
            .O(N__38386),
            .I(N__38377));
    LocalMux I__4075 (
            .O(N__38383),
            .I(N__38374));
    LocalMux I__4074 (
            .O(N__38380),
            .I(\c0.data_in_frame_5_0 ));
    Odrv4 I__4073 (
            .O(N__38377),
            .I(\c0.data_in_frame_5_0 ));
    Odrv4 I__4072 (
            .O(N__38374),
            .I(\c0.data_in_frame_5_0 ));
    InMux I__4071 (
            .O(N__38367),
            .I(N__38363));
    InMux I__4070 (
            .O(N__38366),
            .I(N__38360));
    LocalMux I__4069 (
            .O(N__38363),
            .I(N__38357));
    LocalMux I__4068 (
            .O(N__38360),
            .I(\c0.data_in_frame_9_2 ));
    Odrv4 I__4067 (
            .O(N__38357),
            .I(\c0.data_in_frame_9_2 ));
    CascadeMux I__4066 (
            .O(N__38352),
            .I(N__38349));
    InMux I__4065 (
            .O(N__38349),
            .I(N__38343));
    InMux I__4064 (
            .O(N__38348),
            .I(N__38343));
    LocalMux I__4063 (
            .O(N__38343),
            .I(\c0.data_in_frame_9_6 ));
    CascadeMux I__4062 (
            .O(N__38340),
            .I(\c0.n8_adj_4508_cascade_ ));
    InMux I__4061 (
            .O(N__38337),
            .I(N__38332));
    InMux I__4060 (
            .O(N__38336),
            .I(N__38327));
    InMux I__4059 (
            .O(N__38335),
            .I(N__38327));
    LocalMux I__4058 (
            .O(N__38332),
            .I(N__38324));
    LocalMux I__4057 (
            .O(N__38327),
            .I(N__38320));
    Span4Mux_h I__4056 (
            .O(N__38324),
            .I(N__38317));
    InMux I__4055 (
            .O(N__38323),
            .I(N__38314));
    Span4Mux_h I__4054 (
            .O(N__38320),
            .I(N__38311));
    Odrv4 I__4053 (
            .O(N__38317),
            .I(data_in_3_3));
    LocalMux I__4052 (
            .O(N__38314),
            .I(data_in_3_3));
    Odrv4 I__4051 (
            .O(N__38311),
            .I(data_in_3_3));
    CascadeMux I__4050 (
            .O(N__38304),
            .I(N__38300));
    CascadeMux I__4049 (
            .O(N__38303),
            .I(N__38297));
    InMux I__4048 (
            .O(N__38300),
            .I(N__38294));
    InMux I__4047 (
            .O(N__38297),
            .I(N__38291));
    LocalMux I__4046 (
            .O(N__38294),
            .I(N__38284));
    LocalMux I__4045 (
            .O(N__38291),
            .I(N__38284));
    InMux I__4044 (
            .O(N__38290),
            .I(N__38279));
    InMux I__4043 (
            .O(N__38289),
            .I(N__38279));
    Span4Mux_h I__4042 (
            .O(N__38284),
            .I(N__38276));
    LocalMux I__4041 (
            .O(N__38279),
            .I(data_in_2_3));
    Odrv4 I__4040 (
            .O(N__38276),
            .I(data_in_2_3));
    InMux I__4039 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__4038 (
            .O(N__38268),
            .I(N__38263));
    CascadeMux I__4037 (
            .O(N__38267),
            .I(N__38259));
    InMux I__4036 (
            .O(N__38266),
            .I(N__38256));
    Span4Mux_h I__4035 (
            .O(N__38263),
            .I(N__38253));
    InMux I__4034 (
            .O(N__38262),
            .I(N__38250));
    InMux I__4033 (
            .O(N__38259),
            .I(N__38247));
    LocalMux I__4032 (
            .O(N__38256),
            .I(data_in_1_3));
    Odrv4 I__4031 (
            .O(N__38253),
            .I(data_in_1_3));
    LocalMux I__4030 (
            .O(N__38250),
            .I(data_in_1_3));
    LocalMux I__4029 (
            .O(N__38247),
            .I(data_in_1_3));
    InMux I__4028 (
            .O(N__38238),
            .I(N__38235));
    LocalMux I__4027 (
            .O(N__38235),
            .I(N__38231));
    InMux I__4026 (
            .O(N__38234),
            .I(N__38226));
    Span4Mux_v I__4025 (
            .O(N__38231),
            .I(N__38223));
    InMux I__4024 (
            .O(N__38230),
            .I(N__38218));
    InMux I__4023 (
            .O(N__38229),
            .I(N__38218));
    LocalMux I__4022 (
            .O(N__38226),
            .I(data_in_3_0));
    Odrv4 I__4021 (
            .O(N__38223),
            .I(data_in_3_0));
    LocalMux I__4020 (
            .O(N__38218),
            .I(data_in_3_0));
    InMux I__4019 (
            .O(N__38211),
            .I(N__38206));
    InMux I__4018 (
            .O(N__38210),
            .I(N__38203));
    InMux I__4017 (
            .O(N__38209),
            .I(N__38199));
    LocalMux I__4016 (
            .O(N__38206),
            .I(N__38194));
    LocalMux I__4015 (
            .O(N__38203),
            .I(N__38194));
    InMux I__4014 (
            .O(N__38202),
            .I(N__38191));
    LocalMux I__4013 (
            .O(N__38199),
            .I(data_in_2_0));
    Odrv4 I__4012 (
            .O(N__38194),
            .I(data_in_2_0));
    LocalMux I__4011 (
            .O(N__38191),
            .I(data_in_2_0));
    CascadeMux I__4010 (
            .O(N__38184),
            .I(N__38181));
    InMux I__4009 (
            .O(N__38181),
            .I(N__38174));
    InMux I__4008 (
            .O(N__38180),
            .I(N__38174));
    InMux I__4007 (
            .O(N__38179),
            .I(N__38171));
    LocalMux I__4006 (
            .O(N__38174),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__4005 (
            .O(N__38171),
            .I(\c0.data_in_frame_4_6 ));
    InMux I__4004 (
            .O(N__38166),
            .I(N__38160));
    InMux I__4003 (
            .O(N__38165),
            .I(N__38160));
    LocalMux I__4002 (
            .O(N__38160),
            .I(N__38155));
    InMux I__4001 (
            .O(N__38159),
            .I(N__38152));
    InMux I__4000 (
            .O(N__38158),
            .I(N__38149));
    Span4Mux_h I__3999 (
            .O(N__38155),
            .I(N__38146));
    LocalMux I__3998 (
            .O(N__38152),
            .I(data_in_3_4));
    LocalMux I__3997 (
            .O(N__38149),
            .I(data_in_3_4));
    Odrv4 I__3996 (
            .O(N__38146),
            .I(data_in_3_4));
    InMux I__3995 (
            .O(N__38139),
            .I(N__38136));
    LocalMux I__3994 (
            .O(N__38136),
            .I(N__38132));
    InMux I__3993 (
            .O(N__38135),
            .I(N__38127));
    Span4Mux_h I__3992 (
            .O(N__38132),
            .I(N__38124));
    InMux I__3991 (
            .O(N__38131),
            .I(N__38119));
    InMux I__3990 (
            .O(N__38130),
            .I(N__38119));
    LocalMux I__3989 (
            .O(N__38127),
            .I(data_in_3_6));
    Odrv4 I__3988 (
            .O(N__38124),
            .I(data_in_3_6));
    LocalMux I__3987 (
            .O(N__38119),
            .I(data_in_3_6));
    InMux I__3986 (
            .O(N__38112),
            .I(N__38109));
    LocalMux I__3985 (
            .O(N__38109),
            .I(N__38104));
    CascadeMux I__3984 (
            .O(N__38108),
            .I(N__38100));
    InMux I__3983 (
            .O(N__38107),
            .I(N__38097));
    Span4Mux_v I__3982 (
            .O(N__38104),
            .I(N__38094));
    InMux I__3981 (
            .O(N__38103),
            .I(N__38089));
    InMux I__3980 (
            .O(N__38100),
            .I(N__38089));
    LocalMux I__3979 (
            .O(N__38097),
            .I(N__38086));
    Odrv4 I__3978 (
            .O(N__38094),
            .I(data_in_2_6));
    LocalMux I__3977 (
            .O(N__38089),
            .I(data_in_2_6));
    Odrv4 I__3976 (
            .O(N__38086),
            .I(data_in_2_6));
    InMux I__3975 (
            .O(N__38079),
            .I(N__38071));
    InMux I__3974 (
            .O(N__38078),
            .I(N__38071));
    InMux I__3973 (
            .O(N__38077),
            .I(N__38066));
    InMux I__3972 (
            .O(N__38076),
            .I(N__38066));
    LocalMux I__3971 (
            .O(N__38071),
            .I(data_in_3_2));
    LocalMux I__3970 (
            .O(N__38066),
            .I(data_in_3_2));
    InMux I__3969 (
            .O(N__38061),
            .I(N__38051));
    InMux I__3968 (
            .O(N__38060),
            .I(N__38051));
    InMux I__3967 (
            .O(N__38059),
            .I(N__38051));
    InMux I__3966 (
            .O(N__38058),
            .I(N__38048));
    LocalMux I__3965 (
            .O(N__38051),
            .I(N__38045));
    LocalMux I__3964 (
            .O(N__38048),
            .I(data_in_2_2));
    Odrv4 I__3963 (
            .O(N__38045),
            .I(data_in_2_2));
    InMux I__3962 (
            .O(N__38040),
            .I(N__38034));
    InMux I__3961 (
            .O(N__38039),
            .I(N__38034));
    LocalMux I__3960 (
            .O(N__38034),
            .I(N__38030));
    InMux I__3959 (
            .O(N__38033),
            .I(N__38027));
    Odrv4 I__3958 (
            .O(N__38030),
            .I(\c0.n33266 ));
    LocalMux I__3957 (
            .O(N__38027),
            .I(\c0.n33266 ));
    InMux I__3956 (
            .O(N__38022),
            .I(N__38016));
    InMux I__3955 (
            .O(N__38021),
            .I(N__38016));
    LocalMux I__3954 (
            .O(N__38016),
            .I(N__38013));
    Odrv4 I__3953 (
            .O(N__38013),
            .I(\c0.n63 ));
    CascadeMux I__3952 (
            .O(N__38010),
            .I(N__38005));
    InMux I__3951 (
            .O(N__38009),
            .I(N__38000));
    InMux I__3950 (
            .O(N__38008),
            .I(N__38000));
    InMux I__3949 (
            .O(N__38005),
            .I(N__37997));
    LocalMux I__3948 (
            .O(N__38000),
            .I(N__37994));
    LocalMux I__3947 (
            .O(N__37997),
            .I(N__37991));
    Odrv4 I__3946 (
            .O(N__37994),
            .I(\c0.n107 ));
    Odrv4 I__3945 (
            .O(N__37991),
            .I(\c0.n107 ));
    CascadeMux I__3944 (
            .O(N__37986),
            .I(N__37983));
    InMux I__3943 (
            .O(N__37983),
            .I(N__37977));
    InMux I__3942 (
            .O(N__37982),
            .I(N__37977));
    LocalMux I__3941 (
            .O(N__37977),
            .I(N__37972));
    InMux I__3940 (
            .O(N__37976),
            .I(N__37967));
    InMux I__3939 (
            .O(N__37975),
            .I(N__37967));
    Span4Mux_v I__3938 (
            .O(N__37972),
            .I(N__37962));
    LocalMux I__3937 (
            .O(N__37967),
            .I(N__37962));
    Odrv4 I__3936 (
            .O(N__37962),
            .I(\c0.n14_adj_4784 ));
    InMux I__3935 (
            .O(N__37959),
            .I(N__37953));
    InMux I__3934 (
            .O(N__37958),
            .I(N__37950));
    InMux I__3933 (
            .O(N__37957),
            .I(N__37945));
    InMux I__3932 (
            .O(N__37956),
            .I(N__37945));
    LocalMux I__3931 (
            .O(N__37953),
            .I(\c0.n13_adj_4785 ));
    LocalMux I__3930 (
            .O(N__37950),
            .I(\c0.n13_adj_4785 ));
    LocalMux I__3929 (
            .O(N__37945),
            .I(\c0.n13_adj_4785 ));
    CascadeMux I__3928 (
            .O(N__37938),
            .I(\c0.n19820_cascade_ ));
    CascadeMux I__3927 (
            .O(N__37935),
            .I(N__37931));
    CascadeMux I__3926 (
            .O(N__37934),
            .I(N__37928));
    InMux I__3925 (
            .O(N__37931),
            .I(N__37922));
    InMux I__3924 (
            .O(N__37928),
            .I(N__37922));
    InMux I__3923 (
            .O(N__37927),
            .I(N__37918));
    LocalMux I__3922 (
            .O(N__37922),
            .I(N__37915));
    InMux I__3921 (
            .O(N__37921),
            .I(N__37912));
    LocalMux I__3920 (
            .O(N__37918),
            .I(N__37907));
    Span4Mux_h I__3919 (
            .O(N__37915),
            .I(N__37907));
    LocalMux I__3918 (
            .O(N__37912),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv4 I__3917 (
            .O(N__37907),
            .I(\c0.FRAME_MATCHER_state_21 ));
    InMux I__3916 (
            .O(N__37902),
            .I(N__37899));
    LocalMux I__3915 (
            .O(N__37899),
            .I(\c0.n27824 ));
    InMux I__3914 (
            .O(N__37896),
            .I(N__37893));
    LocalMux I__3913 (
            .O(N__37893),
            .I(\c0.n16_adj_4797 ));
    CascadeMux I__3912 (
            .O(N__37890),
            .I(\c0.n15_adj_4798_cascade_ ));
    InMux I__3911 (
            .O(N__37887),
            .I(N__37881));
    InMux I__3910 (
            .O(N__37886),
            .I(N__37881));
    LocalMux I__3909 (
            .O(N__37881),
            .I(N__37878));
    Odrv4 I__3908 (
            .O(N__37878),
            .I(\c0.n19546 ));
    CascadeMux I__3907 (
            .O(N__37875),
            .I(N__37869));
    InMux I__3906 (
            .O(N__37874),
            .I(N__37864));
    InMux I__3905 (
            .O(N__37873),
            .I(N__37864));
    InMux I__3904 (
            .O(N__37872),
            .I(N__37859));
    InMux I__3903 (
            .O(N__37869),
            .I(N__37859));
    LocalMux I__3902 (
            .O(N__37864),
            .I(N__37856));
    LocalMux I__3901 (
            .O(N__37859),
            .I(\c0.FRAME_MATCHER_state_30 ));
    Odrv4 I__3900 (
            .O(N__37856),
            .I(\c0.FRAME_MATCHER_state_30 ));
    CascadeMux I__3899 (
            .O(N__37851),
            .I(N__37847));
    InMux I__3898 (
            .O(N__37850),
            .I(N__37842));
    InMux I__3897 (
            .O(N__37847),
            .I(N__37842));
    LocalMux I__3896 (
            .O(N__37842),
            .I(N__37839));
    Span4Mux_v I__3895 (
            .O(N__37839),
            .I(N__37836));
    Span4Mux_h I__3894 (
            .O(N__37836),
            .I(N__37833));
    Odrv4 I__3893 (
            .O(N__37833),
            .I(\c0.n33163 ));
    CascadeMux I__3892 (
            .O(N__37830),
            .I(N__37827));
    InMux I__3891 (
            .O(N__37827),
            .I(N__37824));
    LocalMux I__3890 (
            .O(N__37824),
            .I(N__37818));
    InMux I__3889 (
            .O(N__37823),
            .I(N__37813));
    InMux I__3888 (
            .O(N__37822),
            .I(N__37813));
    InMux I__3887 (
            .O(N__37821),
            .I(N__37810));
    Span4Mux_v I__3886 (
            .O(N__37818),
            .I(N__37805));
    LocalMux I__3885 (
            .O(N__37813),
            .I(N__37805));
    LocalMux I__3884 (
            .O(N__37810),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv4 I__3883 (
            .O(N__37805),
            .I(\c0.FRAME_MATCHER_state_29 ));
    InMux I__3882 (
            .O(N__37800),
            .I(N__37797));
    LocalMux I__3881 (
            .O(N__37797),
            .I(\c0.n12_adj_4789 ));
    InMux I__3880 (
            .O(N__37794),
            .I(N__37791));
    LocalMux I__3879 (
            .O(N__37791),
            .I(\c0.n35771 ));
    CascadeMux I__3878 (
            .O(N__37788),
            .I(\c0.n35698_cascade_ ));
    InMux I__3877 (
            .O(N__37785),
            .I(N__37780));
    InMux I__3876 (
            .O(N__37784),
            .I(N__37777));
    InMux I__3875 (
            .O(N__37783),
            .I(N__37774));
    LocalMux I__3874 (
            .O(N__37780),
            .I(N__37770));
    LocalMux I__3873 (
            .O(N__37777),
            .I(N__37765));
    LocalMux I__3872 (
            .O(N__37774),
            .I(N__37765));
    InMux I__3871 (
            .O(N__37773),
            .I(N__37762));
    Odrv4 I__3870 (
            .O(N__37770),
            .I(data_in_1_2));
    Odrv4 I__3869 (
            .O(N__37765),
            .I(data_in_1_2));
    LocalMux I__3868 (
            .O(N__37762),
            .I(data_in_1_2));
    CascadeMux I__3867 (
            .O(N__37755),
            .I(\c0.n33263_cascade_ ));
    SRMux I__3866 (
            .O(N__37752),
            .I(N__37749));
    LocalMux I__3865 (
            .O(N__37749),
            .I(N__37746));
    Span4Mux_v I__3864 (
            .O(N__37746),
            .I(N__37743));
    Odrv4 I__3863 (
            .O(N__37743),
            .I(\c0.n32718 ));
    CascadeMux I__3862 (
            .O(N__37740),
            .I(\c0.n79_cascade_ ));
    CascadeMux I__3861 (
            .O(N__37737),
            .I(\c0.n4_adj_4613_cascade_ ));
    SRMux I__3860 (
            .O(N__37734),
            .I(N__37731));
    LocalMux I__3859 (
            .O(N__37731),
            .I(N__37728));
    Span4Mux_h I__3858 (
            .O(N__37728),
            .I(N__37725));
    Odrv4 I__3857 (
            .O(N__37725),
            .I(\c0.n8 ));
    CascadeMux I__3856 (
            .O(N__37722),
            .I(\c0.n10_cascade_ ));
    CascadeMux I__3855 (
            .O(N__37719),
            .I(N__37715));
    CascadeMux I__3854 (
            .O(N__37718),
            .I(N__37711));
    InMux I__3853 (
            .O(N__37715),
            .I(N__37705));
    InMux I__3852 (
            .O(N__37714),
            .I(N__37705));
    InMux I__3851 (
            .O(N__37711),
            .I(N__37700));
    InMux I__3850 (
            .O(N__37710),
            .I(N__37700));
    LocalMux I__3849 (
            .O(N__37705),
            .I(\c0.FRAME_MATCHER_state_23 ));
    LocalMux I__3848 (
            .O(N__37700),
            .I(\c0.FRAME_MATCHER_state_23 ));
    InMux I__3847 (
            .O(N__37695),
            .I(N__37689));
    InMux I__3846 (
            .O(N__37694),
            .I(N__37686));
    InMux I__3845 (
            .O(N__37693),
            .I(N__37683));
    InMux I__3844 (
            .O(N__37692),
            .I(N__37680));
    LocalMux I__3843 (
            .O(N__37689),
            .I(\c0.FRAME_MATCHER_state_18 ));
    LocalMux I__3842 (
            .O(N__37686),
            .I(\c0.FRAME_MATCHER_state_18 ));
    LocalMux I__3841 (
            .O(N__37683),
            .I(\c0.FRAME_MATCHER_state_18 ));
    LocalMux I__3840 (
            .O(N__37680),
            .I(\c0.FRAME_MATCHER_state_18 ));
    CascadeMux I__3839 (
            .O(N__37671),
            .I(N__37667));
    InMux I__3838 (
            .O(N__37670),
            .I(N__37660));
    InMux I__3837 (
            .O(N__37667),
            .I(N__37660));
    InMux I__3836 (
            .O(N__37666),
            .I(N__37655));
    InMux I__3835 (
            .O(N__37665),
            .I(N__37655));
    LocalMux I__3834 (
            .O(N__37660),
            .I(\c0.FRAME_MATCHER_state_19 ));
    LocalMux I__3833 (
            .O(N__37655),
            .I(\c0.FRAME_MATCHER_state_19 ));
    CascadeMux I__3832 (
            .O(N__37650),
            .I(N__37643));
    InMux I__3831 (
            .O(N__37649),
            .I(N__37639));
    InMux I__3830 (
            .O(N__37648),
            .I(N__37634));
    InMux I__3829 (
            .O(N__37647),
            .I(N__37634));
    InMux I__3828 (
            .O(N__37646),
            .I(N__37627));
    InMux I__3827 (
            .O(N__37643),
            .I(N__37627));
    InMux I__3826 (
            .O(N__37642),
            .I(N__37627));
    LocalMux I__3825 (
            .O(N__37639),
            .I(N__37624));
    LocalMux I__3824 (
            .O(N__37634),
            .I(r_SM_Main_2_adj_4818));
    LocalMux I__3823 (
            .O(N__37627),
            .I(r_SM_Main_2_adj_4818));
    Odrv4 I__3822 (
            .O(N__37624),
            .I(r_SM_Main_2_adj_4818));
    CascadeMux I__3821 (
            .O(N__37617),
            .I(\c0.tx.n36215_cascade_ ));
    InMux I__3820 (
            .O(N__37614),
            .I(N__37611));
    LocalMux I__3819 (
            .O(N__37611),
            .I(\c0.n36218 ));
    InMux I__3818 (
            .O(N__37608),
            .I(N__37605));
    LocalMux I__3817 (
            .O(N__37605),
            .I(\c0.tx.n19358 ));
    InMux I__3816 (
            .O(N__37602),
            .I(N__37599));
    LocalMux I__3815 (
            .O(N__37599),
            .I(N__37589));
    CascadeMux I__3814 (
            .O(N__37598),
            .I(N__37583));
    InMux I__3813 (
            .O(N__37597),
            .I(N__37575));
    InMux I__3812 (
            .O(N__37596),
            .I(N__37575));
    InMux I__3811 (
            .O(N__37595),
            .I(N__37575));
    InMux I__3810 (
            .O(N__37594),
            .I(N__37572));
    InMux I__3809 (
            .O(N__37593),
            .I(N__37569));
    InMux I__3808 (
            .O(N__37592),
            .I(N__37566));
    Span4Mux_h I__3807 (
            .O(N__37589),
            .I(N__37563));
    InMux I__3806 (
            .O(N__37588),
            .I(N__37558));
    InMux I__3805 (
            .O(N__37587),
            .I(N__37558));
    InMux I__3804 (
            .O(N__37586),
            .I(N__37551));
    InMux I__3803 (
            .O(N__37583),
            .I(N__37551));
    InMux I__3802 (
            .O(N__37582),
            .I(N__37551));
    LocalMux I__3801 (
            .O(N__37575),
            .I(N__37548));
    LocalMux I__3800 (
            .O(N__37572),
            .I(r_SM_Main_1_adj_4819));
    LocalMux I__3799 (
            .O(N__37569),
            .I(r_SM_Main_1_adj_4819));
    LocalMux I__3798 (
            .O(N__37566),
            .I(r_SM_Main_1_adj_4819));
    Odrv4 I__3797 (
            .O(N__37563),
            .I(r_SM_Main_1_adj_4819));
    LocalMux I__3796 (
            .O(N__37558),
            .I(r_SM_Main_1_adj_4819));
    LocalMux I__3795 (
            .O(N__37551),
            .I(r_SM_Main_1_adj_4819));
    Odrv4 I__3794 (
            .O(N__37548),
            .I(r_SM_Main_1_adj_4819));
    InMux I__3793 (
            .O(N__37533),
            .I(N__37530));
    LocalMux I__3792 (
            .O(N__37530),
            .I(n35927));
    CEMux I__3791 (
            .O(N__37527),
            .I(N__37523));
    CEMux I__3790 (
            .O(N__37526),
            .I(N__37519));
    LocalMux I__3789 (
            .O(N__37523),
            .I(N__37516));
    InMux I__3788 (
            .O(N__37522),
            .I(N__37513));
    LocalMux I__3787 (
            .O(N__37519),
            .I(N__37505));
    Span4Mux_v I__3786 (
            .O(N__37516),
            .I(N__37505));
    LocalMux I__3785 (
            .O(N__37513),
            .I(N__37505));
    InMux I__3784 (
            .O(N__37512),
            .I(N__37502));
    Span4Mux_v I__3783 (
            .O(N__37505),
            .I(N__37498));
    LocalMux I__3782 (
            .O(N__37502),
            .I(N__37495));
    InMux I__3781 (
            .O(N__37501),
            .I(N__37492));
    Odrv4 I__3780 (
            .O(N__37498),
            .I(n19509));
    Odrv4 I__3779 (
            .O(N__37495),
            .I(n19509));
    LocalMux I__3778 (
            .O(N__37492),
            .I(n19509));
    CascadeMux I__3777 (
            .O(N__37485),
            .I(n9_cascade_));
    InMux I__3776 (
            .O(N__37482),
            .I(N__37476));
    CascadeMux I__3775 (
            .O(N__37481),
            .I(N__37473));
    CascadeMux I__3774 (
            .O(N__37480),
            .I(N__37470));
    InMux I__3773 (
            .O(N__37479),
            .I(N__37465));
    LocalMux I__3772 (
            .O(N__37476),
            .I(N__37462));
    InMux I__3771 (
            .O(N__37473),
            .I(N__37459));
    InMux I__3770 (
            .O(N__37470),
            .I(N__37452));
    InMux I__3769 (
            .O(N__37469),
            .I(N__37452));
    InMux I__3768 (
            .O(N__37468),
            .I(N__37452));
    LocalMux I__3767 (
            .O(N__37465),
            .I(n22210));
    Odrv4 I__3766 (
            .O(N__37462),
            .I(n22210));
    LocalMux I__3765 (
            .O(N__37459),
            .I(n22210));
    LocalMux I__3764 (
            .O(N__37452),
            .I(n22210));
    InMux I__3763 (
            .O(N__37443),
            .I(N__37440));
    LocalMux I__3762 (
            .O(N__37440),
            .I(N__37431));
    InMux I__3761 (
            .O(N__37439),
            .I(N__37423));
    InMux I__3760 (
            .O(N__37438),
            .I(N__37423));
    InMux I__3759 (
            .O(N__37437),
            .I(N__37423));
    InMux I__3758 (
            .O(N__37436),
            .I(N__37418));
    InMux I__3757 (
            .O(N__37435),
            .I(N__37418));
    InMux I__3756 (
            .O(N__37434),
            .I(N__37414));
    Span4Mux_h I__3755 (
            .O(N__37431),
            .I(N__37411));
    InMux I__3754 (
            .O(N__37430),
            .I(N__37408));
    LocalMux I__3753 (
            .O(N__37423),
            .I(N__37403));
    LocalMux I__3752 (
            .O(N__37418),
            .I(N__37403));
    InMux I__3751 (
            .O(N__37417),
            .I(N__37400));
    LocalMux I__3750 (
            .O(N__37414),
            .I(r_SM_Main_0));
    Odrv4 I__3749 (
            .O(N__37411),
            .I(r_SM_Main_0));
    LocalMux I__3748 (
            .O(N__37408),
            .I(r_SM_Main_0));
    Odrv4 I__3747 (
            .O(N__37403),
            .I(r_SM_Main_0));
    LocalMux I__3746 (
            .O(N__37400),
            .I(r_SM_Main_0));
    InMux I__3745 (
            .O(N__37389),
            .I(N__37386));
    LocalMux I__3744 (
            .O(N__37386),
            .I(N__37381));
    InMux I__3743 (
            .O(N__37385),
            .I(N__37378));
    InMux I__3742 (
            .O(N__37384),
            .I(N__37375));
    Span4Mux_h I__3741 (
            .O(N__37381),
            .I(N__37372));
    LocalMux I__3740 (
            .O(N__37378),
            .I(\c0.FRAME_MATCHER_state_27 ));
    LocalMux I__3739 (
            .O(N__37375),
            .I(\c0.FRAME_MATCHER_state_27 ));
    Odrv4 I__3738 (
            .O(N__37372),
            .I(\c0.FRAME_MATCHER_state_27 ));
    CascadeMux I__3737 (
            .O(N__37365),
            .I(N__37361));
    InMux I__3736 (
            .O(N__37364),
            .I(N__37357));
    InMux I__3735 (
            .O(N__37361),
            .I(N__37352));
    InMux I__3734 (
            .O(N__37360),
            .I(N__37352));
    LocalMux I__3733 (
            .O(N__37357),
            .I(\c0.FRAME_MATCHER_state_31 ));
    LocalMux I__3732 (
            .O(N__37352),
            .I(\c0.FRAME_MATCHER_state_31 ));
    InMux I__3731 (
            .O(N__37347),
            .I(N__37343));
    InMux I__3730 (
            .O(N__37346),
            .I(N__37340));
    LocalMux I__3729 (
            .O(N__37343),
            .I(\quad_counter0.a_delay_counter_13 ));
    LocalMux I__3728 (
            .O(N__37340),
            .I(\quad_counter0.a_delay_counter_13 ));
    InMux I__3727 (
            .O(N__37335),
            .I(N__37331));
    InMux I__3726 (
            .O(N__37334),
            .I(N__37328));
    LocalMux I__3725 (
            .O(N__37331),
            .I(\quad_counter0.a_delay_counter_9 ));
    LocalMux I__3724 (
            .O(N__37328),
            .I(\quad_counter0.a_delay_counter_9 ));
    CascadeMux I__3723 (
            .O(N__37323),
            .I(N__37320));
    InMux I__3722 (
            .O(N__37320),
            .I(N__37316));
    InMux I__3721 (
            .O(N__37319),
            .I(N__37313));
    LocalMux I__3720 (
            .O(N__37316),
            .I(N__37310));
    LocalMux I__3719 (
            .O(N__37313),
            .I(\quad_counter0.a_delay_counter_6 ));
    Odrv4 I__3718 (
            .O(N__37310),
            .I(\quad_counter0.a_delay_counter_6 ));
    InMux I__3717 (
            .O(N__37305),
            .I(N__37301));
    InMux I__3716 (
            .O(N__37304),
            .I(N__37298));
    LocalMux I__3715 (
            .O(N__37301),
            .I(\quad_counter0.a_delay_counter_12 ));
    LocalMux I__3714 (
            .O(N__37298),
            .I(\quad_counter0.a_delay_counter_12 ));
    InMux I__3713 (
            .O(N__37293),
            .I(N__37290));
    LocalMux I__3712 (
            .O(N__37290),
            .I(N__37287));
    Odrv4 I__3711 (
            .O(N__37287),
            .I(\quad_counter0.n28_adj_4410 ));
    InMux I__3710 (
            .O(N__37284),
            .I(N__37281));
    LocalMux I__3709 (
            .O(N__37281),
            .I(\quad_counter0.n27_adj_4412 ));
    CascadeMux I__3708 (
            .O(N__37278),
            .I(\quad_counter0.n26_adj_4411_cascade_ ));
    InMux I__3707 (
            .O(N__37275),
            .I(N__37272));
    LocalMux I__3706 (
            .O(N__37272),
            .I(N__37269));
    Odrv4 I__3705 (
            .O(N__37269),
            .I(\quad_counter0.n25_adj_4413 ));
    CascadeMux I__3704 (
            .O(N__37266),
            .I(\c0.tx.n4_cascade_ ));
    InMux I__3703 (
            .O(N__37263),
            .I(N__37260));
    LocalMux I__3702 (
            .O(N__37260),
            .I(\c0.tx.n22211 ));
    InMux I__3701 (
            .O(N__37257),
            .I(N__37252));
    CEMux I__3700 (
            .O(N__37256),
            .I(N__37249));
    CEMux I__3699 (
            .O(N__37255),
            .I(N__37246));
    LocalMux I__3698 (
            .O(N__37252),
            .I(N__37243));
    LocalMux I__3697 (
            .O(N__37249),
            .I(N__37240));
    LocalMux I__3696 (
            .O(N__37246),
            .I(N__37237));
    Span4Mux_v I__3695 (
            .O(N__37243),
            .I(N__37234));
    Sp12to4 I__3694 (
            .O(N__37240),
            .I(N__37231));
    Odrv4 I__3693 (
            .O(N__37237),
            .I(n19493));
    Odrv4 I__3692 (
            .O(N__37234),
            .I(n19493));
    Odrv12 I__3691 (
            .O(N__37231),
            .I(n19493));
    InMux I__3690 (
            .O(N__37224),
            .I(N__37218));
    InMux I__3689 (
            .O(N__37223),
            .I(N__37218));
    LocalMux I__3688 (
            .O(N__37218),
            .I(N__37215));
    Span4Mux_h I__3687 (
            .O(N__37215),
            .I(N__37210));
    InMux I__3686 (
            .O(N__37214),
            .I(N__37207));
    InMux I__3685 (
            .O(N__37213),
            .I(N__37204));
    Span4Mux_h I__3684 (
            .O(N__37210),
            .I(N__37199));
    LocalMux I__3683 (
            .O(N__37207),
            .I(N__37199));
    LocalMux I__3682 (
            .O(N__37204),
            .I(N__37196));
    Span4Mux_v I__3681 (
            .O(N__37199),
            .I(N__37193));
    Span12Mux_v I__3680 (
            .O(N__37196),
            .I(N__37190));
    Span4Mux_v I__3679 (
            .O(N__37193),
            .I(N__37187));
    Odrv12 I__3678 (
            .O(N__37190),
            .I(PIN_7_c));
    Odrv4 I__3677 (
            .O(N__37187),
            .I(PIN_7_c));
    InMux I__3676 (
            .O(N__37182),
            .I(N__37176));
    InMux I__3675 (
            .O(N__37181),
            .I(N__37176));
    LocalMux I__3674 (
            .O(N__37176),
            .I(n15010));
    InMux I__3673 (
            .O(N__37173),
            .I(N__37167));
    InMux I__3672 (
            .O(N__37172),
            .I(N__37167));
    LocalMux I__3671 (
            .O(N__37167),
            .I(N__37163));
    InMux I__3670 (
            .O(N__37166),
            .I(N__37160));
    Span4Mux_v I__3669 (
            .O(N__37163),
            .I(N__37155));
    LocalMux I__3668 (
            .O(N__37160),
            .I(N__37155));
    Span4Mux_h I__3667 (
            .O(N__37155),
            .I(N__37152));
    Span4Mux_v I__3666 (
            .O(N__37152),
            .I(N__37149));
    Odrv4 I__3665 (
            .O(N__37149),
            .I(quadA_delayed));
    InMux I__3664 (
            .O(N__37146),
            .I(\quad_counter0.n30025 ));
    InMux I__3663 (
            .O(N__37143),
            .I(N__37139));
    InMux I__3662 (
            .O(N__37142),
            .I(N__37136));
    LocalMux I__3661 (
            .O(N__37139),
            .I(\quad_counter0.a_delay_counter_11 ));
    LocalMux I__3660 (
            .O(N__37136),
            .I(\quad_counter0.a_delay_counter_11 ));
    InMux I__3659 (
            .O(N__37131),
            .I(\quad_counter0.n30026 ));
    InMux I__3658 (
            .O(N__37128),
            .I(\quad_counter0.n30027 ));
    InMux I__3657 (
            .O(N__37125),
            .I(\quad_counter0.n30028 ));
    InMux I__3656 (
            .O(N__37122),
            .I(\quad_counter0.n30029 ));
    InMux I__3655 (
            .O(N__37119),
            .I(\quad_counter0.n30030 ));
    SRMux I__3654 (
            .O(N__37116),
            .I(N__37112));
    SRMux I__3653 (
            .O(N__37115),
            .I(N__37109));
    LocalMux I__3652 (
            .O(N__37112),
            .I(N__37106));
    LocalMux I__3651 (
            .O(N__37109),
            .I(N__37103));
    Span4Mux_h I__3650 (
            .O(N__37106),
            .I(N__37100));
    Span4Mux_h I__3649 (
            .O(N__37103),
            .I(N__37097));
    Odrv4 I__3648 (
            .O(N__37100),
            .I(a_delay_counter_15__N_4220));
    Odrv4 I__3647 (
            .O(N__37097),
            .I(a_delay_counter_15__N_4220));
    CascadeMux I__3646 (
            .O(N__37092),
            .I(N__37086));
    InMux I__3645 (
            .O(N__37091),
            .I(N__37083));
    InMux I__3644 (
            .O(N__37090),
            .I(N__37080));
    InMux I__3643 (
            .O(N__37089),
            .I(N__37075));
    InMux I__3642 (
            .O(N__37086),
            .I(N__37075));
    LocalMux I__3641 (
            .O(N__37083),
            .I(\c0.n19530 ));
    LocalMux I__3640 (
            .O(N__37080),
            .I(\c0.n19530 ));
    LocalMux I__3639 (
            .O(N__37075),
            .I(\c0.n19530 ));
    InMux I__3638 (
            .O(N__37068),
            .I(N__37064));
    InMux I__3637 (
            .O(N__37067),
            .I(N__37061));
    LocalMux I__3636 (
            .O(N__37064),
            .I(\quad_counter0.a_delay_counter_10 ));
    LocalMux I__3635 (
            .O(N__37061),
            .I(\quad_counter0.a_delay_counter_10 ));
    InMux I__3634 (
            .O(N__37056),
            .I(N__37052));
    InMux I__3633 (
            .O(N__37055),
            .I(N__37049));
    LocalMux I__3632 (
            .O(N__37052),
            .I(\quad_counter0.a_delay_counter_14 ));
    LocalMux I__3631 (
            .O(N__37049),
            .I(\quad_counter0.a_delay_counter_14 ));
    CascadeMux I__3630 (
            .O(N__37044),
            .I(N__37040));
    InMux I__3629 (
            .O(N__37043),
            .I(N__37037));
    InMux I__3628 (
            .O(N__37040),
            .I(N__37034));
    LocalMux I__3627 (
            .O(N__37037),
            .I(\quad_counter0.a_delay_counter_15 ));
    LocalMux I__3626 (
            .O(N__37034),
            .I(\quad_counter0.a_delay_counter_15 ));
    InMux I__3625 (
            .O(N__37029),
            .I(N__37025));
    InMux I__3624 (
            .O(N__37028),
            .I(N__37022));
    LocalMux I__3623 (
            .O(N__37025),
            .I(N__37019));
    LocalMux I__3622 (
            .O(N__37022),
            .I(\quad_counter0.a_delay_counter_7 ));
    Odrv4 I__3621 (
            .O(N__37019),
            .I(\quad_counter0.a_delay_counter_7 ));
    InMux I__3620 (
            .O(N__37014),
            .I(N__37010));
    InMux I__3619 (
            .O(N__37013),
            .I(N__37007));
    LocalMux I__3618 (
            .O(N__37010),
            .I(\quad_counter0.a_delay_counter_1 ));
    LocalMux I__3617 (
            .O(N__37007),
            .I(\quad_counter0.a_delay_counter_1 ));
    InMux I__3616 (
            .O(N__37002),
            .I(\quad_counter0.n30016 ));
    CascadeMux I__3615 (
            .O(N__36999),
            .I(N__36995));
    InMux I__3614 (
            .O(N__36998),
            .I(N__36992));
    InMux I__3613 (
            .O(N__36995),
            .I(N__36989));
    LocalMux I__3612 (
            .O(N__36992),
            .I(\quad_counter0.a_delay_counter_2 ));
    LocalMux I__3611 (
            .O(N__36989),
            .I(\quad_counter0.a_delay_counter_2 ));
    InMux I__3610 (
            .O(N__36984),
            .I(\quad_counter0.n30017 ));
    InMux I__3609 (
            .O(N__36981),
            .I(N__36977));
    InMux I__3608 (
            .O(N__36980),
            .I(N__36974));
    LocalMux I__3607 (
            .O(N__36977),
            .I(\quad_counter0.a_delay_counter_3 ));
    LocalMux I__3606 (
            .O(N__36974),
            .I(\quad_counter0.a_delay_counter_3 ));
    InMux I__3605 (
            .O(N__36969),
            .I(\quad_counter0.n30018 ));
    CascadeMux I__3604 (
            .O(N__36966),
            .I(N__36962));
    InMux I__3603 (
            .O(N__36965),
            .I(N__36959));
    InMux I__3602 (
            .O(N__36962),
            .I(N__36956));
    LocalMux I__3601 (
            .O(N__36959),
            .I(\quad_counter0.a_delay_counter_4 ));
    LocalMux I__3600 (
            .O(N__36956),
            .I(\quad_counter0.a_delay_counter_4 ));
    InMux I__3599 (
            .O(N__36951),
            .I(\quad_counter0.n30019 ));
    InMux I__3598 (
            .O(N__36948),
            .I(N__36944));
    InMux I__3597 (
            .O(N__36947),
            .I(N__36941));
    LocalMux I__3596 (
            .O(N__36944),
            .I(\quad_counter0.a_delay_counter_5 ));
    LocalMux I__3595 (
            .O(N__36941),
            .I(\quad_counter0.a_delay_counter_5 ));
    InMux I__3594 (
            .O(N__36936),
            .I(\quad_counter0.n30020 ));
    InMux I__3593 (
            .O(N__36933),
            .I(\quad_counter0.n30021 ));
    InMux I__3592 (
            .O(N__36930),
            .I(\quad_counter0.n30022 ));
    InMux I__3591 (
            .O(N__36927),
            .I(N__36923));
    InMux I__3590 (
            .O(N__36926),
            .I(N__36920));
    LocalMux I__3589 (
            .O(N__36923),
            .I(\quad_counter0.a_delay_counter_8 ));
    LocalMux I__3588 (
            .O(N__36920),
            .I(\quad_counter0.a_delay_counter_8 ));
    InMux I__3587 (
            .O(N__36915),
            .I(bfn_7_10_0_));
    InMux I__3586 (
            .O(N__36912),
            .I(\quad_counter0.n30024 ));
    InMux I__3585 (
            .O(N__36909),
            .I(N__36906));
    LocalMux I__3584 (
            .O(N__36906),
            .I(N__36902));
    InMux I__3583 (
            .O(N__36905),
            .I(N__36899));
    Span4Mux_v I__3582 (
            .O(N__36902),
            .I(N__36896));
    LocalMux I__3581 (
            .O(N__36899),
            .I(n27744));
    Odrv4 I__3580 (
            .O(N__36896),
            .I(n27744));
    InMux I__3579 (
            .O(N__36891),
            .I(N__36887));
    InMux I__3578 (
            .O(N__36890),
            .I(N__36884));
    LocalMux I__3577 (
            .O(N__36887),
            .I(n4_adj_4808));
    LocalMux I__3576 (
            .O(N__36884),
            .I(n4_adj_4808));
    InMux I__3575 (
            .O(N__36879),
            .I(N__36874));
    InMux I__3574 (
            .O(N__36878),
            .I(N__36869));
    InMux I__3573 (
            .O(N__36877),
            .I(N__36869));
    LocalMux I__3572 (
            .O(N__36874),
            .I(a_delay_counter_0));
    LocalMux I__3571 (
            .O(N__36869),
            .I(a_delay_counter_0));
    InMux I__3570 (
            .O(N__36864),
            .I(N__36861));
    LocalMux I__3569 (
            .O(N__36861),
            .I(n39));
    InMux I__3568 (
            .O(N__36858),
            .I(bfn_7_9_0_));
    InMux I__3567 (
            .O(N__36855),
            .I(N__36851));
    InMux I__3566 (
            .O(N__36854),
            .I(N__36848));
    LocalMux I__3565 (
            .O(N__36851),
            .I(data_in_0_0));
    LocalMux I__3564 (
            .O(N__36848),
            .I(data_in_0_0));
    InMux I__3563 (
            .O(N__36843),
            .I(N__36835));
    InMux I__3562 (
            .O(N__36842),
            .I(N__36835));
    InMux I__3561 (
            .O(N__36841),
            .I(N__36830));
    InMux I__3560 (
            .O(N__36840),
            .I(N__36830));
    LocalMux I__3559 (
            .O(N__36835),
            .I(data_in_1_0));
    LocalMux I__3558 (
            .O(N__36830),
            .I(data_in_1_0));
    CascadeMux I__3557 (
            .O(N__36825),
            .I(N__36821));
    InMux I__3556 (
            .O(N__36824),
            .I(N__36815));
    InMux I__3555 (
            .O(N__36821),
            .I(N__36815));
    InMux I__3554 (
            .O(N__36820),
            .I(N__36812));
    LocalMux I__3553 (
            .O(N__36815),
            .I(N__36809));
    LocalMux I__3552 (
            .O(N__36812),
            .I(data_in_0_3));
    Odrv4 I__3551 (
            .O(N__36809),
            .I(data_in_0_3));
    CascadeMux I__3550 (
            .O(N__36804),
            .I(N__36800));
    InMux I__3549 (
            .O(N__36803),
            .I(N__36793));
    InMux I__3548 (
            .O(N__36800),
            .I(N__36793));
    InMux I__3547 (
            .O(N__36799),
            .I(N__36790));
    InMux I__3546 (
            .O(N__36798),
            .I(N__36787));
    LocalMux I__3545 (
            .O(N__36793),
            .I(N__36784));
    LocalMux I__3544 (
            .O(N__36790),
            .I(data_in_2_4));
    LocalMux I__3543 (
            .O(N__36787),
            .I(data_in_2_4));
    Odrv4 I__3542 (
            .O(N__36784),
            .I(data_in_2_4));
    CascadeMux I__3541 (
            .O(N__36777),
            .I(N__36774));
    InMux I__3540 (
            .O(N__36774),
            .I(N__36770));
    InMux I__3539 (
            .O(N__36773),
            .I(N__36766));
    LocalMux I__3538 (
            .O(N__36770),
            .I(N__36763));
    CascadeMux I__3537 (
            .O(N__36769),
            .I(N__36759));
    LocalMux I__3536 (
            .O(N__36766),
            .I(N__36756));
    Span4Mux_v I__3535 (
            .O(N__36763),
            .I(N__36753));
    InMux I__3534 (
            .O(N__36762),
            .I(N__36748));
    InMux I__3533 (
            .O(N__36759),
            .I(N__36748));
    Odrv4 I__3532 (
            .O(N__36756),
            .I(data_in_2_1));
    Odrv4 I__3531 (
            .O(N__36753),
            .I(data_in_2_1));
    LocalMux I__3530 (
            .O(N__36748),
            .I(data_in_2_1));
    InMux I__3529 (
            .O(N__36741),
            .I(N__36736));
    InMux I__3528 (
            .O(N__36740),
            .I(N__36733));
    InMux I__3527 (
            .O(N__36739),
            .I(N__36730));
    LocalMux I__3526 (
            .O(N__36736),
            .I(data_in_1_1));
    LocalMux I__3525 (
            .O(N__36733),
            .I(data_in_1_1));
    LocalMux I__3524 (
            .O(N__36730),
            .I(data_in_1_1));
    CascadeMux I__3523 (
            .O(N__36723),
            .I(N__36718));
    InMux I__3522 (
            .O(N__36722),
            .I(N__36715));
    InMux I__3521 (
            .O(N__36721),
            .I(N__36710));
    InMux I__3520 (
            .O(N__36718),
            .I(N__36710));
    LocalMux I__3519 (
            .O(N__36715),
            .I(data_in_0_5));
    LocalMux I__3518 (
            .O(N__36710),
            .I(data_in_0_5));
    InMux I__3517 (
            .O(N__36705),
            .I(N__36699));
    InMux I__3516 (
            .O(N__36704),
            .I(N__36696));
    InMux I__3515 (
            .O(N__36703),
            .I(N__36691));
    InMux I__3514 (
            .O(N__36702),
            .I(N__36691));
    LocalMux I__3513 (
            .O(N__36699),
            .I(data_in_1_6));
    LocalMux I__3512 (
            .O(N__36696),
            .I(data_in_1_6));
    LocalMux I__3511 (
            .O(N__36691),
            .I(data_in_1_6));
    InMux I__3510 (
            .O(N__36684),
            .I(N__36676));
    InMux I__3509 (
            .O(N__36683),
            .I(N__36676));
    InMux I__3508 (
            .O(N__36682),
            .I(N__36671));
    InMux I__3507 (
            .O(N__36681),
            .I(N__36671));
    LocalMux I__3506 (
            .O(N__36676),
            .I(N__36668));
    LocalMux I__3505 (
            .O(N__36671),
            .I(data_in_3_7));
    Odrv4 I__3504 (
            .O(N__36668),
            .I(data_in_3_7));
    CascadeMux I__3503 (
            .O(N__36663),
            .I(\c0.n17_adj_4791_cascade_ ));
    InMux I__3502 (
            .O(N__36660),
            .I(N__36657));
    LocalMux I__3501 (
            .O(N__36657),
            .I(\c0.n16_adj_4790 ));
    CascadeMux I__3500 (
            .O(N__36654),
            .I(N__36650));
    InMux I__3499 (
            .O(N__36653),
            .I(N__36647));
    InMux I__3498 (
            .O(N__36650),
            .I(N__36644));
    LocalMux I__3497 (
            .O(N__36647),
            .I(\c0.n18094 ));
    LocalMux I__3496 (
            .O(N__36644),
            .I(\c0.n18094 ));
    InMux I__3495 (
            .O(N__36639),
            .I(N__36633));
    InMux I__3494 (
            .O(N__36638),
            .I(N__36630));
    InMux I__3493 (
            .O(N__36637),
            .I(N__36627));
    InMux I__3492 (
            .O(N__36636),
            .I(N__36624));
    LocalMux I__3491 (
            .O(N__36633),
            .I(N__36619));
    LocalMux I__3490 (
            .O(N__36630),
            .I(N__36619));
    LocalMux I__3489 (
            .O(N__36627),
            .I(data_in_1_5));
    LocalMux I__3488 (
            .O(N__36624),
            .I(data_in_1_5));
    Odrv4 I__3487 (
            .O(N__36619),
            .I(data_in_1_5));
    InMux I__3486 (
            .O(N__36612),
            .I(N__36609));
    LocalMux I__3485 (
            .O(N__36609),
            .I(N__36605));
    InMux I__3484 (
            .O(N__36608),
            .I(N__36602));
    Span4Mux_v I__3483 (
            .O(N__36605),
            .I(N__36596));
    LocalMux I__3482 (
            .O(N__36602),
            .I(N__36596));
    InMux I__3481 (
            .O(N__36601),
            .I(N__36593));
    Span4Mux_v I__3480 (
            .O(N__36596),
            .I(N__36590));
    LocalMux I__3479 (
            .O(N__36593),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__3478 (
            .O(N__36590),
            .I(\c0.FRAME_MATCHER_state_9 ));
    SRMux I__3477 (
            .O(N__36585),
            .I(N__36582));
    LocalMux I__3476 (
            .O(N__36582),
            .I(N__36579));
    Span4Mux_h I__3475 (
            .O(N__36579),
            .I(N__36576));
    Span4Mux_v I__3474 (
            .O(N__36576),
            .I(N__36573));
    Odrv4 I__3473 (
            .O(N__36573),
            .I(\c0.n8_adj_4496 ));
    SRMux I__3472 (
            .O(N__36570),
            .I(N__36567));
    LocalMux I__3471 (
            .O(N__36567),
            .I(\c0.n32798 ));
    CascadeMux I__3470 (
            .O(N__36564),
            .I(N__36559));
    InMux I__3469 (
            .O(N__36563),
            .I(N__36556));
    InMux I__3468 (
            .O(N__36562),
            .I(N__36550));
    InMux I__3467 (
            .O(N__36559),
            .I(N__36550));
    LocalMux I__3466 (
            .O(N__36556),
            .I(N__36547));
    InMux I__3465 (
            .O(N__36555),
            .I(N__36544));
    LocalMux I__3464 (
            .O(N__36550),
            .I(N__36541));
    Odrv4 I__3463 (
            .O(N__36547),
            .I(data_in_1_4));
    LocalMux I__3462 (
            .O(N__36544),
            .I(data_in_1_4));
    Odrv4 I__3461 (
            .O(N__36541),
            .I(data_in_1_4));
    CascadeMux I__3460 (
            .O(N__36534),
            .I(N__36531));
    InMux I__3459 (
            .O(N__36531),
            .I(N__36527));
    InMux I__3458 (
            .O(N__36530),
            .I(N__36524));
    LocalMux I__3457 (
            .O(N__36527),
            .I(N__36521));
    LocalMux I__3456 (
            .O(N__36524),
            .I(data_in_0_4));
    Odrv4 I__3455 (
            .O(N__36521),
            .I(data_in_0_4));
    InMux I__3454 (
            .O(N__36516),
            .I(N__36510));
    InMux I__3453 (
            .O(N__36515),
            .I(N__36510));
    LocalMux I__3452 (
            .O(N__36510),
            .I(N__36506));
    InMux I__3451 (
            .O(N__36509),
            .I(N__36503));
    Span4Mux_h I__3450 (
            .O(N__36506),
            .I(N__36500));
    LocalMux I__3449 (
            .O(N__36503),
            .I(data_in_0_1));
    Odrv4 I__3448 (
            .O(N__36500),
            .I(data_in_0_1));
    InMux I__3447 (
            .O(N__36495),
            .I(N__36490));
    InMux I__3446 (
            .O(N__36494),
            .I(N__36487));
    InMux I__3445 (
            .O(N__36493),
            .I(N__36484));
    LocalMux I__3444 (
            .O(N__36490),
            .I(N__36479));
    LocalMux I__3443 (
            .O(N__36487),
            .I(N__36479));
    LocalMux I__3442 (
            .O(N__36484),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv12 I__3441 (
            .O(N__36479),
            .I(\c0.FRAME_MATCHER_state_14 ));
    CascadeMux I__3440 (
            .O(N__36474),
            .I(N__36471));
    InMux I__3439 (
            .O(N__36471),
            .I(N__36467));
    CascadeMux I__3438 (
            .O(N__36470),
            .I(N__36463));
    LocalMux I__3437 (
            .O(N__36467),
            .I(N__36460));
    InMux I__3436 (
            .O(N__36466),
            .I(N__36457));
    InMux I__3435 (
            .O(N__36463),
            .I(N__36454));
    Span4Mux_h I__3434 (
            .O(N__36460),
            .I(N__36451));
    LocalMux I__3433 (
            .O(N__36457),
            .I(\c0.FRAME_MATCHER_state_15 ));
    LocalMux I__3432 (
            .O(N__36454),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__3431 (
            .O(N__36451),
            .I(\c0.FRAME_MATCHER_state_15 ));
    InMux I__3430 (
            .O(N__36444),
            .I(N__36439));
    InMux I__3429 (
            .O(N__36443),
            .I(N__36436));
    InMux I__3428 (
            .O(N__36442),
            .I(N__36433));
    LocalMux I__3427 (
            .O(N__36439),
            .I(\c0.FRAME_MATCHER_state_11 ));
    LocalMux I__3426 (
            .O(N__36436),
            .I(\c0.FRAME_MATCHER_state_11 ));
    LocalMux I__3425 (
            .O(N__36433),
            .I(\c0.FRAME_MATCHER_state_11 ));
    InMux I__3424 (
            .O(N__36426),
            .I(N__36423));
    LocalMux I__3423 (
            .O(N__36423),
            .I(\c0.n16_adj_4787 ));
    InMux I__3422 (
            .O(N__36420),
            .I(N__36415));
    InMux I__3421 (
            .O(N__36419),
            .I(N__36410));
    InMux I__3420 (
            .O(N__36418),
            .I(N__36410));
    LocalMux I__3419 (
            .O(N__36415),
            .I(\c0.FRAME_MATCHER_state_7 ));
    LocalMux I__3418 (
            .O(N__36410),
            .I(\c0.FRAME_MATCHER_state_7 ));
    SRMux I__3417 (
            .O(N__36405),
            .I(N__36402));
    LocalMux I__3416 (
            .O(N__36402),
            .I(\c0.n32840 ));
    InMux I__3415 (
            .O(N__36399),
            .I(N__36395));
    InMux I__3414 (
            .O(N__36398),
            .I(N__36391));
    LocalMux I__3413 (
            .O(N__36395),
            .I(N__36388));
    InMux I__3412 (
            .O(N__36394),
            .I(N__36385));
    LocalMux I__3411 (
            .O(N__36391),
            .I(\c0.FRAME_MATCHER_state_22 ));
    Odrv12 I__3410 (
            .O(N__36388),
            .I(\c0.FRAME_MATCHER_state_22 ));
    LocalMux I__3409 (
            .O(N__36385),
            .I(\c0.FRAME_MATCHER_state_22 ));
    CascadeMux I__3408 (
            .O(N__36378),
            .I(\c0.n45_adj_4637_cascade_ ));
    SRMux I__3407 (
            .O(N__36375),
            .I(N__36372));
    LocalMux I__3406 (
            .O(N__36372),
            .I(N__36369));
    Odrv12 I__3405 (
            .O(N__36369),
            .I(\c0.n32714 ));
    CascadeMux I__3404 (
            .O(N__36366),
            .I(N__36363));
    InMux I__3403 (
            .O(N__36363),
            .I(N__36359));
    InMux I__3402 (
            .O(N__36362),
            .I(N__36355));
    LocalMux I__3401 (
            .O(N__36359),
            .I(N__36352));
    InMux I__3400 (
            .O(N__36358),
            .I(N__36349));
    LocalMux I__3399 (
            .O(N__36355),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv12 I__3398 (
            .O(N__36352),
            .I(\c0.FRAME_MATCHER_state_20 ));
    LocalMux I__3397 (
            .O(N__36349),
            .I(\c0.FRAME_MATCHER_state_20 ));
    SRMux I__3396 (
            .O(N__36342),
            .I(N__36339));
    LocalMux I__3395 (
            .O(N__36339),
            .I(N__36336));
    Span4Mux_h I__3394 (
            .O(N__36336),
            .I(N__36333));
    Odrv4 I__3393 (
            .O(N__36333),
            .I(\c0.n32804 ));
    SRMux I__3392 (
            .O(N__36330),
            .I(N__36327));
    LocalMux I__3391 (
            .O(N__36327),
            .I(N__36324));
    Odrv4 I__3390 (
            .O(N__36324),
            .I(\c0.n32712 ));
    InMux I__3389 (
            .O(N__36321),
            .I(N__36317));
    InMux I__3388 (
            .O(N__36320),
            .I(N__36314));
    LocalMux I__3387 (
            .O(N__36317),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__3386 (
            .O(N__36314),
            .I(\c0.tx.r_Clock_Count_5 ));
    InMux I__3385 (
            .O(N__36309),
            .I(N__36305));
    InMux I__3384 (
            .O(N__36308),
            .I(N__36302));
    LocalMux I__3383 (
            .O(N__36305),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__3382 (
            .O(N__36302),
            .I(\c0.tx.r_Clock_Count_7 ));
    CascadeMux I__3381 (
            .O(N__36297),
            .I(N__36293));
    InMux I__3380 (
            .O(N__36296),
            .I(N__36290));
    InMux I__3379 (
            .O(N__36293),
            .I(N__36287));
    LocalMux I__3378 (
            .O(N__36290),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__3377 (
            .O(N__36287),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__3376 (
            .O(N__36282),
            .I(N__36278));
    InMux I__3375 (
            .O(N__36281),
            .I(N__36275));
    LocalMux I__3374 (
            .O(N__36278),
            .I(\c0.tx.r_Clock_Count_8 ));
    LocalMux I__3373 (
            .O(N__36275),
            .I(\c0.tx.r_Clock_Count_8 ));
    InMux I__3372 (
            .O(N__36270),
            .I(N__36267));
    LocalMux I__3371 (
            .O(N__36267),
            .I(\c0.n47_adj_4651 ));
    CascadeMux I__3370 (
            .O(N__36264),
            .I(\c0.n10_adj_4504_cascade_ ));
    InMux I__3369 (
            .O(N__36261),
            .I(N__36258));
    LocalMux I__3368 (
            .O(N__36258),
            .I(N__36255));
    Odrv4 I__3367 (
            .O(N__36255),
            .I(\c0.n35 ));
    InMux I__3366 (
            .O(N__36252),
            .I(N__36240));
    InMux I__3365 (
            .O(N__36251),
            .I(N__36240));
    InMux I__3364 (
            .O(N__36250),
            .I(N__36240));
    InMux I__3363 (
            .O(N__36249),
            .I(N__36240));
    LocalMux I__3362 (
            .O(N__36240),
            .I(r_Bit_Index_2));
    SRMux I__3361 (
            .O(N__36237),
            .I(N__36234));
    LocalMux I__3360 (
            .O(N__36234),
            .I(N__36231));
    Span4Mux_v I__3359 (
            .O(N__36231),
            .I(N__36228));
    Span4Mux_v I__3358 (
            .O(N__36228),
            .I(N__36225));
    Odrv4 I__3357 (
            .O(N__36225),
            .I(\c0.n32762 ));
    CascadeMux I__3356 (
            .O(N__36222),
            .I(N__36218));
    CascadeMux I__3355 (
            .O(N__36221),
            .I(N__36215));
    InMux I__3354 (
            .O(N__36218),
            .I(N__36212));
    InMux I__3353 (
            .O(N__36215),
            .I(N__36208));
    LocalMux I__3352 (
            .O(N__36212),
            .I(N__36205));
    InMux I__3351 (
            .O(N__36211),
            .I(N__36202));
    LocalMux I__3350 (
            .O(N__36208),
            .I(N__36197));
    Span4Mux_h I__3349 (
            .O(N__36205),
            .I(N__36197));
    LocalMux I__3348 (
            .O(N__36202),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv4 I__3347 (
            .O(N__36197),
            .I(\c0.FRAME_MATCHER_state_6 ));
    CascadeMux I__3346 (
            .O(N__36192),
            .I(N__36188));
    InMux I__3345 (
            .O(N__36191),
            .I(N__36185));
    InMux I__3344 (
            .O(N__36188),
            .I(N__36181));
    LocalMux I__3343 (
            .O(N__36185),
            .I(N__36178));
    InMux I__3342 (
            .O(N__36184),
            .I(N__36175));
    LocalMux I__3341 (
            .O(N__36181),
            .I(N__36170));
    Span4Mux_h I__3340 (
            .O(N__36178),
            .I(N__36170));
    LocalMux I__3339 (
            .O(N__36175),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__3338 (
            .O(N__36170),
            .I(\c0.FRAME_MATCHER_state_4 ));
    CascadeMux I__3337 (
            .O(N__36165),
            .I(N__36162));
    InMux I__3336 (
            .O(N__36162),
            .I(N__36156));
    InMux I__3335 (
            .O(N__36161),
            .I(N__36156));
    LocalMux I__3334 (
            .O(N__36156),
            .I(N__36152));
    InMux I__3333 (
            .O(N__36155),
            .I(N__36149));
    Span12Mux_h I__3332 (
            .O(N__36152),
            .I(N__36146));
    LocalMux I__3331 (
            .O(N__36149),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv12 I__3330 (
            .O(N__36146),
            .I(\c0.FRAME_MATCHER_state_8 ));
    InMux I__3329 (
            .O(N__36141),
            .I(N__36138));
    LocalMux I__3328 (
            .O(N__36138),
            .I(N__36133));
    InMux I__3327 (
            .O(N__36137),
            .I(N__36130));
    InMux I__3326 (
            .O(N__36136),
            .I(N__36127));
    Span4Mux_h I__3325 (
            .O(N__36133),
            .I(N__36124));
    LocalMux I__3324 (
            .O(N__36130),
            .I(\c0.FRAME_MATCHER_state_13 ));
    LocalMux I__3323 (
            .O(N__36127),
            .I(\c0.FRAME_MATCHER_state_13 ));
    Odrv4 I__3322 (
            .O(N__36124),
            .I(\c0.FRAME_MATCHER_state_13 ));
    CascadeMux I__3321 (
            .O(N__36117),
            .I(\c0.n17_adj_4788_cascade_ ));
    CascadeMux I__3320 (
            .O(N__36114),
            .I(a_delay_counter_15__N_4220_cascade_));
    InMux I__3319 (
            .O(N__36111),
            .I(N__36107));
    InMux I__3318 (
            .O(N__36110),
            .I(N__36104));
    LocalMux I__3317 (
            .O(N__36107),
            .I(\c0.tx.r_Clock_Count_0 ));
    LocalMux I__3316 (
            .O(N__36104),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__3315 (
            .O(N__36099),
            .I(N__36095));
    InMux I__3314 (
            .O(N__36098),
            .I(N__36092));
    LocalMux I__3313 (
            .O(N__36095),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__3312 (
            .O(N__36092),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__3311 (
            .O(N__36087),
            .I(N__36083));
    InMux I__3310 (
            .O(N__36086),
            .I(N__36080));
    LocalMux I__3309 (
            .O(N__36083),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__3308 (
            .O(N__36080),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__3307 (
            .O(N__36075),
            .I(N__36071));
    InMux I__3306 (
            .O(N__36074),
            .I(N__36068));
    LocalMux I__3305 (
            .O(N__36071),
            .I(\c0.r_Clock_Count_2 ));
    LocalMux I__3304 (
            .O(N__36068),
            .I(\c0.r_Clock_Count_2 ));
    InMux I__3303 (
            .O(N__36063),
            .I(N__36059));
    InMux I__3302 (
            .O(N__36062),
            .I(N__36056));
    LocalMux I__3301 (
            .O(N__36059),
            .I(\c0.r_Clock_Count_4 ));
    LocalMux I__3300 (
            .O(N__36056),
            .I(\c0.r_Clock_Count_4 ));
    CascadeMux I__3299 (
            .O(N__36051),
            .I(\c0.n8_adj_4652_cascade_ ));
    CascadeMux I__3298 (
            .O(N__36048),
            .I(n22210_cascade_));
    SRMux I__3297 (
            .O(N__36045),
            .I(N__36042));
    LocalMux I__3296 (
            .O(N__36042),
            .I(N__36038));
    SRMux I__3295 (
            .O(N__36041),
            .I(N__36035));
    Sp12to4 I__3294 (
            .O(N__36038),
            .I(N__36032));
    LocalMux I__3293 (
            .O(N__36035),
            .I(N__36029));
    Odrv12 I__3292 (
            .O(N__36032),
            .I(\c0.tx.n19946 ));
    Odrv12 I__3291 (
            .O(N__36029),
            .I(\c0.tx.n19946 ));
    InMux I__3290 (
            .O(N__36024),
            .I(N__36016));
    InMux I__3289 (
            .O(N__36023),
            .I(N__36016));
    InMux I__3288 (
            .O(N__36022),
            .I(N__36011));
    InMux I__3287 (
            .O(N__36021),
            .I(N__36011));
    LocalMux I__3286 (
            .O(N__36016),
            .I(data_in_2_7));
    LocalMux I__3285 (
            .O(N__36011),
            .I(data_in_2_7));
    InMux I__3284 (
            .O(N__36006),
            .I(N__36002));
    InMux I__3283 (
            .O(N__36005),
            .I(N__35998));
    LocalMux I__3282 (
            .O(N__36002),
            .I(N__35995));
    InMux I__3281 (
            .O(N__36001),
            .I(N__35992));
    LocalMux I__3280 (
            .O(N__35998),
            .I(N__35989));
    Span4Mux_h I__3279 (
            .O(N__35995),
            .I(N__35986));
    LocalMux I__3278 (
            .O(N__35992),
            .I(data_in_0_7));
    Odrv4 I__3277 (
            .O(N__35989),
            .I(data_in_0_7));
    Odrv4 I__3276 (
            .O(N__35986),
            .I(data_in_0_7));
    InMux I__3275 (
            .O(N__35979),
            .I(N__35974));
    InMux I__3274 (
            .O(N__35978),
            .I(N__35971));
    InMux I__3273 (
            .O(N__35977),
            .I(N__35968));
    LocalMux I__3272 (
            .O(N__35974),
            .I(N__35963));
    LocalMux I__3271 (
            .O(N__35971),
            .I(N__35963));
    LocalMux I__3270 (
            .O(N__35968),
            .I(data_in_0_2));
    Odrv4 I__3269 (
            .O(N__35963),
            .I(data_in_0_2));
    InMux I__3268 (
            .O(N__35958),
            .I(N__35953));
    InMux I__3267 (
            .O(N__35957),
            .I(N__35948));
    InMux I__3266 (
            .O(N__35956),
            .I(N__35948));
    LocalMux I__3265 (
            .O(N__35953),
            .I(data_in_0_6));
    LocalMux I__3264 (
            .O(N__35948),
            .I(data_in_0_6));
    InMux I__3263 (
            .O(N__35943),
            .I(N__35934));
    InMux I__3262 (
            .O(N__35942),
            .I(N__35934));
    InMux I__3261 (
            .O(N__35941),
            .I(N__35934));
    LocalMux I__3260 (
            .O(N__35934),
            .I(data_in_1_7));
    InMux I__3259 (
            .O(N__35931),
            .I(N__35925));
    InMux I__3258 (
            .O(N__35930),
            .I(N__35925));
    LocalMux I__3257 (
            .O(N__35925),
            .I(\c0.n10_adj_4531 ));
    IoInMux I__3256 (
            .O(N__35922),
            .I(N__35919));
    LocalMux I__3255 (
            .O(N__35919),
            .I(N__35916));
    Span12Mux_s6_v I__3254 (
            .O(N__35916),
            .I(N__35913));
    Odrv12 I__3253 (
            .O(N__35913),
            .I(LED_c));
    InMux I__3252 (
            .O(N__35910),
            .I(N__35907));
    LocalMux I__3251 (
            .O(N__35907),
            .I(\c0.n6_adj_4532 ));
    InMux I__3250 (
            .O(N__35904),
            .I(N__35901));
    LocalMux I__3249 (
            .O(N__35901),
            .I(\c0.n15_adj_4796 ));
    CascadeMux I__3248 (
            .O(N__35898),
            .I(\c0.n18_adj_4794_cascade_ ));
    CascadeMux I__3247 (
            .O(N__35895),
            .I(N__35892));
    InMux I__3246 (
            .O(N__35892),
            .I(N__35889));
    LocalMux I__3245 (
            .O(N__35889),
            .I(N__35886));
    Odrv4 I__3244 (
            .O(N__35886),
            .I(\c0.n20_adj_4795 ));
    InMux I__3243 (
            .O(N__35883),
            .I(N__35880));
    LocalMux I__3242 (
            .O(N__35880),
            .I(\c0.n18086 ));
    InMux I__3241 (
            .O(N__35877),
            .I(N__35871));
    InMux I__3240 (
            .O(N__35876),
            .I(N__35871));
    LocalMux I__3239 (
            .O(N__35871),
            .I(\c0.n115 ));
    SRMux I__3238 (
            .O(N__35868),
            .I(N__35865));
    LocalMux I__3237 (
            .O(N__35865),
            .I(N__35862));
    Odrv12 I__3236 (
            .O(N__35862),
            .I(\c0.n32734 ));
    SRMux I__3235 (
            .O(N__35859),
            .I(N__35856));
    LocalMux I__3234 (
            .O(N__35856),
            .I(N__35853));
    Odrv4 I__3233 (
            .O(N__35853),
            .I(\c0.n32716 ));
    InMux I__3232 (
            .O(N__35850),
            .I(N__35847));
    LocalMux I__3231 (
            .O(N__35847),
            .I(\c0.n14_adj_4792 ));
    CascadeMux I__3230 (
            .O(N__35844),
            .I(\c0.n15_adj_4793_cascade_ ));
    CascadeMux I__3229 (
            .O(N__35841),
            .I(\c0.n63_cascade_ ));
    InMux I__3228 (
            .O(N__35838),
            .I(N__35832));
    InMux I__3227 (
            .O(N__35837),
            .I(N__35832));
    LocalMux I__3226 (
            .O(N__35832),
            .I(\c0.n118_adj_4786 ));
    InMux I__3225 (
            .O(N__35829),
            .I(\c0.tx.n30071 ));
    InMux I__3224 (
            .O(N__35826),
            .I(\c0.tx.n30072 ));
    InMux I__3223 (
            .O(N__35823),
            .I(\c0.tx.n30073 ));
    InMux I__3222 (
            .O(N__35820),
            .I(\c0.tx.n30074 ));
    InMux I__3221 (
            .O(N__35817),
            .I(bfn_5_12_0_));
    InMux I__3220 (
            .O(N__35814),
            .I(N__35810));
    CascadeMux I__3219 (
            .O(N__35813),
            .I(N__35806));
    LocalMux I__3218 (
            .O(N__35810),
            .I(N__35803));
    InMux I__3217 (
            .O(N__35809),
            .I(N__35798));
    InMux I__3216 (
            .O(N__35806),
            .I(N__35798));
    Span4Mux_v I__3215 (
            .O(N__35803),
            .I(N__35795));
    LocalMux I__3214 (
            .O(N__35798),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__3213 (
            .O(N__35795),
            .I(\c0.FRAME_MATCHER_state_24 ));
    SRMux I__3212 (
            .O(N__35790),
            .I(N__35787));
    LocalMux I__3211 (
            .O(N__35787),
            .I(N__35784));
    Span4Mux_h I__3210 (
            .O(N__35784),
            .I(N__35781));
    Odrv4 I__3209 (
            .O(N__35781),
            .I(\c0.n32810 ));
    SRMux I__3208 (
            .O(N__35778),
            .I(N__35775));
    LocalMux I__3207 (
            .O(N__35775),
            .I(\c0.n32722 ));
    CascadeMux I__3206 (
            .O(N__35772),
            .I(N__35768));
    CascadeMux I__3205 (
            .O(N__35771),
            .I(N__35765));
    InMux I__3204 (
            .O(N__35768),
            .I(N__35761));
    InMux I__3203 (
            .O(N__35765),
            .I(N__35756));
    InMux I__3202 (
            .O(N__35764),
            .I(N__35756));
    LocalMux I__3201 (
            .O(N__35761),
            .I(\c0.FRAME_MATCHER_state_28 ));
    LocalMux I__3200 (
            .O(N__35756),
            .I(\c0.FRAME_MATCHER_state_28 ));
    SRMux I__3199 (
            .O(N__35751),
            .I(N__35748));
    LocalMux I__3198 (
            .O(N__35748),
            .I(N__35745));
    Span4Mux_h I__3197 (
            .O(N__35745),
            .I(N__35742));
    Odrv4 I__3196 (
            .O(N__35742),
            .I(\c0.n32828 ));
    InMux I__3195 (
            .O(N__35739),
            .I(N__35735));
    InMux I__3194 (
            .O(N__35738),
            .I(N__35731));
    LocalMux I__3193 (
            .O(N__35735),
            .I(N__35728));
    InMux I__3192 (
            .O(N__35734),
            .I(N__35725));
    LocalMux I__3191 (
            .O(N__35731),
            .I(\c0.FRAME_MATCHER_state_26 ));
    Odrv4 I__3190 (
            .O(N__35728),
            .I(\c0.FRAME_MATCHER_state_26 ));
    LocalMux I__3189 (
            .O(N__35725),
            .I(\c0.FRAME_MATCHER_state_26 ));
    SRMux I__3188 (
            .O(N__35718),
            .I(N__35715));
    LocalMux I__3187 (
            .O(N__35715),
            .I(N__35712));
    Odrv12 I__3186 (
            .O(N__35712),
            .I(\c0.n32822 ));
    InMux I__3185 (
            .O(N__35709),
            .I(bfn_5_11_0_));
    InMux I__3184 (
            .O(N__35706),
            .I(\c0.tx.n30068 ));
    InMux I__3183 (
            .O(N__35703),
            .I(\c0.tx.n30069 ));
    InMux I__3182 (
            .O(N__35700),
            .I(\c0.tx.n30070 ));
    SRMux I__3181 (
            .O(N__35697),
            .I(N__35694));
    LocalMux I__3180 (
            .O(N__35694),
            .I(N__35691));
    Span4Mux_h I__3179 (
            .O(N__35691),
            .I(N__35688));
    Odrv4 I__3178 (
            .O(N__35688),
            .I(\c0.n32834 ));
    CascadeMux I__3177 (
            .O(N__35685),
            .I(\c0.n3_adj_4636_cascade_ ));
    SRMux I__3176 (
            .O(N__35682),
            .I(N__35679));
    LocalMux I__3175 (
            .O(N__35679),
            .I(\c0.n32710 ));
    SRMux I__3174 (
            .O(N__35676),
            .I(N__35673));
    LocalMux I__3173 (
            .O(N__35673),
            .I(N__35670));
    Span4Mux_s3_h I__3172 (
            .O(N__35670),
            .I(N__35667));
    Odrv4 I__3171 (
            .O(N__35667),
            .I(\c0.n32816 ));
    CascadeMux I__3170 (
            .O(N__35664),
            .I(N__35660));
    InMux I__3169 (
            .O(N__35663),
            .I(N__35657));
    InMux I__3168 (
            .O(N__35660),
            .I(N__35654));
    LocalMux I__3167 (
            .O(N__35657),
            .I(N__35650));
    LocalMux I__3166 (
            .O(N__35654),
            .I(N__35647));
    InMux I__3165 (
            .O(N__35653),
            .I(N__35644));
    Span4Mux_h I__3164 (
            .O(N__35650),
            .I(N__35641));
    Span4Mux_h I__3163 (
            .O(N__35647),
            .I(N__35638));
    LocalMux I__3162 (
            .O(N__35644),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__3161 (
            .O(N__35641),
            .I(\c0.FRAME_MATCHER_state_25 ));
    Odrv4 I__3160 (
            .O(N__35638),
            .I(\c0.FRAME_MATCHER_state_25 ));
    CascadeMux I__3159 (
            .O(N__35631),
            .I(n3_cascade_));
    IoInMux I__3158 (
            .O(N__35628),
            .I(N__35625));
    LocalMux I__3157 (
            .O(N__35625),
            .I(N__35622));
    Span4Mux_s3_h I__3156 (
            .O(N__35622),
            .I(N__35618));
    InMux I__3155 (
            .O(N__35621),
            .I(N__35615));
    Span4Mux_v I__3154 (
            .O(N__35618),
            .I(N__35612));
    LocalMux I__3153 (
            .O(N__35615),
            .I(N__35609));
    Span4Mux_v I__3152 (
            .O(N__35612),
            .I(N__35605));
    Span12Mux_s3_h I__3151 (
            .O(N__35609),
            .I(N__35602));
    InMux I__3150 (
            .O(N__35608),
            .I(N__35599));
    Odrv4 I__3149 (
            .O(N__35605),
            .I(tx_o));
    Odrv12 I__3148 (
            .O(N__35602),
            .I(tx_o));
    LocalMux I__3147 (
            .O(N__35599),
            .I(tx_o));
    SRMux I__3146 (
            .O(N__35592),
            .I(N__35589));
    LocalMux I__3145 (
            .O(N__35589),
            .I(N__35586));
    Span4Mux_h I__3144 (
            .O(N__35586),
            .I(N__35583));
    Odrv4 I__3143 (
            .O(N__35583),
            .I(\c0.n32792 ));
    CascadeMux I__3142 (
            .O(N__35580),
            .I(N__35575));
    CascadeMux I__3141 (
            .O(N__35579),
            .I(N__35572));
    InMux I__3140 (
            .O(N__35578),
            .I(N__35565));
    InMux I__3139 (
            .O(N__35575),
            .I(N__35565));
    InMux I__3138 (
            .O(N__35572),
            .I(N__35565));
    LocalMux I__3137 (
            .O(N__35565),
            .I(\c0.FRAME_MATCHER_state_17 ));
    InMux I__3136 (
            .O(N__35562),
            .I(N__35556));
    InMux I__3135 (
            .O(N__35561),
            .I(N__35556));
    LocalMux I__3134 (
            .O(N__35556),
            .I(N__35552));
    InMux I__3133 (
            .O(N__35555),
            .I(N__35549));
    Span4Mux_h I__3132 (
            .O(N__35552),
            .I(N__35546));
    LocalMux I__3131 (
            .O(N__35549),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv4 I__3130 (
            .O(N__35546),
            .I(\c0.FRAME_MATCHER_state_16 ));
    SRMux I__3129 (
            .O(N__35541),
            .I(N__35538));
    LocalMux I__3128 (
            .O(N__35538),
            .I(N__35535));
    Span4Mux_s3_h I__3127 (
            .O(N__35535),
            .I(N__35532));
    Odrv4 I__3126 (
            .O(N__35532),
            .I(\c0.n32786 ));
    SRMux I__3125 (
            .O(N__35529),
            .I(N__35526));
    LocalMux I__3124 (
            .O(N__35526),
            .I(\c0.n32780 ));
    SRMux I__3123 (
            .O(N__35523),
            .I(N__35520));
    LocalMux I__3122 (
            .O(N__35520),
            .I(N__35517));
    Odrv12 I__3121 (
            .O(N__35517),
            .I(\c0.n32774 ));
    InMux I__3120 (
            .O(N__35514),
            .I(N__35510));
    InMux I__3119 (
            .O(N__35513),
            .I(N__35507));
    LocalMux I__3118 (
            .O(N__35510),
            .I(\quad_counter0.b_delay_counter_11 ));
    LocalMux I__3117 (
            .O(N__35507),
            .I(\quad_counter0.b_delay_counter_11 ));
    InMux I__3116 (
            .O(N__35502),
            .I(\quad_counter0.n30011 ));
    CascadeMux I__3115 (
            .O(N__35499),
            .I(N__35495));
    InMux I__3114 (
            .O(N__35498),
            .I(N__35492));
    InMux I__3113 (
            .O(N__35495),
            .I(N__35489));
    LocalMux I__3112 (
            .O(N__35492),
            .I(\quad_counter0.b_delay_counter_12 ));
    LocalMux I__3111 (
            .O(N__35489),
            .I(\quad_counter0.b_delay_counter_12 ));
    InMux I__3110 (
            .O(N__35484),
            .I(\quad_counter0.n30012 ));
    CascadeMux I__3109 (
            .O(N__35481),
            .I(N__35477));
    InMux I__3108 (
            .O(N__35480),
            .I(N__35474));
    InMux I__3107 (
            .O(N__35477),
            .I(N__35471));
    LocalMux I__3106 (
            .O(N__35474),
            .I(\quad_counter0.b_delay_counter_13 ));
    LocalMux I__3105 (
            .O(N__35471),
            .I(\quad_counter0.b_delay_counter_13 ));
    InMux I__3104 (
            .O(N__35466),
            .I(\quad_counter0.n30013 ));
    InMux I__3103 (
            .O(N__35463),
            .I(N__35459));
    InMux I__3102 (
            .O(N__35462),
            .I(N__35456));
    LocalMux I__3101 (
            .O(N__35459),
            .I(\quad_counter0.b_delay_counter_14 ));
    LocalMux I__3100 (
            .O(N__35456),
            .I(\quad_counter0.b_delay_counter_14 ));
    InMux I__3099 (
            .O(N__35451),
            .I(\quad_counter0.n30014 ));
    InMux I__3098 (
            .O(N__35448),
            .I(\quad_counter0.n30015 ));
    InMux I__3097 (
            .O(N__35445),
            .I(N__35441));
    InMux I__3096 (
            .O(N__35444),
            .I(N__35438));
    LocalMux I__3095 (
            .O(N__35441),
            .I(\quad_counter0.b_delay_counter_15 ));
    LocalMux I__3094 (
            .O(N__35438),
            .I(\quad_counter0.b_delay_counter_15 ));
    CascadeMux I__3093 (
            .O(N__35433),
            .I(N__35430));
    InMux I__3092 (
            .O(N__35430),
            .I(N__35427));
    LocalMux I__3091 (
            .O(N__35427),
            .I(N__35422));
    InMux I__3090 (
            .O(N__35426),
            .I(N__35417));
    InMux I__3089 (
            .O(N__35425),
            .I(N__35417));
    Odrv4 I__3088 (
            .O(N__35422),
            .I(quadB_delayed));
    LocalMux I__3087 (
            .O(N__35417),
            .I(quadB_delayed));
    InMux I__3086 (
            .O(N__35412),
            .I(N__35405));
    InMux I__3085 (
            .O(N__35411),
            .I(N__35405));
    InMux I__3084 (
            .O(N__35410),
            .I(N__35401));
    LocalMux I__3083 (
            .O(N__35405),
            .I(N__35398));
    InMux I__3082 (
            .O(N__35404),
            .I(N__35395));
    LocalMux I__3081 (
            .O(N__35401),
            .I(N__35392));
    Span4Mux_v I__3080 (
            .O(N__35398),
            .I(N__35387));
    LocalMux I__3079 (
            .O(N__35395),
            .I(N__35387));
    Span4Mux_v I__3078 (
            .O(N__35392),
            .I(N__35384));
    Span4Mux_h I__3077 (
            .O(N__35387),
            .I(N__35381));
    Span4Mux_v I__3076 (
            .O(N__35384),
            .I(N__35378));
    Span4Mux_v I__3075 (
            .O(N__35381),
            .I(N__35375));
    Odrv4 I__3074 (
            .O(N__35378),
            .I(PIN_8_c));
    Odrv4 I__3073 (
            .O(N__35375),
            .I(PIN_8_c));
    CascadeMux I__3072 (
            .O(N__35370),
            .I(b_delay_counter_15__N_4237_cascade_));
    InMux I__3071 (
            .O(N__35367),
            .I(N__35364));
    LocalMux I__3070 (
            .O(N__35364),
            .I(N__35360));
    InMux I__3069 (
            .O(N__35363),
            .I(N__35357));
    Odrv4 I__3068 (
            .O(N__35360),
            .I(n17987));
    LocalMux I__3067 (
            .O(N__35357),
            .I(n17987));
    CEMux I__3066 (
            .O(N__35352),
            .I(N__35348));
    CEMux I__3065 (
            .O(N__35351),
            .I(N__35345));
    LocalMux I__3064 (
            .O(N__35348),
            .I(N__35342));
    LocalMux I__3063 (
            .O(N__35345),
            .I(N__35339));
    Span4Mux_v I__3062 (
            .O(N__35342),
            .I(N__35336));
    Odrv4 I__3061 (
            .O(N__35339),
            .I(n19282));
    Odrv4 I__3060 (
            .O(N__35336),
            .I(n19282));
    InMux I__3059 (
            .O(N__35331),
            .I(N__35328));
    LocalMux I__3058 (
            .O(N__35328),
            .I(N__35325));
    Odrv4 I__3057 (
            .O(N__35325),
            .I(n187));
    SRMux I__3056 (
            .O(N__35322),
            .I(N__35319));
    LocalMux I__3055 (
            .O(N__35319),
            .I(N__35315));
    SRMux I__3054 (
            .O(N__35318),
            .I(N__35312));
    Span4Mux_v I__3053 (
            .O(N__35315),
            .I(N__35306));
    LocalMux I__3052 (
            .O(N__35312),
            .I(N__35306));
    InMux I__3051 (
            .O(N__35311),
            .I(N__35303));
    Odrv4 I__3050 (
            .O(N__35306),
            .I(b_delay_counter_15__N_4237));
    LocalMux I__3049 (
            .O(N__35303),
            .I(b_delay_counter_15__N_4237));
    CascadeMux I__3048 (
            .O(N__35298),
            .I(n19282_cascade_));
    InMux I__3047 (
            .O(N__35295),
            .I(N__35290));
    CascadeMux I__3046 (
            .O(N__35294),
            .I(N__35287));
    InMux I__3045 (
            .O(N__35293),
            .I(N__35284));
    LocalMux I__3044 (
            .O(N__35290),
            .I(N__35281));
    InMux I__3043 (
            .O(N__35287),
            .I(N__35278));
    LocalMux I__3042 (
            .O(N__35284),
            .I(b_delay_counter_0));
    Odrv4 I__3041 (
            .O(N__35281),
            .I(b_delay_counter_0));
    LocalMux I__3040 (
            .O(N__35278),
            .I(b_delay_counter_0));
    InMux I__3039 (
            .O(N__35271),
            .I(\quad_counter0.n30002 ));
    InMux I__3038 (
            .O(N__35268),
            .I(N__35264));
    InMux I__3037 (
            .O(N__35267),
            .I(N__35261));
    LocalMux I__3036 (
            .O(N__35264),
            .I(\quad_counter0.b_delay_counter_3 ));
    LocalMux I__3035 (
            .O(N__35261),
            .I(\quad_counter0.b_delay_counter_3 ));
    InMux I__3034 (
            .O(N__35256),
            .I(\quad_counter0.n30003 ));
    InMux I__3033 (
            .O(N__35253),
            .I(N__35249));
    InMux I__3032 (
            .O(N__35252),
            .I(N__35246));
    LocalMux I__3031 (
            .O(N__35249),
            .I(\quad_counter0.b_delay_counter_4 ));
    LocalMux I__3030 (
            .O(N__35246),
            .I(\quad_counter0.b_delay_counter_4 ));
    InMux I__3029 (
            .O(N__35241),
            .I(\quad_counter0.n30004 ));
    InMux I__3028 (
            .O(N__35238),
            .I(N__35234));
    InMux I__3027 (
            .O(N__35237),
            .I(N__35231));
    LocalMux I__3026 (
            .O(N__35234),
            .I(\quad_counter0.b_delay_counter_5 ));
    LocalMux I__3025 (
            .O(N__35231),
            .I(\quad_counter0.b_delay_counter_5 ));
    InMux I__3024 (
            .O(N__35226),
            .I(\quad_counter0.n30005 ));
    CascadeMux I__3023 (
            .O(N__35223),
            .I(N__35219));
    InMux I__3022 (
            .O(N__35222),
            .I(N__35216));
    InMux I__3021 (
            .O(N__35219),
            .I(N__35213));
    LocalMux I__3020 (
            .O(N__35216),
            .I(\quad_counter0.b_delay_counter_6 ));
    LocalMux I__3019 (
            .O(N__35213),
            .I(\quad_counter0.b_delay_counter_6 ));
    InMux I__3018 (
            .O(N__35208),
            .I(\quad_counter0.n30006 ));
    InMux I__3017 (
            .O(N__35205),
            .I(N__35201));
    InMux I__3016 (
            .O(N__35204),
            .I(N__35198));
    LocalMux I__3015 (
            .O(N__35201),
            .I(\quad_counter0.b_delay_counter_7 ));
    LocalMux I__3014 (
            .O(N__35198),
            .I(\quad_counter0.b_delay_counter_7 ));
    InMux I__3013 (
            .O(N__35193),
            .I(\quad_counter0.n30007 ));
    InMux I__3012 (
            .O(N__35190),
            .I(N__35186));
    InMux I__3011 (
            .O(N__35189),
            .I(N__35183));
    LocalMux I__3010 (
            .O(N__35186),
            .I(\quad_counter0.b_delay_counter_8 ));
    LocalMux I__3009 (
            .O(N__35183),
            .I(\quad_counter0.b_delay_counter_8 ));
    InMux I__3008 (
            .O(N__35178),
            .I(bfn_4_11_0_));
    InMux I__3007 (
            .O(N__35175),
            .I(N__35171));
    InMux I__3006 (
            .O(N__35174),
            .I(N__35168));
    LocalMux I__3005 (
            .O(N__35171),
            .I(\quad_counter0.b_delay_counter_9 ));
    LocalMux I__3004 (
            .O(N__35168),
            .I(\quad_counter0.b_delay_counter_9 ));
    InMux I__3003 (
            .O(N__35163),
            .I(\quad_counter0.n30009 ));
    InMux I__3002 (
            .O(N__35160),
            .I(N__35156));
    InMux I__3001 (
            .O(N__35159),
            .I(N__35153));
    LocalMux I__3000 (
            .O(N__35156),
            .I(\quad_counter0.b_delay_counter_10 ));
    LocalMux I__2999 (
            .O(N__35153),
            .I(\quad_counter0.b_delay_counter_10 ));
    InMux I__2998 (
            .O(N__35148),
            .I(\quad_counter0.n30010 ));
    SRMux I__2997 (
            .O(N__35145),
            .I(N__35142));
    LocalMux I__2996 (
            .O(N__35142),
            .I(N__35139));
    Odrv12 I__2995 (
            .O(N__35139),
            .I(\c0.n8_adj_4498 ));
    SRMux I__2994 (
            .O(N__35136),
            .I(N__35133));
    LocalMux I__2993 (
            .O(N__35133),
            .I(N__35130));
    Span4Mux_v I__2992 (
            .O(N__35130),
            .I(N__35127));
    Odrv4 I__2991 (
            .O(N__35127),
            .I(\c0.n8_adj_4494 ));
    InMux I__2990 (
            .O(N__35124),
            .I(bfn_4_10_0_));
    InMux I__2989 (
            .O(N__35121),
            .I(N__35117));
    InMux I__2988 (
            .O(N__35120),
            .I(N__35114));
    LocalMux I__2987 (
            .O(N__35117),
            .I(\quad_counter0.b_delay_counter_1 ));
    LocalMux I__2986 (
            .O(N__35114),
            .I(\quad_counter0.b_delay_counter_1 ));
    InMux I__2985 (
            .O(N__35109),
            .I(\quad_counter0.n30001 ));
    InMux I__2984 (
            .O(N__35106),
            .I(N__35102));
    InMux I__2983 (
            .O(N__35105),
            .I(N__35099));
    LocalMux I__2982 (
            .O(N__35102),
            .I(\quad_counter0.b_delay_counter_2 ));
    LocalMux I__2981 (
            .O(N__35099),
            .I(\quad_counter0.b_delay_counter_2 ));
    InMux I__2980 (
            .O(N__35094),
            .I(N__35091));
    LocalMux I__2979 (
            .O(N__35091),
            .I(\quad_counter0.n28_adj_4414 ));
    InMux I__2978 (
            .O(N__35088),
            .I(N__35085));
    LocalMux I__2977 (
            .O(N__35085),
            .I(\quad_counter0.n26_adj_4415 ));
    CascadeMux I__2976 (
            .O(N__35082),
            .I(\quad_counter0.n25_adj_4417_cascade_ ));
    InMux I__2975 (
            .O(N__35079),
            .I(N__35076));
    LocalMux I__2974 (
            .O(N__35076),
            .I(\quad_counter0.n27_adj_4416 ));
    SRMux I__2973 (
            .O(N__35073),
            .I(N__35070));
    LocalMux I__2972 (
            .O(N__35070),
            .I(N__35067));
    Odrv4 I__2971 (
            .O(N__35067),
            .I(\c0.n32768 ));
    SRMux I__2970 (
            .O(N__35064),
            .I(N__35061));
    LocalMux I__2969 (
            .O(N__35061),
            .I(N__35058));
    Span4Mux_s3_h I__2968 (
            .O(N__35058),
            .I(N__35055));
    Odrv4 I__2967 (
            .O(N__35055),
            .I(\c0.n32756 ));
    IoInMux I__2966 (
            .O(N__35052),
            .I(N__35049));
    LocalMux I__2965 (
            .O(N__35049),
            .I(N__35046));
    Span4Mux_s1_v I__2964 (
            .O(N__35046),
            .I(N__35043));
    Span4Mux_v I__2963 (
            .O(N__35043),
            .I(N__35040));
    Sp12to4 I__2962 (
            .O(N__35040),
            .I(N__35037));
    Span12Mux_h I__2961 (
            .O(N__35037),
            .I(N__35034));
    Span12Mux_v I__2960 (
            .O(N__35034),
            .I(N__35031));
    Span12Mux_v I__2959 (
            .O(N__35031),
            .I(N__35028));
    Odrv12 I__2958 (
            .O(N__35028),
            .I(CLK_c));
    IoInMux I__2957 (
            .O(N__35025),
            .I(N__35022));
    LocalMux I__2956 (
            .O(N__35022),
            .I(N__35019));
    IoSpan4Mux I__2955 (
            .O(N__35019),
            .I(N__35016));
    Odrv4 I__2954 (
            .O(N__35016),
            .I(tx_enable));
    IoInMux I__2953 (
            .O(N__35013),
            .I(N__35010));
    LocalMux I__2952 (
            .O(N__35010),
            .I(GB_BUFFER_PIN_9_c_THRU_CO));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\quad_counter1.n30083 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\quad_counter1.n30091 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\quad_counter1.n30099 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\quad_counter1.n30107 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(\quad_counter0.n30115 ),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(\quad_counter0.n30123 ),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(\quad_counter0.n30131 ),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(\quad_counter0.n30139 ),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_23_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_12_0_));
    defparam IN_MUX_bfv_23_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_13_0_ (
            .carryinitin(\quad_counter1.n30682 ),
            .carryinitout(bfn_23_13_0_));
    defparam IN_MUX_bfv_23_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_14_0_ (
            .carryinitin(\quad_counter1.n30690 ),
            .carryinitout(bfn_23_14_0_));
    defparam IN_MUX_bfv_22_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_13_0_));
    defparam IN_MUX_bfv_22_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_14_0_ (
            .carryinitin(\quad_counter1.n30661 ),
            .carryinitout(bfn_22_14_0_));
    defparam IN_MUX_bfv_22_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_15_0_ (
            .carryinitin(\quad_counter1.n30669 ),
            .carryinitout(bfn_22_15_0_));
    defparam IN_MUX_bfv_19_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_11_0_));
    defparam IN_MUX_bfv_19_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_12_0_ (
            .carryinitin(\quad_counter1.n30641 ),
            .carryinitout(bfn_19_12_0_));
    defparam IN_MUX_bfv_19_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_13_0_ (
            .carryinitin(\quad_counter1.n30649 ),
            .carryinitout(bfn_19_13_0_));
    defparam IN_MUX_bfv_20_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_8_0_));
    defparam IN_MUX_bfv_20_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_9_0_ (
            .carryinitin(\quad_counter1.n30622 ),
            .carryinitout(bfn_20_9_0_));
    defparam IN_MUX_bfv_20_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_10_0_ (
            .carryinitin(\quad_counter1.n30630 ),
            .carryinitout(bfn_20_10_0_));
    defparam IN_MUX_bfv_19_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_5_0_));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(\quad_counter1.n30604 ),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(\quad_counter1.n30612 ),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_18_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_3_0_));
    defparam IN_MUX_bfv_18_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_4_0_ (
            .carryinitin(\quad_counter1.n30587 ),
            .carryinitout(bfn_18_4_0_));
    defparam IN_MUX_bfv_18_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_5_0_ (
            .carryinitin(\quad_counter1.n30595 ),
            .carryinitout(bfn_18_5_0_));
    defparam IN_MUX_bfv_19_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_2_0_));
    defparam IN_MUX_bfv_19_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_3_0_ (
            .carryinitin(\quad_counter1.n30571 ),
            .carryinitout(bfn_19_3_0_));
    defparam IN_MUX_bfv_19_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_4_0_ (
            .carryinitin(\quad_counter1.n30579 ),
            .carryinitout(bfn_19_4_0_));
    defparam IN_MUX_bfv_20_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_4_0_));
    defparam IN_MUX_bfv_20_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_5_0_ (
            .carryinitin(\quad_counter1.n30556 ),
            .carryinitout(bfn_20_5_0_));
    defparam IN_MUX_bfv_21_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_5_0_));
    defparam IN_MUX_bfv_21_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_6_0_ (
            .carryinitin(\quad_counter1.n30542 ),
            .carryinitout(bfn_21_6_0_));
    defparam IN_MUX_bfv_23_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_7_0_));
    defparam IN_MUX_bfv_23_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_8_0_ (
            .carryinitin(\quad_counter1.n30529 ),
            .carryinitout(bfn_23_8_0_));
    defparam IN_MUX_bfv_21_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_9_0_));
    defparam IN_MUX_bfv_21_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_10_0_ (
            .carryinitin(\quad_counter1.n30517 ),
            .carryinitout(bfn_21_10_0_));
    defparam IN_MUX_bfv_23_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_9_0_));
    defparam IN_MUX_bfv_23_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_10_0_ (
            .carryinitin(\quad_counter1.n30506 ),
            .carryinitout(bfn_23_10_0_));
    defparam IN_MUX_bfv_26_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_11_0_));
    defparam IN_MUX_bfv_26_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_12_0_ (
            .carryinitin(\quad_counter1.n30496 ),
            .carryinitout(bfn_26_12_0_));
    defparam IN_MUX_bfv_27_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_27_11_0_));
    defparam IN_MUX_bfv_27_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_12_0_ (
            .carryinitin(\quad_counter1.n30487 ),
            .carryinitout(bfn_27_12_0_));
    defparam IN_MUX_bfv_28_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_28_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_28_9_0_));
    defparam IN_MUX_bfv_28_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_28_10_0_ (
            .carryinitin(\quad_counter1.n30479 ),
            .carryinitout(bfn_28_10_0_));
    defparam IN_MUX_bfv_26_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_9_0_));
    defparam IN_MUX_bfv_26_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_8_0_));
    defparam IN_MUX_bfv_22_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_7_0_));
    defparam IN_MUX_bfv_22_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_8_0_ (
            .carryinitin(\quad_counter1.n30178 ),
            .carryinitout(bfn_22_8_0_));
    defparam IN_MUX_bfv_22_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_9_0_ (
            .carryinitin(\quad_counter1.n30186 ),
            .carryinitout(bfn_22_9_0_));
    defparam IN_MUX_bfv_22_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_10_0_ (
            .carryinitin(\quad_counter1.n30194 ),
            .carryinitout(bfn_22_10_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\quad_counter1.n30038 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\quad_counter1.n30053 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_22_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_11_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\quad_counter0.n30432 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\quad_counter0.n30440 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\quad_counter0.n30411 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\quad_counter0.n30419 ),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\quad_counter0.n30391 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(\quad_counter0.n30399 ),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(\quad_counter0.n30372 ),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\quad_counter0.n30380 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\quad_counter0.n30354 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\quad_counter0.n30362 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\quad_counter0.n30337 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\quad_counter0.n30345 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\quad_counter0.n30321 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\quad_counter0.n30329 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\quad_counter0.n30306 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\quad_counter0.n30292 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\quad_counter0.n30279 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\quad_counter0.n30267 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\quad_counter0.n30256 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\quad_counter0.n30246 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(\quad_counter0.n30237 ),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\quad_counter0.n30229 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\quad_counter0.n30147 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\quad_counter0.n30155 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\quad_counter0.n30163 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(\quad_counter0.n30008 ),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(\quad_counter0.n30023 ),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\c0.tx.n30075 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_24_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_1_0_));
    defparam IN_MUX_bfv_24_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_2_0_ (
            .carryinitin(\c0.n29970_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_2_0_));
    defparam IN_MUX_bfv_24_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_3_0_ (
            .carryinitin(\c0.n29971_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_3_0_));
    defparam IN_MUX_bfv_24_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_4_0_ (
            .carryinitin(\c0.n29972_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_4_0_));
    defparam IN_MUX_bfv_24_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_5_0_ (
            .carryinitin(\c0.n29973_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_5_0_));
    defparam IN_MUX_bfv_24_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_6_0_ (
            .carryinitin(\c0.n29974_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_6_0_));
    defparam IN_MUX_bfv_24_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_7_0_ (
            .carryinitin(\c0.n29975_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_7_0_));
    defparam IN_MUX_bfv_24_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_8_0_ (
            .carryinitin(\c0.n29976_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_8_0_));
    defparam IN_MUX_bfv_24_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_9_0_ (
            .carryinitin(\c0.n29977_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_9_0_));
    defparam IN_MUX_bfv_24_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_10_0_ (
            .carryinitin(\c0.n29978_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_10_0_));
    defparam IN_MUX_bfv_24_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_11_0_ (
            .carryinitin(\c0.n29979_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_11_0_));
    defparam IN_MUX_bfv_24_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_12_0_ (
            .carryinitin(\c0.n29980_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_12_0_));
    defparam IN_MUX_bfv_24_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_13_0_ (
            .carryinitin(\c0.n29981_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_13_0_));
    defparam IN_MUX_bfv_24_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_14_0_ (
            .carryinitin(\c0.n29982_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_14_0_));
    defparam IN_MUX_bfv_24_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_15_0_ (
            .carryinitin(\c0.n29983_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_15_0_));
    defparam IN_MUX_bfv_24_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_16_0_ (
            .carryinitin(\c0.n29984_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_16_0_));
    defparam IN_MUX_bfv_24_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_17_0_ (
            .carryinitin(\c0.n29985_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_17_0_));
    defparam IN_MUX_bfv_24_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_18_0_ (
            .carryinitin(\c0.n29986_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_18_0_));
    defparam IN_MUX_bfv_24_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_19_0_ (
            .carryinitin(\c0.n29987_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_19_0_));
    defparam IN_MUX_bfv_24_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_20_0_ (
            .carryinitin(\c0.n29988_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_20_0_));
    defparam IN_MUX_bfv_24_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_21_0_ (
            .carryinitin(\c0.n29989_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_21_0_));
    defparam IN_MUX_bfv_24_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_22_0_ (
            .carryinitin(\c0.n29990_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_22_0_));
    defparam IN_MUX_bfv_24_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_23_0_ (
            .carryinitin(\c0.n29991_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_23_0_));
    defparam IN_MUX_bfv_24_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_24_0_ (
            .carryinitin(\c0.n29992_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_24_0_));
    defparam IN_MUX_bfv_24_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_25_0_ (
            .carryinitin(\c0.n29993_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_25_0_));
    defparam IN_MUX_bfv_24_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_26_0_ (
            .carryinitin(\c0.n29994_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_26_0_));
    defparam IN_MUX_bfv_24_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_27_0_ (
            .carryinitin(\c0.n29995_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_27_0_));
    defparam IN_MUX_bfv_24_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_28_0_ (
            .carryinitin(\c0.n29996_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_28_0_));
    defparam IN_MUX_bfv_24_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_29_0_ (
            .carryinitin(\c0.n29997_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_29_0_));
    defparam IN_MUX_bfv_24_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_30_0_ (
            .carryinitin(\c0.n29998_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_30_0_));
    defparam IN_MUX_bfv_24_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_31_0_ (
            .carryinitin(\c0.n29999_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_31_0_));
    defparam IN_MUX_bfv_24_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_32_0_ (
            .carryinitin(\c0.n30000_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_24_32_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_5_1 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35621),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i16_LC_1_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_1_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_1_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__35555),
            .in2(_gnd_net_),
            .in3(N__71497),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97728),
            .ce(),
            .sr(N__35541));
    defparam \c0.FRAME_MATCHER_state_i14_LC_1_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_1_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_1_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__36493),
            .in2(_gnd_net_),
            .in3(N__71496),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97746),
            .ce(),
            .sr(N__35523));
    defparam GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_21_4.C_ON=1'b0;
    defparam GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_21_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_21_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_21_4 (
            .in0(N__97809),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_PIN_9_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i13_LC_2_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_2_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_2_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__36137),
            .in2(_gnd_net_),
            .in3(N__71495),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97717),
            .ce(),
            .sr(N__35073));
    defparam \c0.FRAME_MATCHER_state_i6_LC_2_14_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_2_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_2_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__36211),
            .in2(_gnd_net_),
            .in3(N__71494),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97733),
            .ce(),
            .sr(N__35145));
    defparam \c0.FRAME_MATCHER_state_i25_LC_2_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_2_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_2_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__35653),
            .in2(_gnd_net_),
            .in3(N__71473),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97752),
            .ce(),
            .sr(N__35676));
    defparam \quad_counter0.i12_4_lut_adj_1236_LC_3_10_2 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1236_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1236_LC_3_10_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1236_LC_3_10_2  (
            .in0(N__35105),
            .in1(N__35120),
            .in2(N__35481),
            .in3(N__35237),
            .lcout(\quad_counter0.n28_adj_4414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1237_LC_3_10_4 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1237_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1237_LC_3_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1237_LC_3_10_4  (
            .in0(N__35513),
            .in1(N__35159),
            .in2(N__35223),
            .in3(N__35189),
            .lcout(\quad_counter0.n26_adj_4415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_1239_LC_3_11_0 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_1239_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_1239_LC_3_11_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter0.i9_4_lut_adj_1239_LC_3_11_0  (
            .in0(N__35174),
            .in1(N__35267),
            .in2(N__35294),
            .in3(N__35252),
            .lcout(),
            .ltout(\quad_counter0.n25_adj_4417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_adj_1240_LC_3_11_1 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_adj_1240_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_adj_1240_LC_3_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_adj_1240_LC_3_11_1  (
            .in0(N__35094),
            .in1(N__35088),
            .in2(N__35082),
            .in3(N__35079),
            .lcout(n17987),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1238_LC_3_11_3 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1238_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1238_LC_3_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1238_LC_3_11_3  (
            .in0(N__35462),
            .in1(N__35204),
            .in2(N__35499),
            .in3(N__35444),
            .lcout(\quad_counter0.n27_adj_4416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadB_delayed_71_LC_3_11_5 .C_ON=1'b0;
    defparam \quad_counter0.quadB_delayed_71_LC_3_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadB_delayed_71_LC_3_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.quadB_delayed_71_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35410),
            .lcout(quadB_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i4_LC_3_12_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_3_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_3_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__36184),
            .in2(_gnd_net_),
            .in3(N__71493),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97682),
            .ce(),
            .sr(N__35064));
    defparam \quad_counter0.B_74_LC_3_13_7 .C_ON=1'b0;
    defparam \quad_counter0.B_74_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_74_LC_3_13_7 .LUT_INIT=16'b1010101011101000;
    LogicCell40 \quad_counter0.B_74_LC_3_13_7  (
            .in0(N__39416),
            .in1(N__35404),
            .in2(N__35433),
            .in3(N__35367),
            .lcout(B_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1609_LC_3_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1609_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1609_LC_3_14_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1609_LC_3_14_0  (
            .in0(N__46201),
            .in1(N__36136),
            .in2(N__45915),
            .in3(N__46029),
            .lcout(\c0.n32768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1620_LC_3_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1620_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1620_LC_3_14_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1620_LC_3_14_5  (
            .in0(N__46027),
            .in1(N__45910),
            .in2(N__36192),
            .in3(N__46199),
            .lcout(\c0.n32756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadA_delayed_70_LC_3_14_6 .C_ON=1'b0;
    defparam \quad_counter0.quadA_delayed_70_LC_3_14_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.quadA_delayed_70_LC_3_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.quadA_delayed_70_LC_3_14_6  (
            .in0(N__37214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadA_delayed),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97718),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1672_LC_3_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1672_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1672_LC_3_14_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1672_LC_3_14_7  (
            .in0(N__46028),
            .in1(N__45911),
            .in2(N__36221),
            .in3(N__46200),
            .lcout(\c0.n8_adj_4498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i22_LC_3_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_3_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_3_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__36398),
            .in2(_gnd_net_),
            .in3(N__71472),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97734),
            .ce(),
            .sr(N__36375));
    defparam \c0.FRAME_MATCHER_state_i27_LC_3_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_3_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_3_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__37385),
            .in2(_gnd_net_),
            .in3(N__71491),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97753),
            .ce(),
            .sr(N__35682));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1612_LC_3_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1612_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1612_LC_3_17_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1612_LC_3_17_1  (
            .in0(N__45894),
            .in1(N__45985),
            .in2(N__46300),
            .in3(N__46148),
            .lcout(\c0.n8_adj_4494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i12_LC_3_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_3_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_3_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__71490),
            .in2(_gnd_net_),
            .in3(N__46293),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97783),
            .ce(),
            .sr(N__35136));
    defparam \c0.FRAME_MATCHER_state_i8_LC_4_9_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_4_9_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_4_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__36155),
            .in2(_gnd_net_),
            .in3(N__71474),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97623),
            .ce(),
            .sr(N__36237));
    defparam \quad_counter0.add_98_2_lut_LC_4_10_0 .C_ON=1'b1;
    defparam \quad_counter0.add_98_2_lut_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_98_2_lut_LC_4_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_98_2_lut_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__35295),
            .in2(_gnd_net_),
            .in3(N__35124),
            .lcout(n187),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\quad_counter0.n30001 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i1_LC_4_10_1 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i1_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i1_LC_4_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i1_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__35121),
            .in2(_gnd_net_),
            .in3(N__35109),
            .lcout(\quad_counter0.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n30001 ),
            .carryout(\quad_counter0.n30002 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i2_LC_4_10_2 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i2_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i2_LC_4_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i2_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__35106),
            .in2(_gnd_net_),
            .in3(N__35271),
            .lcout(\quad_counter0.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n30002 ),
            .carryout(\quad_counter0.n30003 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i3_LC_4_10_3 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i3_LC_4_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i3_LC_4_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i3_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__35268),
            .in2(_gnd_net_),
            .in3(N__35256),
            .lcout(\quad_counter0.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n30003 ),
            .carryout(\quad_counter0.n30004 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i4_LC_4_10_4 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i4_LC_4_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i4_LC_4_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i4_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__35253),
            .in2(_gnd_net_),
            .in3(N__35241),
            .lcout(\quad_counter0.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n30004 ),
            .carryout(\quad_counter0.n30005 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i5_LC_4_10_5 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i5_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i5_LC_4_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i5_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(N__35238),
            .in2(_gnd_net_),
            .in3(N__35226),
            .lcout(\quad_counter0.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n30005 ),
            .carryout(\quad_counter0.n30006 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i6_LC_4_10_6 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i6_LC_4_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i6_LC_4_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i6_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(N__35222),
            .in2(_gnd_net_),
            .in3(N__35208),
            .lcout(\quad_counter0.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n30006 ),
            .carryout(\quad_counter0.n30007 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i7_LC_4_10_7 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i7_LC_4_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i7_LC_4_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i7_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(N__35205),
            .in2(_gnd_net_),
            .in3(N__35193),
            .lcout(\quad_counter0.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n30007 ),
            .carryout(\quad_counter0.n30008 ),
            .clk(N__97637),
            .ce(N__35351),
            .sr(N__35322));
    defparam \quad_counter0.b_delay_counter__i8_LC_4_11_0 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i8_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i8_LC_4_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i8_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__35190),
            .in2(_gnd_net_),
            .in3(N__35178),
            .lcout(\quad_counter0.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\quad_counter0.n30009 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i9_LC_4_11_1 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i9_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i9_LC_4_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i9_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__35175),
            .in2(_gnd_net_),
            .in3(N__35163),
            .lcout(\quad_counter0.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n30009 ),
            .carryout(\quad_counter0.n30010 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i10_LC_4_11_2 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i10_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i10_LC_4_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i10_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__35160),
            .in2(_gnd_net_),
            .in3(N__35148),
            .lcout(\quad_counter0.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n30010 ),
            .carryout(\quad_counter0.n30011 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i11_LC_4_11_3 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i11_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i11_LC_4_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i11_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__35514),
            .in2(_gnd_net_),
            .in3(N__35502),
            .lcout(\quad_counter0.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n30011 ),
            .carryout(\quad_counter0.n30012 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i12_LC_4_11_4 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i12_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i12_LC_4_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i12_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__35498),
            .in2(_gnd_net_),
            .in3(N__35484),
            .lcout(\quad_counter0.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n30012 ),
            .carryout(\quad_counter0.n30013 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i13_LC_4_11_5 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i13_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i13_LC_4_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i13_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__35480),
            .in2(_gnd_net_),
            .in3(N__35466),
            .lcout(\quad_counter0.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n30013 ),
            .carryout(\quad_counter0.n30014 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i14_LC_4_11_6 .C_ON=1'b1;
    defparam \quad_counter0.b_delay_counter__i14_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i14_LC_4_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i14_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(N__35463),
            .in2(_gnd_net_),
            .in3(N__35451),
            .lcout(\quad_counter0.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n30014 ),
            .carryout(\quad_counter0.n30015 ),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.b_delay_counter__i15_LC_4_11_7 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i15_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i15_LC_4_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.b_delay_counter__i15_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(N__35445),
            .in2(_gnd_net_),
            .in3(N__35448),
            .lcout(\quad_counter0.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97652),
            .ce(N__35352),
            .sr(N__35318));
    defparam \quad_counter0.quadB_I_0_91_2_lut_LC_4_12_0 .C_ON=1'b0;
    defparam \quad_counter0.quadB_I_0_91_2_lut_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadB_I_0_91_2_lut_LC_4_12_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter0.quadB_I_0_91_2_lut_LC_4_12_0  (
            .in0(N__35412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35425),
            .lcout(b_delay_counter_15__N_4237),
            .ltout(b_delay_counter_15__N_4237_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_4_12_1.C_ON=1'b0;
    defparam i1_4_lut_LC_4_12_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_4_12_1.LUT_INIT=16'b1111100111110000;
    LogicCell40 i1_4_lut_LC_4_12_1 (
            .in0(N__35426),
            .in1(N__35411),
            .in2(N__35370),
            .in3(N__35363),
            .lcout(n19282),
            .ltout(n19282_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_delay_counter__i0_LC_4_12_2 .C_ON=1'b0;
    defparam \quad_counter0.b_delay_counter__i0_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_delay_counter__i0_LC_4_12_2 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \quad_counter0.b_delay_counter__i0_LC_4_12_2  (
            .in0(N__35331),
            .in1(N__35311),
            .in2(N__35298),
            .in3(N__35293),
            .lcout(b_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_LC_4_12_4 .C_ON=1'b0;
    defparam \c0.i8_3_lut_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_LC_4_12_4 .LUT_INIT=16'b1011101110011001;
    LogicCell40 \c0.i8_3_lut_LC_4_12_4  (
            .in0(N__37602),
            .in1(N__37443),
            .in2(_gnd_net_),
            .in3(N__36261),
            .lcout(),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_4_12_5 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_4_12_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__35608),
            .in2(N__35631),
            .in3(N__37522),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i15_LC_4_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_4_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_4_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__36466),
            .in2(_gnd_net_),
            .in3(N__71488),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97683),
            .ce(),
            .sr(N__35529));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1605_LC_4_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1605_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1605_LC_4_14_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1605_LC_4_14_0  (
            .in0(N__45896),
            .in1(N__46196),
            .in2(N__35580),
            .in3(N__46019),
            .lcout(\c0.n32792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i17_LC_4_14_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_4_14_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_4_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__35578),
            .in2(_gnd_net_),
            .in3(N__71492),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97700),
            .ce(),
            .sr(N__35592));
    defparam \c0.i3_4_lut_adj_2018_LC_4_14_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_2018_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_2018_LC_4_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_2018_LC_4_14_2  (
            .in0(N__35561),
            .in1(N__36394),
            .in2(N__35579),
            .in3(N__36358),
            .lcout(\c0.n33166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1606_LC_4_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1606_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1606_LC_4_14_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1606_LC_4_14_3  (
            .in0(N__46195),
            .in1(N__35562),
            .in2(N__46053),
            .in3(N__45897),
            .lcout(\c0.n32786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1607_LC_4_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1607_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1607_LC_4_14_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1607_LC_4_14_4  (
            .in0(N__45899),
            .in1(N__46026),
            .in2(N__36470),
            .in3(N__46198),
            .lcout(\c0.n32780 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1608_LC_4_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1608_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1608_LC_4_14_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1608_LC_4_14_5  (
            .in0(N__46197),
            .in1(N__36495),
            .in2(N__46054),
            .in3(N__45898),
            .lcout(\c0.n32774 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i20_LC_4_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_4_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_4_15_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_4_15_0  (
            .in0(N__71445),
            .in1(N__36362),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97719),
            .ce(),
            .sr(N__36342));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1575_LC_4_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1575_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1575_LC_4_16_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1575_LC_4_16_0  (
            .in0(N__45904),
            .in1(N__45986),
            .in2(N__37875),
            .in3(N__46186),
            .lcout(\c0.n32834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i30_LC_4_16_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_4_16_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_4_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__37872),
            .in2(_gnd_net_),
            .in3(N__71505),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97735),
            .ce(),
            .sr(N__35697));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1579_LC_4_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1579_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1579_LC_4_16_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1579_LC_4_16_2  (
            .in0(N__45905),
            .in1(N__45987),
            .in2(N__35772),
            .in3(N__46187),
            .lcout(\c0.n32828 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1721_LC_4_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1721_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1721_LC_4_16_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1721_LC_4_16_3  (
            .in0(N__49050),
            .in1(N__48192),
            .in2(_gnd_net_),
            .in3(N__49262),
            .lcout(\c0.n3_adj_4636 ),
            .ltout(\c0.n3_adj_4636_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1583_LC_4_16_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1583_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1583_LC_4_16_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1583_LC_4_16_4  (
            .in0(N__45906),
            .in1(N__35739),
            .in2(N__35685),
            .in3(N__46188),
            .lcout(\c0.n32822 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1581_LC_4_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1581_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1581_LC_4_16_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1581_LC_4_16_5  (
            .in0(N__46190),
            .in1(N__37384),
            .in2(N__46032),
            .in3(N__45909),
            .lcout(\c0.n32710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1577_LC_4_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1577_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1577_LC_4_16_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1577_LC_4_16_6  (
            .in0(N__45908),
            .in1(N__45991),
            .in2(N__37830),
            .in3(N__46189),
            .lcout(\c0.n32716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1585_LC_4_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1585_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1585_LC_4_16_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1585_LC_4_16_7  (
            .in0(N__46185),
            .in1(N__35663),
            .in2(N__46031),
            .in3(N__45907),
            .lcout(\c0.n32816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_2022_LC_4_17_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_2022_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_2022_LC_4_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_2022_LC_4_17_0  (
            .in0(N__35734),
            .in1(N__35814),
            .in2(N__35664),
            .in3(N__35764),
            .lcout(\c0.n33163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i28_LC_4_17_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_4_17_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_4_17_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35771),
            .in3(N__71502),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97754),
            .ce(),
            .sr(N__35751));
    defparam \c0.i3_4_lut_adj_2029_LC_4_17_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_2029_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_2029_LC_4_17_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i3_4_lut_adj_2029_LC_4_17_4  (
            .in0(N__35978),
            .in1(N__36006),
            .in2(N__38303),
            .in3(N__38335),
            .lcout(\c0.n14_adj_4784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_2037_LC_4_17_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_2037_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_2037_LC_4_17_7 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \c0.i5_3_lut_adj_2037_LC_4_17_7  (
            .in0(N__38336),
            .in1(_gnd_net_),
            .in2(N__36777),
            .in3(N__38139),
            .lcout(\c0.n14_adj_4792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i26_LC_4_18_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_4_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_4_18_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_4_18_0  (
            .in0(N__71503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35738),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97768),
            .ce(),
            .sr(N__35718));
    defparam \c0.FRAME_MATCHER_state_i9_LC_5_10_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_5_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_5_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__36601),
            .in2(_gnd_net_),
            .in3(N__71475),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97624),
            .ce(),
            .sr(N__36585));
    defparam \c0.tx.r_Clock_Count__i0_LC_5_11_0 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i0_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__36111),
            .in2(_gnd_net_),
            .in3(N__35709),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\c0.tx.n30068 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i1_LC_5_11_1 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i1_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__36087),
            .in2(_gnd_net_),
            .in3(N__35706),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx.n30068 ),
            .carryout(\c0.tx.n30069 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i2_LC_5_11_2 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i2_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__36075),
            .in2(_gnd_net_),
            .in3(N__35703),
            .lcout(\c0.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx.n30069 ),
            .carryout(\c0.tx.n30070 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i3_LC_5_11_3 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i3_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__36099),
            .in2(_gnd_net_),
            .in3(N__35700),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx.n30070 ),
            .carryout(\c0.tx.n30071 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i4_LC_5_11_4 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i4_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__36063),
            .in2(_gnd_net_),
            .in3(N__35829),
            .lcout(\c0.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx.n30071 ),
            .carryout(\c0.tx.n30072 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i5_LC_5_11_5 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i5_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__36321),
            .in2(_gnd_net_),
            .in3(N__35826),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx.n30072 ),
            .carryout(\c0.tx.n30073 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i6_LC_5_11_6 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i6_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__36296),
            .in2(_gnd_net_),
            .in3(N__35823),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx.n30073 ),
            .carryout(\c0.tx.n30074 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i7_LC_5_11_7 .C_ON=1'b1;
    defparam \c0.tx.r_Clock_Count__i7_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__36309),
            .in2(_gnd_net_),
            .in3(N__35820),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx.n30074 ),
            .carryout(\c0.tx.n30075 ),
            .clk(N__97638),
            .ce(N__37527),
            .sr(N__36041));
    defparam \c0.tx.r_Clock_Count__i8_LC_5_12_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__36282),
            .in2(_gnd_net_),
            .in3(N__35817),
            .lcout(\c0.tx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97653),
            .ce(N__37526),
            .sr(N__36045));
    defparam \c0.FRAME_MATCHER_state_i11_LC_5_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_5_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_5_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__36444),
            .in2(_gnd_net_),
            .in3(N__71499),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97667),
            .ce(),
            .sr(N__35778));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_5_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_5_14_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_5_14_0  (
            .in0(N__45837),
            .in1(N__46030),
            .in2(N__35813),
            .in3(N__46194),
            .lcout(\c0.n32810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i24_LC_5_14_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_5_14_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_5_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__71489),
            .in2(_gnd_net_),
            .in3(N__35809),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97684),
            .ce(),
            .sr(N__35790));
    defparam \c0.i1_2_lut_adj_1545_LC_5_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1545_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1545_LC_5_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1545_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__36443),
            .in2(_gnd_net_),
            .in3(N__42659),
            .lcout(\c0.n32722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i116_2_lut_LC_5_14_6 .C_ON=1'b0;
    defparam \c0.i116_2_lut_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i116_2_lut_LC_5_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i116_2_lut_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__45809),
            .in2(_gnd_net_),
            .in3(N__46193),
            .lcout(\c0.n93_adj_4634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1567_LC_5_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1567_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1567_LC_5_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1567_LC_5_14_7  (
            .in0(N__42660),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37927),
            .lcout(\c0.n32734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i21_LC_5_15_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_5_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_5_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__37921),
            .in2(_gnd_net_),
            .in3(N__71444),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97701),
            .ce(),
            .sr(N__35868));
    defparam \c0.FRAME_MATCHER_state_i29_LC_5_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_5_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_5_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__37821),
            .in2(_gnd_net_),
            .in3(N__71504),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97720),
            .ce(),
            .sr(N__35859));
    defparam \c0.i1_2_lut_adj_2040_LC_5_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2040_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2040_LC_5_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_2040_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__35876),
            .in2(_gnd_net_),
            .in3(N__35837),
            .lcout(\c0.n107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2038_LC_5_17_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2038_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2038_LC_5_17_1 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i6_4_lut_adj_2038_LC_5_17_1  (
            .in0(N__35979),
            .in1(N__36005),
            .in2(N__38304),
            .in3(N__36653),
            .lcout(),
            .ltout(\c0.n15_adj_4793_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_2039_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_2039_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_2039_LC_5_17_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i8_4_lut_adj_2039_LC_5_17_2  (
            .in0(N__35850),
            .in1(N__48707),
            .in2(N__35844),
            .in3(N__42945),
            .lcout(\c0.n33266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_2027_LC_5_17_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_2027_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_2027_LC_5_17_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i4_4_lut_adj_2027_LC_5_17_4  (
            .in0(N__38059),
            .in1(N__35910),
            .in2(N__36564),
            .in3(N__36638),
            .lcout(\c0.n118_adj_4786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_2044_LC_5_17_5 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_2044_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_2044_LC_5_17_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i10_4_lut_adj_2044_LC_5_17_5  (
            .in0(N__35904),
            .in1(N__38060),
            .in2(N__35895),
            .in3(N__36562),
            .lcout(\c0.n63 ),
            .ltout(\c0.n63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_2016_LC_5_17_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_2016_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_2016_LC_5_17_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_4_lut_adj_2016_LC_5_17_6  (
            .in0(N__38033),
            .in1(N__35877),
            .in2(N__35841),
            .in3(N__35838),
            .lcout(\c0.n11851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_5_17_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_5_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_5_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i11_LC_5_17_7  (
            .in0(N__57977),
            .in1(N__37784),
            .in2(_gnd_net_),
            .in3(N__38061),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_5_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_5_18_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i15_LC_5_18_0  (
            .in0(N__38112),
            .in1(N__57978),
            .in2(_gnd_net_),
            .in3(N__36704),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97755),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1363_LC_5_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1363_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1363_LC_5_18_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1363_LC_5_18_1  (
            .in0(N__36021),
            .in1(N__38165),
            .in2(N__36804),
            .in3(N__35930),
            .lcout(\c0.n6_adj_4532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_adj_2043_LC_5_18_2 .C_ON=1'b0;
    defparam \c0.i4_2_lut_adj_2043_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_adj_2043_LC_5_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i4_2_lut_adj_2043_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__36636),
            .in2(_gnd_net_),
            .in3(N__36841),
            .lcout(\c0.n15_adj_4796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_2041_LC_5_18_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_2041_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_2041_LC_5_18_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i7_4_lut_adj_2041_LC_5_18_3  (
            .in0(N__36803),
            .in1(N__36824),
            .in2(N__36654),
            .in3(N__38230),
            .lcout(),
            .ltout(\c0.n18_adj_4794_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_2042_LC_5_18_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_2042_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_2042_LC_5_18_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i9_4_lut_adj_2042_LC_5_18_4  (
            .in0(N__35883),
            .in1(N__39026),
            .in2(N__35898),
            .in3(N__35957),
            .lcout(\c0.n20_adj_4795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_2032_LC_5_18_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_2032_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_2032_LC_5_18_5 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.i5_3_lut_adj_2032_LC_5_18_5  (
            .in0(N__36022),
            .in1(N__38166),
            .in2(_gnd_net_),
            .in3(N__35931),
            .lcout(\c0.n18086 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_2028_LC_5_18_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_2028_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_2028_LC_5_18_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i3_4_lut_adj_2028_LC_5_18_6  (
            .in0(N__38229),
            .in1(N__36840),
            .in2(N__36825),
            .in3(N__35956),
            .lcout(\c0.n115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_5_19_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i13_LC_5_19_0  (
            .in0(N__36799),
            .in1(N__57952),
            .in2(_gnd_net_),
            .in3(N__36555),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_5_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_5_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i32_LC_5_19_1  (
            .in0(N__80051),
            .in1(N__57966),
            .in2(_gnd_net_),
            .in3(N__36681),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_5_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_5_19_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i24_LC_5_19_2  (
            .in0(N__36682),
            .in1(N__57953),
            .in2(_gnd_net_),
            .in3(N__36023),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_5_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_5_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_5_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i16_LC_5_19_3  (
            .in0(N__36024),
            .in1(N__57965),
            .in2(_gnd_net_),
            .in3(N__35942),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_5_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_5_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i8_LC_5_19_4  (
            .in0(N__35943),
            .in1(N__57954),
            .in2(_gnd_net_),
            .in3(N__36001),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_5_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_5_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i3_LC_5_19_5  (
            .in0(N__57955),
            .in1(N__35977),
            .in2(_gnd_net_),
            .in3(N__37785),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_5_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_5_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_5_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i7_LC_5_19_6  (
            .in0(N__57964),
            .in1(N__36705),
            .in2(_gnd_net_),
            .in3(N__35958),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97769),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_2031_LC_5_19_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_2031_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_2031_LC_5_19_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i4_4_lut_adj_2031_LC_5_19_7  (
            .in0(N__36739),
            .in1(N__36854),
            .in2(N__36534),
            .in3(N__35941),
            .lcout(\c0.n10_adj_4531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rx_i_I_0_1_lut_LC_5_20_6.C_ON=1'b0;
    defparam rx_i_I_0_1_lut_LC_5_20_6.SEQ_MODE=4'b0000;
    defparam rx_i_I_0_1_lut_LC_5_20_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 rx_i_I_0_1_lut_LC_5_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38493),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_5_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_5_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_5_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i2_LC_5_20_7  (
            .in0(N__57900),
            .in1(N__36509),
            .in2(_gnd_net_),
            .in3(N__36741),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97784),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_1231_LC_6_9_2 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1231_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1231_LC_6_9_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1231_LC_6_9_2  (
            .in0(N__36926),
            .in1(N__37013),
            .in2(N__36999),
            .in3(N__36980),
            .lcout(\quad_counter0.n28_adj_4410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.quadA_I_0_85_2_lut_LC_6_9_3 .C_ON=1'b0;
    defparam \quad_counter0.quadA_I_0_85_2_lut_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.quadA_I_0_85_2_lut_LC_6_9_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter0.quadA_I_0_85_2_lut_LC_6_9_3  (
            .in0(N__37213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37166),
            .lcout(a_delay_counter_15__N_4220),
            .ltout(a_delay_counter_15__N_4220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i0_LC_6_9_4 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i0_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i0_LC_6_9_4 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \quad_counter0.a_delay_counter__i0_LC_6_9_4  (
            .in0(N__36878),
            .in1(N__37257),
            .in2(N__36114),
            .in3(N__36864),
            .lcout(a_delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97599),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_1234_LC_6_9_7 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_1234_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_1234_LC_6_9_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \quad_counter0.i9_4_lut_adj_1234_LC_6_9_7  (
            .in0(N__36947),
            .in1(N__37142),
            .in2(N__36966),
            .in3(N__36877),
            .lcout(\quad_counter0.n25_adj_4413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_6_10_0 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_6_10_0 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_6_10_0  (
            .in0(N__37593),
            .in1(N__37091),
            .in2(_gnd_net_),
            .in3(N__42721),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i3_3_lut_LC_6_11_1 .C_ON=1'b0;
    defparam \c0.tx.i3_3_lut_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i3_3_lut_LC_6_11_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i3_3_lut_LC_6_11_1  (
            .in0(N__36110),
            .in1(N__36098),
            .in2(_gnd_net_),
            .in3(N__36086),
            .lcout(),
            .ltout(\c0.n8_adj_4652_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1611_LC_6_11_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1611_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1611_LC_6_11_2 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \c0.i1_4_lut_adj_1611_LC_6_11_2  (
            .in0(N__36074),
            .in1(N__36062),
            .in2(N__36051),
            .in3(N__36270),
            .lcout(n22210),
            .ltout(n22210_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_4_lut_LC_6_11_3 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_4_lut_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_4_lut_LC_6_11_3 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \c0.tx.i1_4_lut_4_lut_LC_6_11_3  (
            .in0(N__37647),
            .in1(N__37582),
            .in2(N__36048),
            .in3(N__37435),
            .lcout(\c0.tx.n19946 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_6_11_5 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_6_11_5 .LUT_INIT=16'b0111100001010000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_6_11_5  (
            .in0(N__37090),
            .in1(N__42720),
            .in2(N__42810),
            .in3(N__37586),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_6_11_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_6_11_6 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_6_11_6  (
            .in0(N__37436),
            .in1(N__37648),
            .in2(N__37598),
            .in3(N__37479),
            .lcout(r_SM_Main_1_adj_4819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97625),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i3_4_lut_LC_6_11_7 .C_ON=1'b0;
    defparam \c0.tx.i3_4_lut_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i3_4_lut_LC_6_11_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i3_4_lut_LC_6_11_7  (
            .in0(N__36320),
            .in1(N__36308),
            .in2(N__36297),
            .in3(N__36281),
            .lcout(\c0.n47_adj_4651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_LC_6_12_0 .C_ON=1'b0;
    defparam \c0.i25_4_lut_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_LC_6_12_0 .LUT_INIT=16'b0111011110000000;
    LogicCell40 \c0.i25_4_lut_LC_6_12_0  (
            .in0(N__42729),
            .in1(N__42803),
            .in2(N__37092),
            .in3(N__36251),
            .lcout(),
            .ltout(\c0.n10_adj_4504_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_6_12_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_6_12_1 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_6_12_1  (
            .in0(N__36252),
            .in1(N__37089),
            .in2(N__36264),
            .in3(N__37594),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97639),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i34_3_lut_LC_6_12_2 .C_ON=1'b0;
    defparam \c0.i34_3_lut_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.i34_3_lut_LC_6_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i34_3_lut_LC_6_12_2  (
            .in0(N__42672),
            .in1(N__37614),
            .in2(_gnd_net_),
            .in3(N__36250),
            .lcout(\c0.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i30580_4_lut_LC_6_12_6.C_ON=1'b0;
    defparam i30580_4_lut_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam i30580_4_lut_LC_6_12_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 i30580_4_lut_LC_6_12_6 (
            .in0(N__42728),
            .in1(N__42802),
            .in2(N__37481),
            .in3(N__36249),
            .lcout(n35927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i7_LC_6_13_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_6_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_6_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__36420),
            .in2(_gnd_net_),
            .in3(N__71498),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97654),
            .ce(),
            .sr(N__36405));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_6_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_6_14_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_6_14_0  (
            .in0(N__45833),
            .in1(N__46038),
            .in2(N__36165),
            .in3(N__46181),
            .lcout(\c0.n32762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_2020_LC_6_14_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_2020_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_2020_LC_6_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_2020_LC_6_14_1  (
            .in0(N__45090),
            .in1(N__36608),
            .in2(N__36222),
            .in3(N__36191),
            .lcout(),
            .ltout(\c0.n17_adj_4788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_2021_LC_6_14_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_2021_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_2021_LC_6_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_2021_LC_6_14_2  (
            .in0(N__36161),
            .in1(N__36141),
            .in2(N__36117),
            .in3(N__36426),
            .lcout(\c0.n33160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2019_LC_6_14_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2019_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2019_LC_6_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_2019_LC_6_14_3  (
            .in0(N__36418),
            .in1(N__36494),
            .in2(N__36474),
            .in3(N__36442),
            .lcout(\c0.n16_adj_4787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1619_LC_6_14_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1619_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1619_LC_6_14_5 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1619_LC_6_14_5  (
            .in0(N__36419),
            .in1(N__45835),
            .in2(N__46060),
            .in3(N__46192),
            .lcout(\c0.n32840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1628_LC_6_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1628_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1628_LC_6_14_7 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1628_LC_6_14_7  (
            .in0(N__46182),
            .in1(N__45834),
            .in2(N__46059),
            .in3(N__37364),
            .lcout(\c0.n32718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1670_LC_6_15_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1670_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1670_LC_6_15_0 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1670_LC_6_15_0  (
            .in0(N__55231),
            .in1(N__38984),
            .in2(N__92616),
            .in3(N__48539),
            .lcout(\c0.n45_adj_4637 ),
            .ltout(\c0.n45_adj_4637_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1590_LC_6_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1590_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1590_LC_6_15_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1590_LC_6_15_1  (
            .in0(N__46047),
            .in1(N__36399),
            .in2(N__36378),
            .in3(N__46204),
            .lcout(\c0.n32714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1593_LC_6_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1593_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1593_LC_6_15_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1593_LC_6_15_3  (
            .in0(N__46046),
            .in1(N__45862),
            .in2(N__36366),
            .in3(N__46203),
            .lcout(\c0.n32804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1604_LC_6_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1604_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1604_LC_6_15_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1604_LC_6_15_4  (
            .in0(N__46206),
            .in1(N__37694),
            .in2(N__45901),
            .in3(N__46049),
            .lcout(\c0.n32798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_15_5 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_15_5 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_6_15_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_6_15_5  (
            .in0(N__71500),
            .in1(_gnd_net_),
            .in2(N__37719),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97685),
            .ce(),
            .sr(N__36330));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_6_15_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_6_15_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_6_15_6  (
            .in0(N__46205),
            .in1(N__37714),
            .in2(N__45900),
            .in3(N__46048),
            .lcout(\c0.n32712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1673_LC_6_15_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1673_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1673_LC_6_15_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1673_LC_6_15_7  (
            .in0(N__46045),
            .in1(N__36612),
            .in2(N__45895),
            .in3(N__46202),
            .lcout(\c0.n8_adj_4496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i18_LC_6_16_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_6_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_6_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__37695),
            .in2(_gnd_net_),
            .in3(N__71501),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97702),
            .ce(),
            .sr(N__36570));
    defparam \c0.data_in_0___i27_LC_6_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_6_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_6_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i27_LC_6_17_0  (
            .in0(N__80537),
            .in1(N__57971),
            .in2(_gnd_net_),
            .in3(N__38077),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_6_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_6_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_6_17_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i6_LC_6_17_3  (
            .in0(N__36721),
            .in1(_gnd_net_),
            .in2(N__57980),
            .in3(N__36639),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_6_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_6_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i5_LC_6_17_5  (
            .in0(N__57967),
            .in1(N__36563),
            .in2(_gnd_net_),
            .in3(N__36530),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97721),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30346_2_lut_LC_6_17_6 .C_ON=1'b0;
    defparam \c0.i30346_2_lut_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30346_2_lut_LC_6_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i30346_2_lut_LC_6_17_6  (
            .in0(N__36516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41149),
            .lcout(\c0.n35771 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2034_LC_6_17_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2034_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2034_LC_6_17_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_2034_LC_6_17_7  (
            .in0(N__38076),
            .in1(N__37773),
            .in2(N__36723),
            .in3(N__36515),
            .lcout(\c0.n16_adj_4790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_2030_LC_6_18_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_2030_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_2030_LC_6_18_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i3_4_lut_adj_2030_LC_6_18_0  (
            .in0(N__48713),
            .in1(N__38130),
            .in2(N__36769),
            .in3(N__42944),
            .lcout(\c0.n13_adj_4785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_6_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_6_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_6_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i18_LC_6_18_1  (
            .in0(N__57972),
            .in1(N__36762),
            .in2(_gnd_net_),
            .in3(N__48714),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i116_LC_6_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i116_LC_6_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i116_LC_6_18_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i116_LC_6_18_2  (
            .in0(N__89796),
            .in1(N__58437),
            .in2(N__52477),
            .in3(N__78908),
            .lcout(\c0.data_in_frame_14_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_2023_LC_6_18_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_2023_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_2023_LC_6_18_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i5_4_lut_adj_2023_LC_6_18_3  (
            .in0(N__36703),
            .in1(N__36684),
            .in2(N__38010),
            .in3(N__36722),
            .lcout(\c0.n12_adj_4789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_2035_LC_6_18_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_2035_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_2035_LC_6_18_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i7_4_lut_adj_2035_LC_6_18_4  (
            .in0(N__41150),
            .in1(N__38202),
            .in2(N__38267),
            .in3(N__36702),
            .lcout(),
            .ltout(\c0.n17_adj_4791_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_2036_LC_6_18_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_2036_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_2036_LC_6_18_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i9_4_lut_adj_2036_LC_6_18_5  (
            .in0(N__38107),
            .in1(N__36683),
            .in2(N__36663),
            .in3(N__36660),
            .lcout(\c0.n18094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_6_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_6_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_6_18_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i31_LC_6_18_7  (
            .in0(N__38131),
            .in1(_gnd_net_),
            .in2(N__57981),
            .in3(N__73522),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_6_19_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_6_19_0  (
            .in0(N__36890),
            .in1(N__80519),
            .in2(N__55935),
            .in3(N__46667),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i23039_2_lut_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.rx.i23039_2_lut_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i23039_2_lut_LC_6_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i23039_2_lut_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(N__55458),
            .in2(_gnd_net_),
            .in3(N__55562),
            .lcout(n27744),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_6_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_6_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i14_LC_6_19_3  (
            .in0(N__57958),
            .in1(N__36637),
            .in2(_gnd_net_),
            .in3(N__41151),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_6_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i25_LC_6_19_4  (
            .in0(N__80923),
            .in1(N__57962),
            .in2(_gnd_net_),
            .in3(N__38234),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_6_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_6_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_6_19_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i1_LC_6_19_5  (
            .in0(N__36843),
            .in1(_gnd_net_),
            .in2(N__57979),
            .in3(N__36855),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_6_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_6_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_6_19_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i9_LC_6_19_6  (
            .in0(N__38209),
            .in1(N__57963),
            .in2(_gnd_net_),
            .in3(N__36842),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i37_LC_6_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i37_LC_6_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i37_LC_6_19_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i37_LC_6_19_7  (
            .in0(N__73942),
            .in1(N__83967),
            .in2(N__39214),
            .in3(N__84031),
            .lcout(\c0.data_in_frame_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97756),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_105_i4_2_lut_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.rx.equal_105_i4_2_lut_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_105_i4_2_lut_LC_6_20_0 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \c0.rx.equal_105_i4_2_lut_LC_6_20_0  (
            .in0(N__55448),
            .in1(N__55558),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n4_adj_4808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_6_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_6_20_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i4_LC_6_20_1  (
            .in0(N__38271),
            .in1(N__57913),
            .in2(_gnd_net_),
            .in3(N__36820),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_6_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_6_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i21_LC_6_20_2  (
            .in0(N__57912),
            .in1(N__36798),
            .in2(_gnd_net_),
            .in3(N__38159),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_6_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_6_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_6_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i10_LC_6_20_4  (
            .in0(N__57911),
            .in1(N__36773),
            .in2(_gnd_net_),
            .in3(N__36740),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_6_20_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_6_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_6_20_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_6_20_5  (
            .in0(N__39170),
            .in1(N__84029),
            .in2(N__55933),
            .in3(N__46665),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i78_LC_6_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i78_LC_6_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i78_LC_6_20_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i78_LC_6_20_6  (
            .in0(N__74893),
            .in1(N__58300),
            .in2(N__87300),
            .in3(N__41600),
            .lcout(\c0.data_in_frame_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_6_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_6_20_7 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_6_20_7  (
            .in0(N__73480),
            .in1(N__36905),
            .in2(N__55934),
            .in3(N__46666),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97770),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i147_LC_6_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i147_LC_6_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i147_LC_6_21_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i147_LC_6_21_0  (
            .in0(N__80617),
            .in1(N__80362),
            .in2(N__47300),
            .in3(N__73050),
            .lcout(\c0.data_in_frame_18_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_6_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_6_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_6_21_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i28_LC_6_21_1  (
            .in0(N__78801),
            .in1(N__57976),
            .in2(_gnd_net_),
            .in3(N__38323),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i102_LC_6_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i102_LC_6_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i102_LC_6_21_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i102_LC_6_21_2  (
            .in0(N__58411),
            .in1(N__73922),
            .in2(N__49858),
            .in3(N__74895),
            .lcout(\c0.data_in_frame_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i104_LC_6_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i104_LC_6_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i104_LC_6_21_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i104_LC_6_21_3  (
            .in0(N__79960),
            .in1(N__58412),
            .in2(N__73947),
            .in3(N__41719),
            .lcout(\c0.data_in_frame_12_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_21_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_6_21_4  (
            .in0(N__52543),
            .in1(N__36909),
            .in2(N__55928),
            .in3(N__79961),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i57_LC_6_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i57_LC_6_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i57_LC_6_21_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i57_LC_6_21_5  (
            .in0(N__62266),
            .in1(N__83974),
            .in2(N__38925),
            .in3(N__80953),
            .lcout(\c0.data_in_frame_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_6_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_6_21_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_6_21_6  (
            .in0(N__52542),
            .in1(N__39174),
            .in2(N__55927),
            .in3(N__74894),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_6_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_6_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_6_21_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_6_21_7  (
            .in0(N__36891),
            .in1(N__55898),
            .in2(N__78851),
            .in3(N__52544),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97785),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_97_2_lut_LC_7_9_0 .C_ON=1'b1;
    defparam \quad_counter0.add_97_2_lut_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_97_2_lut_LC_7_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_97_2_lut_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__36879),
            .in2(_gnd_net_),
            .in3(N__36858),
            .lcout(n39),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\quad_counter0.n30016 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_delay_counter__i1_LC_7_9_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i1_LC_7_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i1_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__37014),
            .in2(_gnd_net_),
            .in3(N__37002),
            .lcout(\quad_counter0.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n30016 ),
            .carryout(\quad_counter0.n30017 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i2_LC_7_9_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i2_LC_7_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__36998),
            .in2(_gnd_net_),
            .in3(N__36984),
            .lcout(\quad_counter0.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n30017 ),
            .carryout(\quad_counter0.n30018 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i3_LC_7_9_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i3_LC_7_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i3_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__36981),
            .in2(_gnd_net_),
            .in3(N__36969),
            .lcout(\quad_counter0.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n30018 ),
            .carryout(\quad_counter0.n30019 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i4_LC_7_9_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i4_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i4_LC_7_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i4_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__36965),
            .in2(_gnd_net_),
            .in3(N__36951),
            .lcout(\quad_counter0.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n30019 ),
            .carryout(\quad_counter0.n30020 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i5_LC_7_9_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i5_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i5_LC_7_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i5_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__36948),
            .in2(_gnd_net_),
            .in3(N__36936),
            .lcout(\quad_counter0.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n30020 ),
            .carryout(\quad_counter0.n30021 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i6_LC_7_9_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i6_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i6_LC_7_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i6_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__37319),
            .in2(_gnd_net_),
            .in3(N__36933),
            .lcout(\quad_counter0.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n30021 ),
            .carryout(\quad_counter0.n30022 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i7_LC_7_9_7 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i7_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i7_LC_7_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i7_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__37028),
            .in2(_gnd_net_),
            .in3(N__36930),
            .lcout(\quad_counter0.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n30022 ),
            .carryout(\quad_counter0.n30023 ),
            .clk(N__97591),
            .ce(N__37256),
            .sr(N__37115));
    defparam \quad_counter0.a_delay_counter__i8_LC_7_10_0 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i8_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i8_LC_7_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i8_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__36927),
            .in2(_gnd_net_),
            .in3(N__36915),
            .lcout(\quad_counter0.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\quad_counter0.n30024 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i9_LC_7_10_1 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i9_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i9_LC_7_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i9_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__37335),
            .in2(_gnd_net_),
            .in3(N__36912),
            .lcout(\quad_counter0.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n30024 ),
            .carryout(\quad_counter0.n30025 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i10_LC_7_10_2 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i10_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i10_LC_7_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i10_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__37068),
            .in2(_gnd_net_),
            .in3(N__37146),
            .lcout(\quad_counter0.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n30025 ),
            .carryout(\quad_counter0.n30026 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i11_LC_7_10_3 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i11_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i11_LC_7_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i11_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__37143),
            .in2(_gnd_net_),
            .in3(N__37131),
            .lcout(\quad_counter0.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n30026 ),
            .carryout(\quad_counter0.n30027 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i12_LC_7_10_4 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i12_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i12_LC_7_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i12_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__37305),
            .in2(_gnd_net_),
            .in3(N__37128),
            .lcout(\quad_counter0.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n30027 ),
            .carryout(\quad_counter0.n30028 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i13_LC_7_10_5 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i13_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i13_LC_7_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i13_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__37347),
            .in2(_gnd_net_),
            .in3(N__37125),
            .lcout(\quad_counter0.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n30028 ),
            .carryout(\quad_counter0.n30029 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i14_LC_7_10_6 .C_ON=1'b1;
    defparam \quad_counter0.a_delay_counter__i14_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i14_LC_7_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i14_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__37056),
            .in2(_gnd_net_),
            .in3(N__37122),
            .lcout(\quad_counter0.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n30029 ),
            .carryout(\quad_counter0.n30030 ),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \quad_counter0.a_delay_counter__i15_LC_7_10_7 .C_ON=1'b0;
    defparam \quad_counter0.a_delay_counter__i15_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_delay_counter__i15_LC_7_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.a_delay_counter__i15_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__37043),
            .in2(_gnd_net_),
            .in3(N__37119),
            .lcout(\quad_counter0.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97600),
            .ce(N__37255),
            .sr(N__37116));
    defparam \c0.tx.r_SM_Main_i2_LC_7_11_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_7_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_7_11_0  (
            .in0(N__37439),
            .in1(N__37588),
            .in2(N__37480),
            .in3(N__37646),
            .lcout(r_SM_Main_2_adj_4818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97612),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_4_lut_LC_7_11_1 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_4_lut_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_4_lut_LC_7_11_1 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \c0.tx.i2_4_lut_4_lut_LC_7_11_1  (
            .in0(N__37587),
            .in1(N__37438),
            .in2(N__37650),
            .in3(N__37469),
            .lcout(\c0.n19530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1233_LC_7_11_3 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1233_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1233_LC_7_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1233_LC_7_11_3  (
            .in0(N__37067),
            .in1(N__37055),
            .in2(N__37044),
            .in3(N__37029),
            .lcout(\quad_counter0.n27_adj_4412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1353_1_lut_LC_7_11_4 .C_ON=1'b0;
    defparam \c0.tx.i1353_1_lut_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1353_1_lut_LC_7_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx.i1353_1_lut_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37642),
            .lcout(n19509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_7_11_5 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_7_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i1_2_lut_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__37437),
            .in2(_gnd_net_),
            .in3(N__37468),
            .lcout(\c0.tx.n22211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1232_LC_7_11_6 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1232_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1232_LC_7_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1232_LC_7_11_6  (
            .in0(N__37346),
            .in1(N__37334),
            .in2(N__37323),
            .in3(N__37304),
            .lcout(),
            .ltout(\quad_counter0.n26_adj_4411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_adj_1235_LC_7_11_7 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_adj_1235_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_adj_1235_LC_7_11_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_adj_1235_LC_7_11_7  (
            .in0(N__37293),
            .in1(N__37284),
            .in2(N__37278),
            .in3(N__37275),
            .lcout(n15010),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_1333_LC_7_12_1 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_1333_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_1333_LC_7_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_1333_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__37430),
            .in2(_gnd_net_),
            .in3(N__48289),
            .lcout(),
            .ltout(\c0.tx.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_LC_7_12_2 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_LC_7_12_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \c0.tx.i2_4_lut_LC_7_12_2  (
            .in0(N__37592),
            .in1(N__37501),
            .in2(N__37266),
            .in3(N__37263),
            .lcout(\c0.tx.n19358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_2061_LC_7_12_4.C_ON=1'b0;
    defparam i1_3_lut_adj_2061_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_2061_LC_7_12_4.LUT_INIT=16'b1111111101100110;
    LogicCell40 i1_3_lut_adj_2061_LC_7_12_4 (
            .in0(N__37223),
            .in1(N__37172),
            .in2(_gnd_net_),
            .in3(N__37181),
            .lcout(n19493),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_72_LC_7_12_6 .C_ON=1'b0;
    defparam \quad_counter0.A_72_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_72_LC_7_12_6 .LUT_INIT=16'b1111001011100000;
    LogicCell40 \quad_counter0.A_72_LC_7_12_6  (
            .in0(N__37224),
            .in1(N__37182),
            .in2(N__39295),
            .in3(N__37173),
            .lcout(A_filtered),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97626),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_4_lut_LC_7_13_2 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_4_lut_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_4_lut_LC_7_13_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i2_3_lut_4_lut_LC_7_13_2  (
            .in0(N__37417),
            .in1(N__37649),
            .in2(N__48294),
            .in3(N__37595),
            .lcout(n14821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_7_13_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_7_13_3 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_7_13_3  (
            .in0(N__42966),
            .in1(N__42808),
            .in2(N__42746),
            .in3(N__55143),
            .lcout(),
            .ltout(\c0.tx.n36215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n36215_bdd_4_lut_LC_7_13_4 .C_ON=1'b0;
    defparam \c0.tx.n36215_bdd_4_lut_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n36215_bdd_4_lut_LC_7_13_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.tx.n36215_bdd_4_lut_LC_7_13_4  (
            .in0(N__42809),
            .in1(N__55011),
            .in2(N__37617),
            .in3(N__42900),
            .lcout(\c0.n36218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_7_13_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_7_13_5 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_7_13_5  (
            .in0(N__37597),
            .in1(N__48221),
            .in2(_gnd_net_),
            .in3(N__37608),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97640),
            .ce(),
            .sr(_gnd_net_));
    defparam i26_3_lut_LC_7_13_6.C_ON=1'b0;
    defparam i26_3_lut_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam i26_3_lut_LC_7_13_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 i26_3_lut_LC_7_13_6 (
            .in0(N__48293),
            .in1(N__37596),
            .in2(_gnd_net_),
            .in3(N__37533),
            .lcout(),
            .ltout(n9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_7_13_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_7_13_7 .LUT_INIT=16'b0100000011001000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_7_13_7  (
            .in0(N__37434),
            .in1(N__37512),
            .in2(N__37485),
            .in3(N__37482),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97640),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1591_LC_7_14_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1591_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1591_LC_7_14_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i1_2_lut_adj_1591_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__48345),
            .in2(_gnd_net_),
            .in3(N__48480),
            .lcout(\c0.n6_adj_4638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2017_LC_7_14_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2017_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2017_LC_7_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_2017_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__37389),
            .in2(_gnd_net_),
            .in3(N__37360),
            .lcout(\c0.n19546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i31_LC_7_14_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_7_14_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_7_14_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_7_14_4  (
            .in0(N__71446),
            .in1(_gnd_net_),
            .in2(N__37365),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97655),
            .ce(),
            .sr(N__37752));
    defparam \c0.select_369_Select_7_i3_2_lut_LC_7_14_6 .C_ON=1'b0;
    defparam \c0.select_369_Select_7_i3_2_lut_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_7_i3_2_lut_LC_7_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_7_i3_2_lut_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__91713),
            .in2(_gnd_net_),
            .in3(N__94699),
            .lcout(\c0.n3_adj_4586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1674_LC_7_15_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1674_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1674_LC_7_15_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1674_LC_7_15_0  (
            .in0(N__45836),
            .in1(N__46061),
            .in2(N__37671),
            .in3(N__46191),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1950_LC_7_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1950_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1950_LC_7_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_1950_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__51836),
            .in2(_gnd_net_),
            .in3(N__51591),
            .lcout(\c0.n79 ),
            .ltout(\c0.n79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1725_LC_7_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1725_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1725_LC_7_15_2 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1725_LC_7_15_2  (
            .in0(N__49185),
            .in1(N__48531),
            .in2(N__37740),
            .in3(N__51561),
            .lcout(\c0.data_out_frame_0__7__N_2568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1675_LC_7_15_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1675_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1675_LC_7_15_3 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1675_LC_7_15_3  (
            .in0(N__48447),
            .in1(N__48490),
            .in2(_gnd_net_),
            .in3(N__48190),
            .lcout(),
            .ltout(\c0.n4_adj_4613_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1518_LC_7_15_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1518_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1518_LC_7_15_4 .LUT_INIT=16'b1010000010101000;
    LogicCell40 \c0.i1_4_lut_adj_1518_LC_7_15_4  (
            .in0(N__51837),
            .in1(N__51520),
            .in2(N__37737),
            .in3(N__55370),
            .lcout(\c0.n11_adj_4614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_15_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_15_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_7_15_6  (
            .in0(N__37670),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71447),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97668),
            .ce(),
            .sr(N__37734));
    defparam \c0.i1_2_lut_4_lut_adj_1334_LC_7_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1334_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1334_LC_7_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1334_LC_7_16_0  (
            .in0(N__37693),
            .in1(N__37666),
            .in2(N__37718),
            .in3(N__37887),
            .lcout(),
            .ltout(\c0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_2046_LC_7_16_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_2046_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_2046_LC_7_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_2046_LC_7_16_1  (
            .in0(N__37902),
            .in1(N__46332),
            .in2(N__37722),
            .in3(N__37823),
            .lcout(\c0.n16_adj_4797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_7_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_7_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_7_16_2  (
            .in0(N__37710),
            .in1(N__37692),
            .in2(N__37934),
            .in3(N__37665),
            .lcout(\c0.n19820 ),
            .ltout(\c0.n19820_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1687_LC_7_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1687_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1687_LC_7_16_3 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1687_LC_7_16_3  (
            .in0(N__49237),
            .in1(N__48592),
            .in2(N__37938),
            .in3(N__49092),
            .lcout(\c0.n93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23550_3_lut_4_lut_LC_7_16_4 .C_ON=1'b0;
    defparam \c0.i23550_3_lut_4_lut_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i23550_3_lut_4_lut_LC_7_16_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \c0.i23550_3_lut_4_lut_LC_7_16_4  (
            .in0(N__37874),
            .in1(N__49091),
            .in2(N__37935),
            .in3(N__49236),
            .lcout(\c0.n27824 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2047_LC_7_16_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2047_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2047_LC_7_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_2047_LC_7_16_5  (
            .in0(N__37850),
            .in1(N__48591),
            .in2(N__46269),
            .in3(N__46308),
            .lcout(),
            .ltout(\c0.n15_adj_4798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28768_4_lut_LC_7_16_6 .C_ON=1'b0;
    defparam \c0.i28768_4_lut_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i28768_4_lut_LC_7_16_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i28768_4_lut_LC_7_16_6  (
            .in0(N__71270),
            .in1(N__37896),
            .in2(N__37890),
            .in3(N__48540),
            .lcout(\c0.n34190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1943_LC_7_16_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1943_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1943_LC_7_16_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1943_LC_7_16_7  (
            .in0(N__37886),
            .in1(N__37873),
            .in2(N__37851),
            .in3(N__37822),
            .lcout(\c0.n30958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2024_LC_7_17_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2024_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2024_LC_7_17_0 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i6_4_lut_adj_2024_LC_7_17_0  (
            .in0(N__38078),
            .in1(N__38210),
            .in2(N__38108),
            .in3(N__37800),
            .lcout(),
            .ltout(\c0.n35698_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_2025_LC_7_17_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_2025_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_2025_LC_7_17_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.i4_4_lut_adj_2025_LC_7_17_1  (
            .in0(N__37794),
            .in1(N__38262),
            .in2(N__37788),
            .in3(N__37783),
            .lcout(\c0.n33263 ),
            .ltout(\c0.n33263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23120_2_lut_3_lut_4_lut_LC_7_17_2 .C_ON=1'b0;
    defparam \c0.i23120_2_lut_3_lut_4_lut_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i23120_2_lut_3_lut_4_lut_LC_7_17_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i23120_2_lut_3_lut_4_lut_LC_7_17_2  (
            .in0(N__37976),
            .in1(N__37957),
            .in2(N__37755),
            .in3(N__46231),
            .lcout(\c0.data_out_frame_29_7_N_1483_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2033_LC_7_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2033_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2033_LC_7_17_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_2033_LC_7_17_3  (
            .in0(N__37956),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37975),
            .lcout(\c0.n29676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_7_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_7_17_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i23_LC_7_17_4  (
            .in0(N__38103),
            .in1(_gnd_net_),
            .in2(N__57957),
            .in3(N__38135),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97703),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_7_17_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_7_17_5 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_7_17_5  (
            .in0(N__38040),
            .in1(N__38022),
            .in2(N__38808),
            .in3(N__38008),
            .lcout(\c0.data_out_frame_29_7_N_2879_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_7_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_7_17_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i19_LC_7_17_6  (
            .in0(N__38079),
            .in1(_gnd_net_),
            .in2(N__57956),
            .in3(N__38058),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97703),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_7_17_7 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_7_17_7  (
            .in0(N__38039),
            .in1(N__38021),
            .in2(N__38937),
            .in3(N__38009),
            .lcout(\c0.n22387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2051_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2051_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2051_LC_7_18_0 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_2051_LC_7_18_0  (
            .in0(N__37959),
            .in1(N__39041),
            .in2(N__37986),
            .in3(N__38962),
            .lcout(\c0.data_out_frame_29_7_N_1483_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1967_LC_7_18_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1967_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1967_LC_7_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1967_LC_7_18_1  (
            .in0(N__38179),
            .in1(N__39079),
            .in2(_gnd_net_),
            .in3(N__39241),
            .lcout(\c0.n33341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i107_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i107_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i107_LC_7_18_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i107_LC_7_18_3  (
            .in0(N__68600),
            .in1(N__78594),
            .in2(N__50062),
            .in3(N__80498),
            .lcout(\c0.data_in_frame_13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_2015_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_2015_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_2015_LC_7_18_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_2015_LC_7_18_4  (
            .in0(N__37982),
            .in1(N__39040),
            .in2(_gnd_net_),
            .in3(N__37958),
            .lcout(\c0.n29668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_7_18_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i20_LC_7_18_5  (
            .in0(N__38289),
            .in1(N__57907),
            .in2(_gnd_net_),
            .in3(N__38337),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_7_18_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i12_LC_7_18_6  (
            .in0(N__57908),
            .in1(N__38290),
            .in2(_gnd_net_),
            .in3(N__38266),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i108_LC_7_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i108_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i108_LC_7_18_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i108_LC_7_18_7  (
            .in0(N__78907),
            .in1(N__78595),
            .in2(N__68604),
            .in3(N__50011),
            .lcout(\c0.data_in_frame_13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97722),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1341_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1341_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1341_LC_7_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1341_LC_7_19_0  (
            .in0(N__38180),
            .in1(N__49365),
            .in2(N__38399),
            .in3(N__41466),
            .lcout(\c0.n9_adj_4509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_7_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i17_LC_7_19_1  (
            .in0(N__38238),
            .in1(N__57909),
            .in2(_gnd_net_),
            .in3(N__38211),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1418_LC_7_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1418_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1418_LC_7_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1418_LC_7_19_2  (
            .in0(N__44318),
            .in1(N__52519),
            .in2(_gnd_net_),
            .in3(N__38348),
            .lcout(\c0.n4_adj_4548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i72_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i72_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i72_LC_7_19_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i72_LC_7_19_3  (
            .in0(N__80052),
            .in1(N__81223),
            .in2(N__58440),
            .in3(N__44260),
            .lcout(\c0.data_in_frame_8_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i39_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i39_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i39_LC_7_19_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i39_LC_7_19_4  (
            .in0(N__83963),
            .in1(N__73523),
            .in2(N__38184),
            .in3(N__73936),
            .lcout(\c0.data_in_frame_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_7_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_7_19_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i29_LC_7_19_5  (
            .in0(N__84030),
            .in1(N__57910),
            .in2(_gnd_net_),
            .in3(N__38158),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i38_LC_7_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i38_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i38_LC_7_19_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i38_LC_7_19_6  (
            .in0(N__83962),
            .in1(N__73935),
            .in2(N__39090),
            .in3(N__75061),
            .lcout(\c0.data_in_frame_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i79_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i79_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i79_LC_7_19_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i79_LC_7_19_7  (
            .in0(N__58432),
            .in1(N__73524),
            .in2(N__38352),
            .in3(N__87274),
            .lcout(\c0.data_in_frame_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97738),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_7_20_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.i1_2_lut_LC_7_20_0  (
            .in0(N__58037),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55624),
            .lcout(n18026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_7_20_1 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_7_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_7_20_1  (
            .in0(N__41382),
            .in1(N__43356),
            .in2(N__38400),
            .in3(N__41464),
            .lcout(),
            .ltout(\c0.n8_adj_4508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1833_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1833_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1833_LC_7_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1833_LC_7_20_2  (
            .in0(N__38367),
            .in1(N__41394),
            .in2(N__38340),
            .in3(N__39246),
            .lcout(\c0.n33444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i58_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i58_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i58_LC_7_20_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \c0.data_in_frame_0__i58_LC_7_20_4  (
            .in0(N__75360),
            .in1(N__83966),
            .in2(N__62265),
            .in3(N__38424),
            .lcout(\c0.data_in_frame_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i59_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i59_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i59_LC_7_20_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i59_LC_7_20_5  (
            .in0(N__83964),
            .in1(N__62245),
            .in2(N__44139),
            .in3(N__80499),
            .lcout(\c0.data_in_frame_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_7_20_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_7_20_6  (
            .in0(N__90630),
            .in1(N__42761),
            .in2(N__71163),
            .in3(N__71662),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i60_LC_7_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i60_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i60_LC_7_20_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i60_LC_7_20_7  (
            .in0(N__83965),
            .in1(N__62246),
            .in2(N__41899),
            .in3(N__78808),
            .lcout(\c0.data_in_frame_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97757),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_7_21_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i5_LC_7_21_1  (
            .in0(N__81224),
            .in1(N__83909),
            .in2(N__43830),
            .in3(N__84032),
            .lcout(\c0.data_in_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97771),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1328_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1328_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1328_LC_7_21_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.i1_2_lut_adj_1328_LC_7_21_2  (
            .in0(N__55625),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58038),
            .lcout(n18031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1447_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1447_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1447_LC_7_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1447_LC_7_21_3  (
            .in0(N__46625),
            .in1(N__46940),
            .in2(N__38881),
            .in3(N__41965),
            .lcout(\c0.n33985 ),
            .ltout(\c0.n33985_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1825_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1825_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1825_LC_7_21_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1825_LC_7_21_4  (
            .in0(N__38423),
            .in1(_gnd_net_),
            .in2(N__38427),
            .in3(N__38409),
            .lcout(\c0.n33781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1870_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1870_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1870_LC_7_21_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1870_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__58098),
            .in2(_gnd_net_),
            .in3(N__38422),
            .lcout(\c0.n33758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1834_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1834_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1834_LC_7_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1834_LC_7_21_6  (
            .in0(N__38917),
            .in1(N__42001),
            .in2(_gnd_net_),
            .in3(N__38408),
            .lcout(\c0.n33778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i92_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i92_LC_7_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i92_LC_7_21_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i92_LC_7_21_7  (
            .in0(N__58410),
            .in1(N__78259),
            .in2(N__78852),
            .in3(N__41966),
            .lcout(\c0.data_in_frame_11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97771),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_7_22_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i41_LC_7_22_0  (
            .in0(N__80976),
            .in1(N__78581),
            .in2(N__38398),
            .in3(N__68297),
            .lcout(\c0.data_in_frame_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97786),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i75_LC_7_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i75_LC_7_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i75_LC_7_22_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i75_LC_7_22_1  (
            .in0(N__58382),
            .in1(N__87221),
            .in2(N__80618),
            .in3(N__38366),
            .lcout(\c0.data_in_frame_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97786),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1840_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1840_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1840_LC_7_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1840_LC_7_22_3  (
            .in0(N__58097),
            .in1(N__41844),
            .in2(N__46645),
            .in3(N__41558),
            .lcout(\c0.n18368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i74_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i74_LC_7_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i74_LC_7_22_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i74_LC_7_22_4  (
            .in0(N__75364),
            .in1(N__87220),
            .in2(N__38885),
            .in3(N__58383),
            .lcout(\c0.data_in_frame_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97786),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1866_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1866_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1866_LC_7_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1866_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(N__38877),
            .in2(_gnd_net_),
            .in3(N__38916),
            .lcout(\c0.n34000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3181_2_lut_LC_7_22_6 .C_ON=1'b0;
    defparam \c0.i3181_2_lut_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3181_2_lut_LC_7_22_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3181_2_lut_LC_7_22_6  (
            .in0(N__50233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41713),
            .lcout(\c0.n5860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i93_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i93_LC_7_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i93_LC_7_23_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i93_LC_7_23_1  (
            .in0(N__78260),
            .in1(N__58429),
            .in2(N__42005),
            .in3(N__84071),
            .lcout(\c0.data_in_frame_11_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i88_LC_7_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i88_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i88_LC_7_23_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i88_LC_7_23_6  (
            .in0(N__58427),
            .in1(N__80009),
            .in2(N__80396),
            .in3(N__39327),
            .lcout(\c0.data_in_frame_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i103_LC_7_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i103_LC_7_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i103_LC_7_23_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i103_LC_7_23_7  (
            .in0(N__73934),
            .in1(N__58428),
            .in2(N__50250),
            .in3(N__73545),
            .lcout(\c0.data_in_frame_12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97792),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_7_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_7_24_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i55_LC_7_24_0  (
            .in0(N__73640),
            .in1(N__83961),
            .in2(N__89808),
            .in3(N__46618),
            .lcout(\c0.data_in_frame_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97795),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i125_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i125_LC_7_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i125_LC_7_24_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i125_LC_7_24_2  (
            .in0(N__62253),
            .in1(N__58431),
            .in2(N__44110),
            .in3(N__84117),
            .lcout(\c0.data_in_frame_15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97795),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i120_LC_7_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i120_LC_7_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i120_LC_7_24_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i120_LC_7_24_4  (
            .in0(N__80008),
            .in1(N__58430),
            .in2(N__89807),
            .in3(N__44448),
            .lcout(\c0.data_in_frame_14_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97795),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_97_2_lut_LC_9_7_0 .C_ON=1'b1;
    defparam \quad_counter1.add_97_2_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_97_2_lut_LC_9_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_97_2_lut_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__39566),
            .in2(_gnd_net_),
            .in3(N__38433),
            .lcout(n39_adj_4816),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\quad_counter1.n30046 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i1_LC_9_7_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i1_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i1_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i1_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__39611),
            .in2(_gnd_net_),
            .in3(N__38430),
            .lcout(\quad_counter1.a_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n30046 ),
            .carryout(\quad_counter1.n30047 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i2_LC_9_7_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i2_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i2_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i2_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__39624),
            .in2(_gnd_net_),
            .in3(N__38460),
            .lcout(\quad_counter1.a_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n30047 ),
            .carryout(\quad_counter1.n30048 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i3_LC_9_7_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i3_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i3_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i3_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__39548),
            .in2(_gnd_net_),
            .in3(N__38457),
            .lcout(\quad_counter1.a_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n30048 ),
            .carryout(\quad_counter1.n30049 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i4_LC_9_7_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i4_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i4_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i4_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__39534),
            .in2(_gnd_net_),
            .in3(N__38454),
            .lcout(\quad_counter1.a_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n30049 ),
            .carryout(\quad_counter1.n30050 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i5_LC_9_7_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i5_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i5_LC_9_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i5_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__39597),
            .in2(_gnd_net_),
            .in3(N__38451),
            .lcout(\quad_counter1.a_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n30050 ),
            .carryout(\quad_counter1.n30051 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i6_LC_9_7_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i6_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i6_LC_9_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i6_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__39738),
            .in2(_gnd_net_),
            .in3(N__38448),
            .lcout(\quad_counter1.a_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n30051 ),
            .carryout(\quad_counter1.n30052 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i7_LC_9_7_7 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i7_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i7_LC_9_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i7_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__39510),
            .in2(_gnd_net_),
            .in3(N__38445),
            .lcout(\quad_counter1.a_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n30052 ),
            .carryout(\quad_counter1.n30053 ),
            .clk(N__97560),
            .ce(N__39768),
            .sr(N__39668));
    defparam \quad_counter1.a_delay_counter__i8_LC_9_8_0 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i8_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i8_LC_9_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i8_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__39708),
            .in2(_gnd_net_),
            .in3(N__38442),
            .lcout(\quad_counter1.a_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\quad_counter1.n30054 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i9_LC_9_8_1 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i9_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i9_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i9_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__39585),
            .in2(_gnd_net_),
            .in3(N__38439),
            .lcout(\quad_counter1.a_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n30054 ),
            .carryout(\quad_counter1.n30055 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i10_LC_9_8_2 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i10_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i10_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i10_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__39722),
            .in2(_gnd_net_),
            .in3(N__38436),
            .lcout(\quad_counter1.a_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n30055 ),
            .carryout(\quad_counter1.n30056 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i11_LC_9_8_3 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i11_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i11_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i11_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__39750),
            .in2(_gnd_net_),
            .in3(N__38508),
            .lcout(\quad_counter1.a_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n30056 ),
            .carryout(\quad_counter1.n30057 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i12_LC_9_8_4 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i12_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i12_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i12_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__39497),
            .in2(_gnd_net_),
            .in3(N__38505),
            .lcout(\quad_counter1.a_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n30057 ),
            .carryout(\quad_counter1.n30058 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i13_LC_9_8_5 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i13_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i13_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i13_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__39636),
            .in2(_gnd_net_),
            .in3(N__38502),
            .lcout(\quad_counter1.a_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n30058 ),
            .carryout(\quad_counter1.n30059 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i14_LC_9_8_6 .C_ON=1'b1;
    defparam \quad_counter1.a_delay_counter__i14_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i14_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i14_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__39522),
            .in2(_gnd_net_),
            .in3(N__38499),
            .lcout(\quad_counter1.a_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n30059 ),
            .carryout(\quad_counter1.n30060 ),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \quad_counter1.a_delay_counter__i15_LC_9_8_7 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i15_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i15_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.a_delay_counter__i15_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__39483),
            .in2(_gnd_net_),
            .in3(N__38496),
            .lcout(\quad_counter1.a_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97567),
            .ce(N__39767),
            .sr(N__39669));
    defparam \c0.rx.r_Rx_Data_R_49_LC_9_9_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_R_49_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_R_49_LC_9_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_R_49_LC_9_9_4  (
            .in0(N__38483),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_Rx_Data_R ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97576),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1173_LC_9_9_5 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1173_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1173_LC_9_9_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1173_LC_9_9_5  (
            .in0(N__40257),
            .in1(N__40201),
            .in2(N__42291),
            .in3(N__40461),
            .lcout(\quad_counter0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_1182_LC_9_10_0 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_1182_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_1182_LC_9_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i9_4_lut_adj_1182_LC_9_10_0  (
            .in0(N__44719),
            .in1(N__44983),
            .in2(N__44776),
            .in3(N__47781),
            .lcout(),
            .ltout(\quad_counter0.n25_adj_4367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_adj_1183_LC_9_10_1 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_adj_1183_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_adj_1183_LC_9_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_adj_1183_LC_9_10_1  (
            .in0(N__38547),
            .in1(N__38553),
            .in2(N__38463),
            .in3(N__38541),
            .lcout(\quad_counter0.n3332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1181_LC_9_10_2 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1181_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1181_LC_9_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1181_LC_9_10_2  (
            .in0(N__45007),
            .in1(N__44884),
            .in2(N__44866),
            .in3(N__45259),
            .lcout(\quad_counter0.n27_adj_4366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_1179_LC_9_10_3 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1179_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1179_LC_9_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1179_LC_9_10_3  (
            .in0(N__44906),
            .in1(N__44741),
            .in2(N__44701),
            .in3(N__45283),
            .lcout(\quad_counter0.n28_adj_4364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1180_LC_9_10_5 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1180_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1180_LC_9_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1180_LC_9_10_5  (
            .in0(N__44959),
            .in1(N__44935),
            .in2(N__45040),
            .in3(N__45235),
            .lcout(\quad_counter0.n26_adj_4365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_1174_LC_9_11_0 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_1174_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_1174_LC_9_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i9_4_lut_adj_1174_LC_9_11_0  (
            .in0(N__40597),
            .in1(N__40105),
            .in2(N__40713),
            .in3(N__40639),
            .lcout(\quad_counter0.n24_adj_4360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i13_4_lut_adj_1175_LC_9_11_1 .C_ON=1'b0;
    defparam \quad_counter0.i13_4_lut_adj_1175_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i13_4_lut_adj_1175_LC_9_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i13_4_lut_adj_1175_LC_9_11_1  (
            .in0(N__40015),
            .in1(N__40405),
            .in2(N__39816),
            .in3(N__38535),
            .lcout(),
            .ltout(\quad_counter0.n28_adj_4361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i14_4_lut_LC_9_11_2 .C_ON=1'b0;
    defparam \quad_counter0.i14_4_lut_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i14_4_lut_LC_9_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i14_4_lut_LC_9_11_2  (
            .in0(N__40917),
            .in1(N__39807),
            .in2(N__38526),
            .in3(N__38523),
            .lcout(\quad_counter0.n3233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30716_1_lut_LC_9_11_3 .C_ON=1'b0;
    defparam \quad_counter0.i30716_1_lut_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30716_1_lut_LC_9_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30716_1_lut_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40758),
            .lcout(\quad_counter0.n36143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_9_11_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_9_11_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_9_11_4  (
            .in0(N__38517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97592),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__7__5446_LC_9_11_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__7__5446_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__7__5446_LC_9_11_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_9__7__5446_LC_9_11_5  (
            .in0(N__85230),
            .in1(N__84703),
            .in2(N__75948),
            .in3(N__57566),
            .lcout(data_out_frame_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97592),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_2_lut_LC_9_12_0 .C_ON=1'b0;
    defparam \quad_counter0.i4_2_lut_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_2_lut_LC_9_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i4_2_lut_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__40575),
            .in2(_gnd_net_),
            .in3(N__40887),
            .lcout(),
            .ltout(\quad_counter0.n18_adj_4353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_1170_LC_9_12_1 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1170_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1170_LC_9_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1170_LC_9_12_1  (
            .in0(N__40344),
            .in1(N__40668),
            .in2(N__38583),
            .in3(N__38718),
            .lcout(\quad_counter0.n26_adj_4356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_3_lut_LC_9_12_2 .C_ON=1'b0;
    defparam \quad_counter0.i1_3_lut_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_3_lut_LC_9_12_2 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \quad_counter0.i1_3_lut_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__59845),
            .in2(N__40281),
            .in3(N__40300),
            .lcout(),
            .ltout(\quad_counter0.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1167_LC_9_12_3 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1167_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1167_LC_9_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1167_LC_9_12_3  (
            .in0(N__40216),
            .in1(N__40174),
            .in2(N__38580),
            .in3(N__70647),
            .lcout(),
            .ltout(\quad_counter0.n34617_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_adj_1169_LC_9_12_4 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_adj_1169_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_adj_1169_LC_9_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_adj_1169_LC_9_12_4  (
            .in0(N__40386),
            .in1(N__40081),
            .in2(N__38577),
            .in3(N__40845),
            .lcout(),
            .ltout(\quad_counter0.n22_adj_4355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i13_4_lut_LC_9_12_5 .C_ON=1'b0;
    defparam \quad_counter0.i13_4_lut_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i13_4_lut_LC_9_12_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i13_4_lut_LC_9_12_5  (
            .in0(N__40036),
            .in1(N__40620),
            .in2(N__38574),
            .in3(N__38571),
            .lcout(\quad_counter0.n3134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_2_lut_LC_9_13_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_2_lut_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_2_lut_LC_9_13_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2085_2_lut_LC_9_13_0  (
            .in0(N__59811),
            .in1(N__59810),
            .in2(N__38758),
            .in3(N__38565),
            .lcout(\quad_counter0.n3119 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\quad_counter0.n30347 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_3_lut_LC_9_13_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_3_lut_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_3_lut_LC_9_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_3_lut_LC_9_13_1  (
            .in0(N__42842),
            .in1(N__42841),
            .in2(N__38708),
            .in3(N__38562),
            .lcout(\quad_counter0.n3118 ),
            .ltout(),
            .carryin(\quad_counter0.n30347 ),
            .carryout(\quad_counter0.n30348 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_4_lut_LC_9_13_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_4_lut_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_4_lut_LC_9_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2085_4_lut_LC_9_13_2  (
            .in0(N__42639),
            .in1(N__42638),
            .in2(N__38759),
            .in3(N__38559),
            .lcout(\quad_counter0.n3117 ),
            .ltout(),
            .carryin(\quad_counter0.n30348 ),
            .carryout(\quad_counter0.n30349 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_5_lut_LC_9_13_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_5_lut_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_5_lut_LC_9_13_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2085_5_lut_LC_9_13_3  (
            .in0(N__42590),
            .in1(N__42589),
            .in2(N__38762),
            .in3(N__38556),
            .lcout(\quad_counter0.n3116 ),
            .ltout(),
            .carryin(\quad_counter0.n30349 ),
            .carryout(\quad_counter0.n30350 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_6_lut_LC_9_13_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_6_lut_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_6_lut_LC_9_13_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2085_6_lut_LC_9_13_4  (
            .in0(N__41118),
            .in1(N__41117),
            .in2(N__38760),
            .in3(N__38610),
            .lcout(\quad_counter0.n3115 ),
            .ltout(),
            .carryin(\quad_counter0.n30350 ),
            .carryout(\quad_counter0.n30351 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_7_lut_LC_9_13_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_7_lut_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_7_lut_LC_9_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2085_7_lut_LC_9_13_5  (
            .in0(N__41088),
            .in1(N__41087),
            .in2(N__38763),
            .in3(N__38607),
            .lcout(\quad_counter0.n3114 ),
            .ltout(),
            .carryin(\quad_counter0.n30351 ),
            .carryout(\quad_counter0.n30352 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_8_lut_LC_9_13_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_8_lut_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_8_lut_LC_9_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2085_8_lut_LC_9_13_6  (
            .in0(N__42615),
            .in1(N__42614),
            .in2(N__38761),
            .in3(N__38604),
            .lcout(\quad_counter0.n3113 ),
            .ltout(),
            .carryin(\quad_counter0.n30352 ),
            .carryout(\quad_counter0.n30353 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_9_lut_LC_9_13_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_9_lut_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_9_lut_LC_9_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_9_lut_LC_9_13_7  (
            .in0(N__41061),
            .in1(N__41057),
            .in2(N__38709),
            .in3(N__38601),
            .lcout(\quad_counter0.n3112 ),
            .ltout(),
            .carryin(\quad_counter0.n30353 ),
            .carryout(\quad_counter0.n30354 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_10_lut_LC_9_14_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_10_lut_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_10_lut_LC_9_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_10_lut_LC_9_14_0  (
            .in0(N__41031),
            .in1(N__41030),
            .in2(N__38699),
            .in3(N__38598),
            .lcout(\quad_counter0.n3111 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\quad_counter0.n30355 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_11_lut_LC_9_14_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_11_lut_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_11_lut_LC_9_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_11_lut_LC_9_14_1  (
            .in0(N__41010),
            .in1(N__41009),
            .in2(N__38703),
            .in3(N__38595),
            .lcout(\quad_counter0.n3110 ),
            .ltout(),
            .carryin(\quad_counter0.n30355 ),
            .carryout(\quad_counter0.n30356 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_12_lut_LC_9_14_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_12_lut_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_12_lut_LC_9_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_12_lut_LC_9_14_2  (
            .in0(N__40986),
            .in1(N__40985),
            .in2(N__38700),
            .in3(N__38592),
            .lcout(\quad_counter0.n3109 ),
            .ltout(),
            .carryin(\quad_counter0.n30356 ),
            .carryout(\quad_counter0.n30357 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_13_lut_LC_9_14_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_13_lut_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_13_lut_LC_9_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_13_lut_LC_9_14_3  (
            .in0(N__40959),
            .in1(N__40958),
            .in2(N__38704),
            .in3(N__38589),
            .lcout(\quad_counter0.n3108 ),
            .ltout(),
            .carryin(\quad_counter0.n30357 ),
            .carryout(\quad_counter0.n30358 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_14_lut_LC_9_14_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_14_lut_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_14_lut_LC_9_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_14_lut_LC_9_14_4  (
            .in0(N__41343),
            .in1(N__41342),
            .in2(N__38701),
            .in3(N__38586),
            .lcout(\quad_counter0.n3107 ),
            .ltout(),
            .carryin(\quad_counter0.n30358 ),
            .carryout(\quad_counter0.n30359 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_15_lut_LC_9_14_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_15_lut_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_15_lut_LC_9_14_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_15_lut_LC_9_14_5  (
            .in0(N__41316),
            .in1(N__41315),
            .in2(N__38705),
            .in3(N__38781),
            .lcout(\quad_counter0.n3106 ),
            .ltout(),
            .carryin(\quad_counter0.n30359 ),
            .carryout(\quad_counter0.n30360 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_16_lut_LC_9_14_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_16_lut_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_16_lut_LC_9_14_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_16_lut_LC_9_14_6  (
            .in0(N__41289),
            .in1(N__41288),
            .in2(N__38702),
            .in3(N__38778),
            .lcout(\quad_counter0.n3105 ),
            .ltout(),
            .carryin(\quad_counter0.n30360 ),
            .carryout(\quad_counter0.n30361 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_17_lut_LC_9_14_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_17_lut_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_17_lut_LC_9_14_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_17_lut_LC_9_14_7  (
            .in0(N__41265),
            .in1(N__41261),
            .in2(N__38706),
            .in3(N__38775),
            .lcout(\quad_counter0.n3104 ),
            .ltout(),
            .carryin(\quad_counter0.n30361 ),
            .carryout(\quad_counter0.n30362 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_18_lut_LC_9_15_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_18_lut_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_18_lut_LC_9_15_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_18_lut_LC_9_15_0  (
            .in0(N__41232),
            .in1(N__41228),
            .in2(N__38691),
            .in3(N__38772),
            .lcout(\quad_counter0.n3103 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\quad_counter0.n30363 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_19_lut_LC_9_15_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2085_19_lut_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_19_lut_LC_9_15_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_19_lut_LC_9_15_1  (
            .in0(N__41204),
            .in1(N__41205),
            .in2(N__38707),
            .in3(N__38769),
            .lcout(\quad_counter0.n3102 ),
            .ltout(),
            .carryin(\quad_counter0.n30363 ),
            .carryout(\quad_counter0.n30364 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2085_20_lut_LC_9_15_2 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_2085_20_lut_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2085_20_lut_LC_9_15_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2085_20_lut_LC_9_15_2  (
            .in0(N__41174),
            .in1(N__41175),
            .in2(N__38692),
            .in3(N__38766),
            .lcout(\quad_counter0.n3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30717_1_lut_LC_9_15_3 .C_ON=1'b0;
    defparam \quad_counter0.i30717_1_lut_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30717_1_lut_LC_9_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30717_1_lut_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38652),
            .lcout(\quad_counter0.n36144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1168_LC_9_15_4 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1168_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1168_LC_9_15_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1168_LC_9_15_4  (
            .in0(N__40525),
            .in1(N__40426),
            .in2(N__40482),
            .in3(N__40933),
            .lcout(\quad_counter0.n24_adj_4354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_1166_LC_9_15_5 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1166_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1166_LC_9_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1166_LC_9_15_5  (
            .in0(N__41050),
            .in1(N__40978),
            .in2(N__38844),
            .in3(N__38826),
            .lcout(\quad_counter0.n3035 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_adj_1164_LC_9_15_6 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_adj_1164_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_adj_1164_LC_9_15_6 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \quad_counter0.i3_4_lut_adj_1164_LC_9_15_6  (
            .in0(N__41029),
            .in1(N__41080),
            .in2(N__41110),
            .in3(N__42555),
            .lcout(\quad_counter0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1515_LC_9_16_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1515_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1515_LC_9_16_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \c0.i1_4_lut_adj_1515_LC_9_16_0  (
            .in0(N__48372),
            .in1(N__92680),
            .in2(N__48755),
            .in3(N__38853),
            .lcout(\c0.n2107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i7_3_lut_LC_9_16_2 .C_ON=1'b0;
    defparam \quad_counter0.i7_3_lut_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i7_3_lut_LC_9_16_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter0.i7_3_lut_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__41197),
            .in2(N__41260),
            .in3(N__41167),
            .lcout(\quad_counter0.n20_adj_4351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_LC_9_16_4 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_LC_9_16_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i9_4_lut_LC_9_16_4  (
            .in0(N__41335),
            .in1(N__41281),
            .in2(N__41314),
            .in3(N__41224),
            .lcout(),
            .ltout(\quad_counter0.n22_adj_4350_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1165_LC_9_16_5 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1165_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1165_LC_9_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1165_LC_9_16_5  (
            .in0(N__40951),
            .in1(N__41002),
            .in2(N__38835),
            .in3(N__38832),
            .lcout(\quad_counter0.n24_adj_4352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23145_2_lut_LC_9_16_6 .C_ON=1'b0;
    defparam \c0.i23145_2_lut_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i23145_2_lut_LC_9_16_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.i23145_2_lut_LC_9_16_6  (
            .in0(N__51381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92618),
            .lcout(\c0.n3844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1519_LC_9_16_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1519_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1519_LC_9_16_7 .LUT_INIT=16'b1111111110001100;
    LogicCell40 \c0.i1_4_lut_adj_1519_LC_9_16_7  (
            .in0(N__38973),
            .in1(N__49008),
            .in2(N__42885),
            .in3(N__38820),
            .lcout(\c0.n4_adj_4615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_9_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_9_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i2_LC_9_17_0 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_9_17_0  (
            .in0(N__51685),
            .in1(N__38787),
            .in2(N__39057),
            .in3(N__48191),
            .lcout(\c0.FRAME_MATCHER_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97669),
            .ce(),
            .sr(N__96949));
    defparam \c0.i2_4_lut_adj_1525_LC_9_17_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1525_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1525_LC_9_17_1 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \c0.i2_4_lut_adj_1525_LC_9_17_1  (
            .in0(N__48624),
            .in1(N__51684),
            .in2(N__38796),
            .in3(N__49007),
            .lcout(\c0.n6_adj_4618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_9_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_9_17_2 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_9_17_2  (
            .in0(N__48492),
            .in1(N__48443),
            .in2(N__39027),
            .in3(N__39047),
            .lcout(),
            .ltout(\c0.n33215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1524_LC_9_17_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1524_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1524_LC_9_17_3 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \c0.i1_4_lut_adj_1524_LC_9_17_3  (
            .in0(N__39000),
            .in1(N__46241),
            .in2(N__39060),
            .in3(N__38993),
            .lcout(\c0.n6_adj_4616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6290_2_lut_3_lut_4_lut_LC_9_17_5 .C_ON=1'b0;
    defparam \c0.i6290_2_lut_3_lut_4_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6290_2_lut_3_lut_4_lut_LC_9_17_5 .LUT_INIT=16'b1110111000001110;
    LogicCell40 \c0.i6290_2_lut_3_lut_4_lut_LC_9_17_5  (
            .in0(N__39048),
            .in1(N__39022),
            .in2(N__55239),
            .in3(N__92622),
            .lcout(\c0.n10800 ),
            .ltout(\c0.n10800_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_9_17_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_9_17_6 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i1_LC_9_17_6 .LUT_INIT=16'b1111111110001010;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_9_17_6  (
            .in0(N__38994),
            .in1(N__38972),
            .in2(N__38946),
            .in3(N__38943),
            .lcout(\c0.FRAME_MATCHER_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97669),
            .ce(),
            .sr(N__96949));
    defparam \c0.i1_2_lut_4_lut_adj_1371_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1371_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1371_LC_9_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1371_LC_9_18_0  (
            .in0(N__52060),
            .in1(N__48787),
            .in2(N__48853),
            .in3(N__39215),
            .lcout(\c0.n33454 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_9_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_9_18_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i19_LC_9_18_2  (
            .in0(N__80268),
            .in1(N__83970),
            .in2(N__48800),
            .in3(N__80554),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1474_LC_9_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1474_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1474_LC_9_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1474_LC_9_18_4  (
            .in0(N__38924),
            .in1(N__61209),
            .in2(N__38889),
            .in3(N__43316),
            .lcout(\c0.n6_adj_4564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1966_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1966_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1966_LC_9_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1966_LC_9_18_5  (
            .in0(N__39112),
            .in1(N__52059),
            .in2(_gnd_net_),
            .in3(N__52149),
            .lcout(\c0.n18671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_9_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_9_18_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i3_LC_9_18_6  (
            .in0(N__81246),
            .in1(N__80553),
            .in2(N__52162),
            .in3(N__83971),
            .lcout(\c0.data_in_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_9_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_9_18_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i20_LC_9_18_7  (
            .in0(N__83969),
            .in1(N__78909),
            .in2(N__39117),
            .in3(N__80269),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30381_4_lut_LC_9_19_0 .C_ON=1'b0;
    defparam \c0.i30381_4_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i30381_4_lut_LC_9_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i30381_4_lut_LC_9_19_0  (
            .in0(N__41357),
            .in1(N__39116),
            .in2(N__48861),
            .in3(N__52154),
            .lcout(\c0.n35808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1613_LC_9_19_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1613_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1613_LC_9_19_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.i2_3_lut_adj_1613_LC_9_19_1  (
            .in0(N__46440),
            .in1(N__51931),
            .in2(_gnd_net_),
            .in3(N__51838),
            .lcout(\c0.n19388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_2000_LC_9_19_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_2000_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_2000_LC_9_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_2000_LC_9_19_2  (
            .in0(N__43351),
            .in1(N__39089),
            .in2(_gnd_net_),
            .in3(N__41505),
            .lcout(\c0.data_out_frame_0__7__N_2747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2773_2_lut_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.i2773_2_lut_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2773_2_lut_LC_9_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2773_2_lut_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__46646),
            .in2(_gnd_net_),
            .in3(N__46941),
            .lcout(),
            .ltout(\c0.n5452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1803_LC_9_19_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1803_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1803_LC_9_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1803_LC_9_19_5  (
            .in0(N__39148),
            .in1(N__39099),
            .in2(N__39093),
            .in3(N__43665),
            .lcout(\c0.n33800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1339_LC_9_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1339_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1339_LC_9_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1339_LC_9_19_6  (
            .in0(N__41356),
            .in1(N__52153),
            .in2(_gnd_net_),
            .in3(N__52120),
            .lcout(\c0.n19030 ),
            .ltout(\c0.n19030_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1412_LC_9_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1412_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1412_LC_9_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1412_LC_9_19_7  (
            .in0(N__39088),
            .in1(N__43350),
            .in2(N__39063),
            .in3(N__52199),
            .lcout(\c0.n33476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1881_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1881_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1881_LC_9_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1881_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__41758),
            .in2(_gnd_net_),
            .in3(N__48897),
            .lcout(\c0.n33695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i91_LC_9_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i91_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i91_LC_9_20_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i91_LC_9_20_2  (
            .in0(N__80547),
            .in1(N__58436),
            .in2(N__39156),
            .in3(N__78286),
            .lcout(\c0.data_in_frame_11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97723),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i40_LC_9_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i40_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i40_LC_9_20_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i40_LC_9_20_5  (
            .in0(N__73926),
            .in1(N__83973),
            .in2(N__41465),
            .in3(N__80053),
            .lcout(\c0.data_in_frame_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97723),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_9_20_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_9_20_6  (
            .in0(N__83972),
            .in1(N__78285),
            .in2(N__41418),
            .in3(N__75324),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97723),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_103_i4_2_lut_LC_9_20_7 .C_ON=1'b0;
    defparam \c0.rx.equal_103_i4_2_lut_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_103_i4_2_lut_LC_9_20_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.equal_103_i4_2_lut_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__55447),
            .in2(_gnd_net_),
            .in3(N__55557),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i89_LC_9_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i89_LC_9_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i89_LC_9_21_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i89_LC_9_21_0  (
            .in0(N__80910),
            .in1(N__58416),
            .in2(N__78320),
            .in3(N__39451),
            .lcout(\c0.data_in_frame_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_1829_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_1829_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_1829_LC_9_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_1829_LC_9_21_1  (
            .in0(N__49609),
            .in1(N__47103),
            .in2(N__39155),
            .in3(N__39342),
            .lcout(\c0.n47_adj_4729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i69_LC_9_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i69_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i69_LC_9_21_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i69_LC_9_21_2  (
            .in0(N__84116),
            .in1(N__58415),
            .in2(N__81260),
            .in3(N__41762),
            .lcout(\c0.data_in_frame_8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i71_LC_9_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i71_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i71_LC_9_21_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i71_LC_9_21_3  (
            .in0(N__58413),
            .in1(N__81240),
            .in2(N__41791),
            .in3(N__73616),
            .lcout(\c0.data_in_frame_8_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97739),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1855_LC_9_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1855_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1855_LC_9_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1855_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__41900),
            .in2(_gnd_net_),
            .in3(N__61176),
            .lcout(\c0.n33404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1490_LC_9_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1490_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1490_LC_9_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1490_LC_9_21_5  (
            .in0(N__41781),
            .in1(N__48965),
            .in2(N__39455),
            .in3(N__46413),
            .lcout(\c0.n33714 ),
            .ltout(\c0.n33714_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1828_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1828_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1828_LC_9_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1828_LC_9_21_6  (
            .in0(N__43761),
            .in1(N__39129),
            .in2(N__39120),
            .in3(N__52200),
            .lcout(\c0.n46_adj_4728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i81_LC_9_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i81_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i81_LC_9_21_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i81_LC_9_21_7  (
            .in0(N__58414),
            .in1(N__80911),
            .in2(N__49616),
            .in3(N__80331),
            .lcout(\c0.data_in_frame_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97739),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_9_22_1 .C_ON=1'b0;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.A_filtered_I_0_2_lut_LC_9_22_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.A_filtered_I_0_2_lut_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__39402),
            .in2(_gnd_net_),
            .in3(N__39289),
            .lcout(\quad_counter0.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1882_LC_9_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1882_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1882_LC_9_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1882_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__44173),
            .in2(_gnd_net_),
            .in3(N__50216),
            .lcout(\c0.n33883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1084_1_lut_2_lut_LC_9_22_3 .C_ON=1'b0;
    defparam \quad_counter0.i1084_1_lut_2_lut_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1084_1_lut_2_lut_LC_9_22_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter0.i1084_1_lut_2_lut_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__39401),
            .in2(_gnd_net_),
            .in3(N__39288),
            .lcout(\quad_counter0.n2300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1983_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1983_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1983_LC_9_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1983_LC_9_22_4  (
            .in0(N__52302),
            .in1(N__39245),
            .in2(N__48927),
            .in3(N__77202),
            .lcout(),
            .ltout(\c0.n10_adj_4769_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1984_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1984_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1984_LC_9_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1984_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__39182),
            .in2(N__39219),
            .in3(N__39216),
            .lcout(\c0.n18330 ),
            .ltout(\c0.n18330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_9_22_6 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_9_22_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i5_2_lut_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39186),
            .in3(N__43719),
            .lcout(\c0.n16_adj_4726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_9_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_9_22_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i54_LC_9_22_7  (
            .in0(N__83867),
            .in1(N__75089),
            .in2(N__89819),
            .in3(N__39183),
            .lcout(\c0.data_in_frame_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97758),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1465_LC_9_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1465_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1465_LC_9_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1465_LC_9_23_0  (
            .in0(N__48974),
            .in1(N__41792),
            .in2(N__41630),
            .in3(N__46414),
            .lcout(\c0.n18364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1436_LC_9_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1436_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1436_LC_9_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1436_LC_9_23_1  (
            .in0(N__42037),
            .in1(N__39328),
            .in2(_gnd_net_),
            .in3(N__52355),
            .lcout(\c0.n33997 ),
            .ltout(\c0.n33997_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1792_LC_9_23_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1792_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1792_LC_9_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1792_LC_9_23_2  (
            .in0(N__39435),
            .in1(N__41823),
            .in2(N__39333),
            .in3(N__39261),
            .lcout(\c0.n33371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i70_LC_9_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i70_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i70_LC_9_23_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i70_LC_9_23_3  (
            .in0(N__75088),
            .in1(N__81247),
            .in2(N__43721),
            .in3(N__58406),
            .lcout(\c0.data_in_frame_8_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97772),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1826_LC_9_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1826_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1826_LC_9_23_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1826_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__42038),
            .in2(_gnd_net_),
            .in3(N__39330),
            .lcout(\c0.n33923 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1404_LC_9_23_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1404_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1404_LC_9_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1404_LC_9_23_5  (
            .in0(N__39329),
            .in1(N__48973),
            .in2(N__43720),
            .in3(N__48905),
            .lcout(\c0.n19190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1898_LC_9_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1898_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1898_LC_9_23_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1898_LC_9_23_6  (
            .in0(N__48975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43712),
            .lcout(\c0.n33705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.A_delayed_76_LC_9_24_0 .C_ON=1'b0;
    defparam \quad_counter0.A_delayed_76_LC_9_24_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.A_delayed_76_LC_9_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.A_delayed_76_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39299),
            .lcout(\quad_counter0.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97787),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_adj_1230_LC_9_24_1 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_adj_1230_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_adj_1230_LC_9_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter0.i3_4_lut_adj_1230_LC_9_24_1  (
            .in0(N__39400),
            .in1(N__39306),
            .in2(N__39300),
            .in3(N__39428),
            .lcout(count_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1455_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1455_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1455_LC_9_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1455_LC_9_24_2  (
            .in0(N__39361),
            .in1(N__39260),
            .in2(N__50127),
            .in3(N__47141),
            .lcout(\c0.n18147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1791_LC_9_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1791_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1791_LC_9_24_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1791_LC_9_24_3  (
            .in0(N__39456),
            .in1(N__44106),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n6_adj_4713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.B_delayed_77_LC_9_24_4 .C_ON=1'b0;
    defparam \quad_counter0.B_delayed_77_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.B_delayed_77_LC_9_24_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.B_delayed_77_LC_9_24_4  (
            .in0(N__39429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1883_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1883_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1883_LC_9_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1883_LC_9_24_5  (
            .in0(N__39384),
            .in1(N__41728),
            .in2(_gnd_net_),
            .in3(N__41652),
            .lcout(\c0.n5896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1425_LC_9_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1425_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1425_LC_9_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1425_LC_9_24_6  (
            .in0(N__39362),
            .in1(N__52359),
            .in2(N__50128),
            .in3(N__47142),
            .lcout(\c0.n33982 ),
            .ltout(\c0.n33982_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1794_LC_9_24_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1794_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1794_LC_9_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1794_LC_9_24_7  (
            .in0(N__39375),
            .in1(N__44223),
            .in2(N__39366),
            .in3(N__41729),
            .lcout(\c0.n18861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i95_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i95_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i95_LC_9_25_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i95_LC_9_25_0  (
            .in0(N__73637),
            .in1(N__58404),
            .in2(N__41952),
            .in3(N__78210),
            .lcout(\c0.data_in_frame_11_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i87_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i87_LC_9_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i87_LC_9_25_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i87_LC_9_25_1  (
            .in0(N__58402),
            .in1(N__80411),
            .in2(N__42039),
            .in3(N__73639),
            .lcout(\c0.data_in_frame_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i86_LC_9_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i86_LC_9_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i86_LC_9_25_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i86_LC_9_25_4  (
            .in0(N__80410),
            .in1(N__58403),
            .in2(N__39363),
            .in3(N__75072),
            .lcout(\c0.data_in_frame_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i119_LC_9_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i119_LC_9_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i119_LC_9_25_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i119_LC_9_25_5  (
            .in0(N__58401),
            .in1(N__73638),
            .in2(N__44344),
            .in3(N__89784),
            .lcout(\c0.data_in_frame_14_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3317_2_lut_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.i3317_2_lut_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3317_2_lut_LC_9_25_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3317_2_lut_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__44335),
            .in2(_gnd_net_),
            .in3(N__44456),
            .lcout(\c0.n5996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1894_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1894_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1894_LC_9_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1894_LC_9_26_6  (
            .in0(N__53225),
            .in1(N__52832),
            .in2(_gnd_net_),
            .in3(N__52761),
            .lcout(\c0.n18431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadA_I_0_85_2_lut_LC_10_5_0 .C_ON=1'b0;
    defparam \quad_counter1.quadA_I_0_85_2_lut_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadA_I_0_85_2_lut_LC_10_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter1.quadA_I_0_85_2_lut_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__44589),
            .in2(_gnd_net_),
            .in3(N__44527),
            .lcout(a_delay_counter_15__N_4220_adj_4817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_delayed_71_LC_10_5_4 .C_ON=1'b0;
    defparam \quad_counter1.quadB_delayed_71_LC_10_5_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadB_delayed_71_LC_10_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter1.quadB_delayed_71_LC_10_5_4  (
            .in0(N__42144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadB_delayed_adj_4813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97544),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.a_delay_counter__i0_LC_10_7_1 .C_ON=1'b0;
    defparam \quad_counter1.a_delay_counter__i0_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.a_delay_counter__i0_LC_10_7_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \quad_counter1.a_delay_counter__i0_LC_10_7_1  (
            .in0(N__39661),
            .in1(N__39642),
            .in2(N__39573),
            .in3(N__39766),
            .lcout(a_delay_counter_0_adj_4811),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97552),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1263_LC_10_7_2 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1263_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1263_LC_10_7_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1263_LC_10_7_2  (
            .in0(N__39635),
            .in1(N__39623),
            .in2(N__39612),
            .in3(N__39596),
            .lcout(\quad_counter1.n28_adj_4440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1266_LC_10_7_5 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1266_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1266_LC_10_7_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1266_LC_10_7_5  (
            .in0(N__39584),
            .in1(N__39565),
            .in2(N__39549),
            .in3(N__39533),
            .lcout(\quad_counter1.n25_adj_4443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1265_LC_10_8_0 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1265_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1265_LC_10_8_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1265_LC_10_8_0  (
            .in0(N__39521),
            .in1(N__39509),
            .in2(N__39498),
            .in3(N__39482),
            .lcout(),
            .ltout(\quad_counter1.n27_adj_4442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_adj_1267_LC_10_8_1 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_adj_1267_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_adj_1267_LC_10_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_adj_1267_LC_10_8_1  (
            .in0(N__39471),
            .in1(N__39696),
            .in2(N__39465),
            .in3(N__39462),
            .lcout(n17985),
            .ltout(n17985_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_10_8_2.C_ON=1'b0;
    defparam i1_3_lut_LC_10_8_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_10_8_2.LUT_INIT=16'b1111010111111010;
    LogicCell40 i1_3_lut_LC_10_8_2 (
            .in0(N__44534),
            .in1(_gnd_net_),
            .in2(N__39771),
            .in3(N__44601),
            .lcout(n19433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1264_LC_10_8_6 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1264_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1264_LC_10_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1264_LC_10_8_6  (
            .in0(N__39749),
            .in1(N__39737),
            .in2(N__39726),
            .in3(N__39707),
            .lcout(\quad_counter1.n26_adj_4441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_2_lut_LC_10_9_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_2_lut_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_2_lut_LC_10_9_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2219_2_lut_LC_10_9_0  (
            .in0(N__59883),
            .in1(N__59882),
            .in2(N__39859),
            .in3(N__39690),
            .lcout(\quad_counter0.n3319 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\quad_counter0.n30384 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_3_lut_LC_10_9_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_3_lut_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_3_lut_LC_10_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_3_lut_LC_10_9_1  (
            .in0(N__42393),
            .in1(N__42389),
            .in2(N__39974),
            .in3(N__39687),
            .lcout(\quad_counter0.n3318 ),
            .ltout(),
            .carryin(\quad_counter0.n30384 ),
            .carryout(\quad_counter0.n30385 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_4_lut_LC_10_9_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_4_lut_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_4_lut_LC_10_9_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2219_4_lut_LC_10_9_2  (
            .in0(N__42365),
            .in1(N__42366),
            .in2(N__39860),
            .in3(N__39684),
            .lcout(\quad_counter0.n3317 ),
            .ltout(),
            .carryin(\quad_counter0.n30385 ),
            .carryout(\quad_counter0.n30386 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_5_lut_LC_10_9_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_5_lut_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_5_lut_LC_10_9_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2219_5_lut_LC_10_9_3  (
            .in0(N__42342),
            .in1(N__42341),
            .in2(N__39863),
            .in3(N__39681),
            .lcout(\quad_counter0.n3316 ),
            .ltout(),
            .carryin(\quad_counter0.n30386 ),
            .carryout(\quad_counter0.n30387 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_6_lut_LC_10_9_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_6_lut_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_6_lut_LC_10_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2219_6_lut_LC_10_9_4  (
            .in0(N__40256),
            .in1(N__40255),
            .in2(N__39861),
            .in3(N__39678),
            .lcout(\quad_counter0.n3315 ),
            .ltout(),
            .carryin(\quad_counter0.n30387 ),
            .carryout(\quad_counter0.n30388 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_7_lut_LC_10_9_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_7_lut_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_7_lut_LC_10_9_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2219_7_lut_LC_10_9_5  (
            .in0(N__40203),
            .in1(N__40202),
            .in2(N__39864),
            .in3(N__39675),
            .lcout(\quad_counter0.n3314 ),
            .ltout(),
            .carryin(\quad_counter0.n30388 ),
            .carryout(\quad_counter0.n30389 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_8_lut_LC_10_9_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_8_lut_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_8_lut_LC_10_9_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2219_8_lut_LC_10_9_6  (
            .in0(N__42315),
            .in1(N__42314),
            .in2(N__39862),
            .in3(N__39672),
            .lcout(\quad_counter0.n3313 ),
            .ltout(),
            .carryin(\quad_counter0.n30389 ),
            .carryout(\quad_counter0.n30390 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_9_lut_LC_10_9_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_9_lut_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_9_lut_LC_10_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_9_lut_LC_10_9_7  (
            .in0(N__40113),
            .in1(N__40112),
            .in2(N__39975),
            .in3(N__39798),
            .lcout(\quad_counter0.n3312 ),
            .ltout(),
            .carryin(\quad_counter0.n30390 ),
            .carryout(\quad_counter0.n30391 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_10_lut_LC_10_10_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_10_lut_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_10_lut_LC_10_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_10_lut_LC_10_10_0  (
            .in0(N__40065),
            .in1(N__40064),
            .in2(N__39964),
            .in3(N__39795),
            .lcout(\quad_counter0.n3311 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\quad_counter0.n30392 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_11_lut_LC_10_10_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_11_lut_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_11_lut_LC_10_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_11_lut_LC_10_10_1  (
            .in0(N__40020),
            .in1(N__40019),
            .in2(N__39968),
            .in3(N__39792),
            .lcout(\quad_counter0.n3310 ),
            .ltout(),
            .carryin(\quad_counter0.n30392 ),
            .carryout(\quad_counter0.n30393 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_12_lut_LC_10_10_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_12_lut_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_12_lut_LC_10_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_12_lut_LC_10_10_2  (
            .in0(N__40647),
            .in1(N__40646),
            .in2(N__39965),
            .in3(N__39789),
            .lcout(\quad_counter0.n3309 ),
            .ltout(),
            .carryin(\quad_counter0.n30393 ),
            .carryout(\quad_counter0.n30394 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_13_lut_LC_10_10_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_13_lut_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_13_lut_LC_10_10_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_13_lut_LC_10_10_3  (
            .in0(N__40599),
            .in1(N__40598),
            .in2(N__39969),
            .in3(N__39786),
            .lcout(\quad_counter0.n3308 ),
            .ltout(),
            .carryin(\quad_counter0.n30394 ),
            .carryout(\quad_counter0.n30395 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_14_lut_LC_10_10_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_14_lut_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_14_lut_LC_10_10_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_14_lut_LC_10_10_4  (
            .in0(N__40554),
            .in1(N__40553),
            .in2(N__39966),
            .in3(N__39783),
            .lcout(\quad_counter0.n3307 ),
            .ltout(),
            .carryin(\quad_counter0.n30395 ),
            .carryout(\quad_counter0.n30396 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_15_lut_LC_10_10_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_15_lut_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_15_lut_LC_10_10_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_15_lut_LC_10_10_5  (
            .in0(N__40508),
            .in1(N__40507),
            .in2(N__39970),
            .in3(N__39780),
            .lcout(\quad_counter0.n3306 ),
            .ltout(),
            .carryin(\quad_counter0.n30396 ),
            .carryout(\quad_counter0.n30397 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_16_lut_LC_10_10_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_16_lut_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_16_lut_LC_10_10_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_16_lut_LC_10_10_6  (
            .in0(N__40460),
            .in1(N__40459),
            .in2(N__39967),
            .in3(N__39777),
            .lcout(\quad_counter0.n3305 ),
            .ltout(),
            .carryin(\quad_counter0.n30397 ),
            .carryout(\quad_counter0.n30398 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_17_lut_LC_10_10_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_17_lut_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_17_lut_LC_10_10_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_17_lut_LC_10_10_7  (
            .in0(N__40413),
            .in1(N__40412),
            .in2(N__39971),
            .in3(N__39774),
            .lcout(\quad_counter0.n3304 ),
            .ltout(),
            .carryin(\quad_counter0.n30398 ),
            .carryout(\quad_counter0.n30399 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_18_lut_LC_10_11_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_18_lut_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_18_lut_LC_10_11_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_18_lut_LC_10_11_0  (
            .in0(N__40365),
            .in1(N__40364),
            .in2(N__39955),
            .in3(N__39990),
            .lcout(\quad_counter0.n3303 ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\quad_counter0.n30400 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_19_lut_LC_10_11_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_19_lut_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_19_lut_LC_10_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_19_lut_LC_10_11_1  (
            .in0(N__40322),
            .in1(N__40323),
            .in2(N__39972),
            .in3(N__39987),
            .lcout(\quad_counter0.n3302 ),
            .ltout(),
            .carryin(\quad_counter0.n30400 ),
            .carryout(\quad_counter0.n30401 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_20_lut_LC_10_11_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_20_lut_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_20_lut_LC_10_11_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_20_lut_LC_10_11_2  (
            .in0(N__40916),
            .in1(N__40915),
            .in2(N__39956),
            .in3(N__39984),
            .lcout(\quad_counter0.n3301 ),
            .ltout(),
            .carryin(\quad_counter0.n30401 ),
            .carryout(\quad_counter0.n30402 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_21_lut_LC_10_11_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2219_21_lut_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_21_lut_LC_10_11_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_21_lut_LC_10_11_3  (
            .in0(N__40866),
            .in1(N__40865),
            .in2(N__39973),
            .in3(N__39981),
            .lcout(\quad_counter0.n3300 ),
            .ltout(),
            .carryin(\quad_counter0.n30402 ),
            .carryout(\quad_counter0.n30403 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2219_22_lut_LC_10_11_4 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_2219_22_lut_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2219_22_lut_LC_10_11_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2219_22_lut_LC_10_11_4  (
            .in0(N__40711),
            .in1(N__40712),
            .in2(N__39957),
            .in3(N__39978),
            .lcout(\quad_counter0.n3299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30714_1_lut_LC_10_11_5 .C_ON=1'b0;
    defparam \quad_counter0.i30714_1_lut_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30714_1_lut_LC_10_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30714_1_lut_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39910),
            .lcout(\quad_counter0.n36141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1172_LC_10_11_6 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1172_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1172_LC_10_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1172_LC_10_11_6  (
            .in0(N__40552),
            .in1(N__40363),
            .in2(N__40509),
            .in3(N__40321),
            .lcout(\quad_counter0.n26_adj_4358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_2_lut_LC_10_11_7 .C_ON=1'b0;
    defparam \quad_counter0.i1_2_lut_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_2_lut_LC_10_11_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i1_2_lut_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40063),
            .in3(N__40864),
            .lcout(\quad_counter0.n16_adj_4359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_2_lut_LC_10_12_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_2_lut_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_2_lut_LC_10_12_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2152_2_lut_LC_10_12_0  (
            .in0(N__59853),
            .in1(N__59852),
            .in2(N__40150),
            .in3(N__39801),
            .lcout(\quad_counter0.n3219 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\quad_counter0.n30365 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_3_lut_LC_10_12_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_3_lut_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_3_lut_LC_10_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_3_lut_LC_10_12_1  (
            .in0(N__40302),
            .in1(N__40301),
            .in2(N__40799),
            .in3(N__40284),
            .lcout(\quad_counter0.n3218 ),
            .ltout(),
            .carryin(\quad_counter0.n30365 ),
            .carryout(\quad_counter0.n30366 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_4_lut_LC_10_12_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_4_lut_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_4_lut_LC_10_12_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2152_4_lut_LC_10_12_2  (
            .in0(N__40280),
            .in1(N__40279),
            .in2(N__40151),
            .in3(N__40260),
            .lcout(\quad_counter0.n3217 ),
            .ltout(),
            .carryin(\quad_counter0.n30366 ),
            .carryout(\quad_counter0.n30367 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_5_lut_LC_10_12_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_5_lut_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_5_lut_LC_10_12_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2152_5_lut_LC_10_12_3  (
            .in0(N__70697),
            .in1(N__70696),
            .in2(N__40154),
            .in3(N__40227),
            .lcout(\quad_counter0.n3216 ),
            .ltout(),
            .carryin(\quad_counter0.n30367 ),
            .carryout(\quad_counter0.n30368 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_6_lut_LC_10_12_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_6_lut_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_6_lut_LC_10_12_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2152_6_lut_LC_10_12_4  (
            .in0(N__40224),
            .in1(N__40223),
            .in2(N__40152),
            .in3(N__40179),
            .lcout(\quad_counter0.n3215 ),
            .ltout(),
            .carryin(\quad_counter0.n30368 ),
            .carryout(\quad_counter0.n30369 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_7_lut_LC_10_12_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_7_lut_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_7_lut_LC_10_12_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2152_7_lut_LC_10_12_5  (
            .in0(N__40176),
            .in1(N__40175),
            .in2(N__40155),
            .in3(N__40158),
            .lcout(\quad_counter0.n3214 ),
            .ltout(),
            .carryin(\quad_counter0.n30369 ),
            .carryout(\quad_counter0.n30370 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_8_lut_LC_10_12_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_8_lut_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_8_lut_LC_10_12_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2152_8_lut_LC_10_12_6  (
            .in0(N__70667),
            .in1(N__70666),
            .in2(N__40153),
            .in3(N__40086),
            .lcout(\quad_counter0.n3213 ),
            .ltout(),
            .carryin(\quad_counter0.n30370 ),
            .carryout(\quad_counter0.n30371 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_9_lut_LC_10_12_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_9_lut_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_9_lut_LC_10_12_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_9_lut_LC_10_12_7  (
            .in0(N__40083),
            .in1(N__40082),
            .in2(N__40800),
            .in3(N__40041),
            .lcout(\quad_counter0.n3212 ),
            .ltout(),
            .carryin(\quad_counter0.n30371 ),
            .carryout(\quad_counter0.n30372 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_10_lut_LC_10_13_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_10_lut_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_10_lut_LC_10_13_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_10_lut_LC_10_13_0  (
            .in0(N__40038),
            .in1(N__40037),
            .in2(N__40801),
            .in3(N__39993),
            .lcout(\quad_counter0.n3211 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\quad_counter0.n30373 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_11_lut_LC_10_13_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_11_lut_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_11_lut_LC_10_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_11_lut_LC_10_13_1  (
            .in0(N__40667),
            .in1(N__40666),
            .in2(N__40805),
            .in3(N__40623),
            .lcout(\quad_counter0.n3210 ),
            .ltout(),
            .carryin(\quad_counter0.n30373 ),
            .carryout(\quad_counter0.n30374 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_12_lut_LC_10_13_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_12_lut_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_12_lut_LC_10_13_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_12_lut_LC_10_13_2  (
            .in0(N__40619),
            .in1(N__40618),
            .in2(N__40802),
            .in3(N__40578),
            .lcout(\quad_counter0.n3209 ),
            .ltout(),
            .carryin(\quad_counter0.n30374 ),
            .carryout(\quad_counter0.n30375 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_13_lut_LC_10_13_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_13_lut_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_13_lut_LC_10_13_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_13_lut_LC_10_13_3  (
            .in0(N__40574),
            .in1(N__40573),
            .in2(N__40806),
            .in3(N__40530),
            .lcout(\quad_counter0.n3208 ),
            .ltout(),
            .carryin(\quad_counter0.n30375 ),
            .carryout(\quad_counter0.n30376 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_14_lut_LC_10_13_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_14_lut_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_14_lut_LC_10_13_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_14_lut_LC_10_13_4  (
            .in0(N__40527),
            .in1(N__40526),
            .in2(N__40803),
            .in3(N__40485),
            .lcout(\quad_counter0.n3207 ),
            .ltout(),
            .carryin(\quad_counter0.n30376 ),
            .carryout(\quad_counter0.n30377 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_15_lut_LC_10_13_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_15_lut_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_15_lut_LC_10_13_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_15_lut_LC_10_13_5  (
            .in0(N__40481),
            .in1(N__40480),
            .in2(N__40807),
            .in3(N__40437),
            .lcout(\quad_counter0.n3206 ),
            .ltout(),
            .carryin(\quad_counter0.n30377 ),
            .carryout(\quad_counter0.n30378 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_16_lut_LC_10_13_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_16_lut_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_16_lut_LC_10_13_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_16_lut_LC_10_13_6  (
            .in0(N__40434),
            .in1(N__40433),
            .in2(N__40804),
            .in3(N__40389),
            .lcout(\quad_counter0.n3205 ),
            .ltout(),
            .carryin(\quad_counter0.n30378 ),
            .carryout(\quad_counter0.n30379 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_17_lut_LC_10_13_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_17_lut_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_17_lut_LC_10_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_17_lut_LC_10_13_7  (
            .in0(N__40385),
            .in1(N__40384),
            .in2(N__40808),
            .in3(N__40347),
            .lcout(\quad_counter0.n3204 ),
            .ltout(),
            .carryin(\quad_counter0.n30379 ),
            .carryout(\quad_counter0.n30380 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_18_lut_LC_10_14_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_18_lut_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_18_lut_LC_10_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_18_lut_LC_10_14_0  (
            .in0(N__40343),
            .in1(N__40342),
            .in2(N__40821),
            .in3(N__40305),
            .lcout(\quad_counter0.n3203 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\quad_counter0.n30381 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_19_lut_LC_10_14_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_19_lut_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_19_lut_LC_10_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_19_lut_LC_10_14_1  (
            .in0(N__40935),
            .in1(N__40934),
            .in2(N__40823),
            .in3(N__40890),
            .lcout(\quad_counter0.n3202 ),
            .ltout(),
            .carryin(\quad_counter0.n30381 ),
            .carryout(\quad_counter0.n30382 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_20_lut_LC_10_14_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2152_20_lut_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_20_lut_LC_10_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_20_lut_LC_10_14_2  (
            .in0(N__40886),
            .in1(N__40885),
            .in2(N__40822),
            .in3(N__40848),
            .lcout(\quad_counter0.n3201 ),
            .ltout(),
            .carryin(\quad_counter0.n30382 ),
            .carryout(\quad_counter0.n30383 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2152_21_lut_LC_10_14_3 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_2152_21_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2152_21_lut_LC_10_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2152_21_lut_LC_10_14_3  (
            .in0(N__40843),
            .in1(N__40844),
            .in2(N__40824),
            .in3(N__40716),
            .lcout(\quad_counter0.n3200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1342_LC_10_14_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1342_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1342_LC_10_14_4 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1342_LC_10_14_4  (
            .in0(N__49122),
            .in1(N__51821),
            .in2(N__49184),
            .in3(N__49263),
            .lcout(\c0.n111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1566_LC_10_14_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1566_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1566_LC_10_14_6 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \c0.i1_4_lut_adj_1566_LC_10_14_6  (
            .in0(N__48538),
            .in1(N__48312),
            .in2(N__48491),
            .in3(N__40689),
            .lcout(\c0.n10_adj_4629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1560_LC_10_14_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1560_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1560_LC_10_14_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1560_LC_10_14_7  (
            .in0(N__49264),
            .in1(N__51437),
            .in2(N__49120),
            .in3(N__49180),
            .lcout(\c0.n29678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_2_lut_LC_10_15_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_2_lut_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_2_lut_LC_10_15_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2018_2_lut_LC_10_15_0  (
            .in0(N__59768),
            .in1(N__59767),
            .in2(N__43087),
            .in3(N__40677),
            .lcout(\quad_counter0.n3019 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\quad_counter0.n30330 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_3_lut_LC_10_15_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_3_lut_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_3_lut_LC_10_15_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_3_lut_LC_10_15_1  (
            .in0(N__43112),
            .in1(N__43111),
            .in2(N__43595),
            .in3(N__40674),
            .lcout(\quad_counter0.n3018 ),
            .ltout(),
            .carryin(\quad_counter0.n30330 ),
            .carryout(\quad_counter0.n30331 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_4_lut_LC_10_15_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_4_lut_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_4_lut_LC_10_15_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2018_4_lut_LC_10_15_2  (
            .in0(N__43478),
            .in1(N__43477),
            .in2(N__43088),
            .in3(N__40671),
            .lcout(\quad_counter0.n3017 ),
            .ltout(),
            .carryin(\quad_counter0.n30331 ),
            .carryout(\quad_counter0.n30332 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_5_lut_LC_10_15_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_5_lut_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_5_lut_LC_10_15_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2018_5_lut_LC_10_15_3  (
            .in0(N__43499),
            .in1(N__43498),
            .in2(N__43091),
            .in3(N__41091),
            .lcout(\quad_counter0.n3016 ),
            .ltout(),
            .carryin(\quad_counter0.n30332 ),
            .carryout(\quad_counter0.n30333 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_6_lut_LC_10_15_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_6_lut_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_6_lut_LC_10_15_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2018_6_lut_LC_10_15_4  (
            .in0(N__43427),
            .in1(N__43426),
            .in2(N__43089),
            .in3(N__41067),
            .lcout(\quad_counter0.n3015 ),
            .ltout(),
            .carryin(\quad_counter0.n30333 ),
            .carryout(\quad_counter0.n30334 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_7_lut_LC_10_15_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_7_lut_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_7_lut_LC_10_15_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2018_7_lut_LC_10_15_5  (
            .in0(N__43405),
            .in1(N__43406),
            .in2(N__43092),
            .in3(N__41064),
            .lcout(\quad_counter0.n3014 ),
            .ltout(),
            .carryin(\quad_counter0.n30334 ),
            .carryout(\quad_counter0.n30335 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_8_lut_LC_10_15_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_8_lut_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_8_lut_LC_10_15_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2018_8_lut_LC_10_15_6  (
            .in0(N__43454),
            .in1(N__43453),
            .in2(N__43090),
            .in3(N__41034),
            .lcout(\quad_counter0.n3013 ),
            .ltout(),
            .carryin(\quad_counter0.n30335 ),
            .carryout(\quad_counter0.n30336 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_9_lut_LC_10_15_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_9_lut_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_9_lut_LC_10_15_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_9_lut_LC_10_15_7  (
            .in0(N__43172),
            .in1(N__43171),
            .in2(N__43596),
            .in3(N__41013),
            .lcout(\quad_counter0.n3012 ),
            .ltout(),
            .carryin(\quad_counter0.n30336 ),
            .carryout(\quad_counter0.n30337 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_10_lut_LC_10_16_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_10_lut_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_10_lut_LC_10_16_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_10_lut_LC_10_16_0  (
            .in0(N__43050),
            .in1(N__43046),
            .in2(N__43585),
            .in3(N__40989),
            .lcout(\quad_counter0.n3011 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\quad_counter0.n30338 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_11_lut_LC_10_16_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_11_lut_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_11_lut_LC_10_16_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_11_lut_LC_10_16_1  (
            .in0(N__43625),
            .in1(N__43624),
            .in2(N__43589),
            .in3(N__40962),
            .lcout(\quad_counter0.n3010 ),
            .ltout(),
            .carryin(\quad_counter0.n30338 ),
            .carryout(\quad_counter0.n30339 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_12_lut_LC_10_16_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_12_lut_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_12_lut_LC_10_16_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_12_lut_LC_10_16_2  (
            .in0(N__43191),
            .in1(N__43190),
            .in2(N__43586),
            .in3(N__40938),
            .lcout(\quad_counter0.n3009 ),
            .ltout(),
            .carryin(\quad_counter0.n30339 ),
            .carryout(\quad_counter0.n30340 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_13_lut_LC_10_16_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_13_lut_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_13_lut_LC_10_16_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_13_lut_LC_10_16_3  (
            .in0(N__43646),
            .in1(N__43645),
            .in2(N__43590),
            .in3(N__41319),
            .lcout(\quad_counter0.n3008 ),
            .ltout(),
            .carryin(\quad_counter0.n30340 ),
            .carryout(\quad_counter0.n30341 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_14_lut_LC_10_16_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_14_lut_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_14_lut_LC_10_16_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_14_lut_LC_10_16_4  (
            .in0(N__43238),
            .in1(N__43237),
            .in2(N__43587),
            .in3(N__41292),
            .lcout(\quad_counter0.n3007 ),
            .ltout(),
            .carryin(\quad_counter0.n30341 ),
            .carryout(\quad_counter0.n30342 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_15_lut_LC_10_16_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_15_lut_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_15_lut_LC_10_16_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_15_lut_LC_10_16_5  (
            .in0(N__43151),
            .in1(N__43150),
            .in2(N__43591),
            .in3(N__41268),
            .lcout(\quad_counter0.n3006 ),
            .ltout(),
            .carryin(\quad_counter0.n30342 ),
            .carryout(\quad_counter0.n30343 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_16_lut_LC_10_16_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_16_lut_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_16_lut_LC_10_16_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_16_lut_LC_10_16_6  (
            .in0(N__43382),
            .in1(N__43381),
            .in2(N__43588),
            .in3(N__41235),
            .lcout(\quad_counter0.n3005 ),
            .ltout(),
            .carryin(\quad_counter0.n30343 ),
            .carryout(\quad_counter0.n30344 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_17_lut_LC_10_16_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_17_lut_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_17_lut_LC_10_16_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_17_lut_LC_10_16_7  (
            .in0(N__43131),
            .in1(N__43130),
            .in2(N__43592),
            .in3(N__41208),
            .lcout(\quad_counter0.n3004 ),
            .ltout(),
            .carryin(\quad_counter0.n30344 ),
            .carryout(\quad_counter0.n30345 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_18_lut_LC_10_17_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2018_18_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_18_lut_LC_10_17_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_18_lut_LC_10_17_0  (
            .in0(N__43218),
            .in1(N__43214),
            .in2(N__43593),
            .in3(N__41181),
            .lcout(\quad_counter0.n3003 ),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\quad_counter0.n30346 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2018_19_lut_LC_10_17_1 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_2018_19_lut_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2018_19_lut_LC_10_17_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2018_19_lut_LC_10_17_1  (
            .in0(N__43019),
            .in1(N__43020),
            .in2(N__43594),
            .in3(N__41178),
            .lcout(\quad_counter0.n3002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i113_3_lut_LC_10_17_3 .C_ON=1'b0;
    defparam \c0.i113_3_lut_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i113_3_lut_LC_10_17_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i113_3_lut_LC_10_17_3  (
            .in0(N__42881),
            .in1(N__49073),
            .in2(_gnd_net_),
            .in3(N__49003),
            .lcout(\c0.n99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_10_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_10_17_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i22_LC_10_17_5  (
            .in0(N__42943),
            .in1(N__57945),
            .in2(_gnd_net_),
            .in3(N__41142),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97642),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1987_LC_10_17_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1987_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1987_LC_10_17_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1987_LC_10_17_7  (
            .in0(N__46746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46530),
            .lcout(\c0.n33451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1963_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1963_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1963_LC_10_18_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1963_LC_10_18_0  (
            .in0(N__52103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41491),
            .lcout(\c0.n33473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1369_LC_10_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1369_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1369_LC_10_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1369_LC_10_18_1  (
            .in0(N__41490),
            .in1(N__43831),
            .in2(_gnd_net_),
            .in3(N__52102),
            .lcout(\c0.n18627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_2003_LC_10_18_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_2003_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_2003_LC_10_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i5_4_lut_adj_2003_LC_10_18_2  (
            .in0(N__52104),
            .in1(N__52061),
            .in2(N__52166),
            .in3(N__48845),
            .lcout(\c0.n13_adj_4773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_2004_LC_10_18_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_2004_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_2004_LC_10_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_2004_LC_10_18_3  (
            .in0(N__52062),
            .in1(N__52158),
            .in2(N__48854),
            .in3(N__52105),
            .lcout(\c0.n13_adj_4774 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1338_LC_10_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1338_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1338_LC_10_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1338_LC_10_18_4  (
            .in0(N__43832),
            .in1(N__61452),
            .in2(_gnd_net_),
            .in3(N__49424),
            .lcout(),
            .ltout(\c0.n6_adj_4503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1989_LC_10_18_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1989_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1989_LC_10_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1989_LC_10_18_5  (
            .in0(N__41375),
            .in1(N__41475),
            .in2(N__41364),
            .in3(N__41417),
            .lcout(\c0.n17582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_10_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_10_18_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i22_LC_10_18_6  (
            .in0(N__83891),
            .in1(N__75093),
            .in2(N__80319),
            .in3(N__41492),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97656),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_10_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_10_18_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i21_LC_10_18_7  (
            .in0(N__84121),
            .in1(N__83892),
            .in2(N__41361),
            .in3(N__80273),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97656),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1958_2_lut_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.rx.i1958_2_lut_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1958_2_lut_LC_10_19_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.rx.i1958_2_lut_LC_10_19_0  (
            .in0(N__55563),
            .in1(N__55626),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.n3821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1964_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1964_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1964_LC_10_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1964_LC_10_19_1  (
            .in0(N__46524),
            .in1(N__43836),
            .in2(N__46745),
            .in3(N__41504),
            .lcout(\c0.n33804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1405_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1405_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1405_LC_10_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1405_LC_10_19_2  (
            .in0(N__43837),
            .in1(N__43320),
            .in2(N__52122),
            .in3(N__41493),
            .lcout(\c0.data_out_frame_0__7__N_2744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1988_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1988_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1988_LC_10_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1988_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__41426),
            .in2(_gnd_net_),
            .in3(N__76122),
            .lcout(\c0.n33386 ),
            .ltout(\c0.n33386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1978_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1978_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1978_LC_10_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1978_LC_10_19_4  (
            .in0(N__49433),
            .in1(N__46793),
            .in2(N__41469),
            .in3(N__41451),
            .lcout(\c0.n10_adj_4768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_10_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_10_19_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i25_LC_10_19_6  (
            .in0(N__80865),
            .in1(N__78270),
            .in2(N__41430),
            .in3(N__83958),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_10_19_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i9_LC_10_19_7  (
            .in0(N__83957),
            .in1(N__80866),
            .in2(N__76143),
            .in3(N__87198),
            .lcout(data_in_frame_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1844_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1844_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1844_LC_10_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1844_LC_10_20_1  (
            .in0(N__52523),
            .in1(N__44311),
            .in2(_gnd_net_),
            .in3(N__46463),
            .lcout(\c0.n33836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1430_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1430_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1430_LC_10_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1430_LC_10_20_2  (
            .in0(N__49569),
            .in1(N__41522),
            .in2(N__41580),
            .in3(N__65273),
            .lcout(\c0.n7_adj_4554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1985_LC_10_20_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1985_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1985_LC_10_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1985_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__46864),
            .in2(_gnd_net_),
            .in3(N__41410),
            .lcout(\c0.n33720 ),
            .ltout(\c0.n33720_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1986_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1986_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1986_LC_10_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1986_LC_10_20_4  (
            .in0(N__46789),
            .in1(N__43863),
            .in2(N__41607),
            .in3(N__68093),
            .lcout(\c0.n17559 ),
            .ltout(\c0.n17559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1997_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1997_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1997_LC_10_20_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1997_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41604),
            .in3(N__65272),
            .lcout(\c0.n18544 ),
            .ltout(\c0.n18544_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1857_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1857_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1857_LC_10_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1857_LC_10_20_6  (
            .in0(N__49648),
            .in1(N__41601),
            .in2(N__41586),
            .in3(N__41687),
            .lcout(\c0.n31505 ),
            .ltout(\c0.n31505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1860_LC_10_20_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1860_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1860_LC_10_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1860_LC_10_20_7  (
            .in0(N__43757),
            .in1(N__49689),
            .in2(N__41583),
            .in3(N__41576),
            .lcout(\c0.n32325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1832_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1832_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1832_LC_10_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_1832_LC_10_21_1  (
            .in0(N__44036),
            .in1(N__52604),
            .in2(N__49859),
            .in3(N__41670),
            .lcout(),
            .ltout(\c0.n43_adj_4732_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_LC_10_21_2 .C_ON=1'b0;
    defparam \c0.i27_4_lut_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_LC_10_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i27_4_lut_LC_10_21_2  (
            .in0(N__43689),
            .in1(N__41529),
            .in2(N__41562),
            .in3(N__41637),
            .lcout(\c0.n35077 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1830_LC_10_21_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1830_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1830_LC_10_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1830_LC_10_21_3  (
            .in0(N__65277),
            .in1(N__41559),
            .in2(N__43935),
            .in3(N__43887),
            .lcout(),
            .ltout(\c0.n45_adj_4730_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i26_4_lut_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.i26_4_lut_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i26_4_lut_LC_10_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i26_4_lut_LC_10_21_4  (
            .in0(N__41544),
            .in1(N__41538),
            .in2(N__41532),
            .in3(N__41697),
            .lcout(\c0.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_1827_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_1827_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_1827_LC_10_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_1827_LC_10_21_5  (
            .in0(N__44011),
            .in1(N__41523),
            .in2(N__41916),
            .in3(N__49959),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1434_LC_10_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1434_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1434_LC_10_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1434_LC_10_22_0  (
            .in0(N__50199),
            .in1(N__43782),
            .in2(_gnd_net_),
            .in3(N__52879),
            .lcout(),
            .ltout(\c0.n6_adj_4556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1848_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1848_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1848_LC_10_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1848_LC_10_22_1  (
            .in0(N__46967),
            .in1(N__55995),
            .in2(N__41691),
            .in3(N__43881),
            .lcout(\c0.n31651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1845_LC_10_22_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1845_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1845_LC_10_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1845_LC_10_22_2  (
            .in0(N__43902),
            .in1(N__41861),
            .in2(N__41934),
            .in3(N__41688),
            .lcout(),
            .ltout(\c0.n12_adj_4735_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1846_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1846_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1846_LC_10_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1846_LC_10_22_3  (
            .in0(N__43930),
            .in1(N__46935),
            .in2(N__41676),
            .in3(N__44015),
            .lcout(\c0.n31526 ),
            .ltout(\c0.n31526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1847_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1847_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1847_LC_10_22_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1847_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41673),
            .in3(N__50198),
            .lcout(\c0.n33624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1831_LC_10_22_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1831_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1831_LC_10_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1831_LC_10_22_5  (
            .in0(N__41664),
            .in1(N__50343),
            .in2(N__43971),
            .in3(N__41648),
            .lcout(\c0.n44_adj_4731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1811_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1811_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1811_LC_10_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1811_LC_10_23_0  (
            .in0(N__50577),
            .in1(N__53136),
            .in2(N__47625),
            .in3(N__50080),
            .lcout(\c0.n37_adj_4720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i77_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i77_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i77_LC_10_23_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i77_LC_10_23_3  (
            .in0(N__58366),
            .in1(N__87302),
            .in2(N__84217),
            .in3(N__41930),
            .lcout(\c0.data_in_frame_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97740),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1790_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1790_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1790_LC_10_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1790_LC_10_23_4  (
            .in0(N__50032),
            .in1(N__50079),
            .in2(_gnd_net_),
            .in3(N__41631),
            .lcout(\c0.n33951 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1838_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1838_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1838_LC_10_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1838_LC_10_23_5  (
            .in0(N__41951),
            .in1(N__44140),
            .in2(_gnd_net_),
            .in3(N__41929),
            .lcout(\c0.n33641 ),
            .ltout(\c0.n33641_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1839_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1839_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1839_LC_10_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1839_LC_10_23_6  (
            .in0(N__41904),
            .in1(N__41874),
            .in2(N__41865),
            .in3(N__41862),
            .lcout(\c0.n32298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1435_LC_10_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1435_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1435_LC_10_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1435_LC_10_23_7  (
            .in0(N__46936),
            .in1(N__44141),
            .in2(_gnd_net_),
            .in3(N__61184),
            .lcout(\c0.n6_adj_4557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1820_LC_10_24_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1820_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1820_LC_10_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1820_LC_10_24_0  (
            .in0(N__50252),
            .in1(N__44481),
            .in2(N__47547),
            .in3(N__41742),
            .lcout(),
            .ltout(\c0.n18_adj_4725_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1821_LC_10_24_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1821_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1821_LC_10_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1821_LC_10_24_1  (
            .in0(N__44112),
            .in1(N__41832),
            .in2(N__41826),
            .in3(N__48906),
            .lcout(),
            .ltout(\c0.n20_adj_4727_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1822_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1822_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1822_LC_10_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1822_LC_10_24_2  (
            .in0(N__41822),
            .in1(N__41808),
            .in2(N__41796),
            .in3(N__41793),
            .lcout(\c0.n6227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1900_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1900_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1900_LC_10_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1900_LC_10_24_4  (
            .in0(N__55734),
            .in1(N__50151),
            .in2(_gnd_net_),
            .in3(N__41763),
            .lcout(\c0.n33723 ),
            .ltout(\c0.n33723_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1385_LC_10_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1385_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1385_LC_10_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1385_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(N__50251),
            .in2(N__41736),
            .in3(N__41733),
            .lcout(),
            .ltout(\c0.n6_adj_4539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1901_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1901_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1901_LC_10_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1901_LC_10_24_6  (
            .in0(N__44505),
            .in1(N__42033),
            .in2(N__42012),
            .in3(N__47208),
            .lcout(\c0.n18582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i156_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i156_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i156_LC_10_25_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i156_LC_10_25_0  (
            .in0(N__78208),
            .in1(N__78963),
            .in2(N__53318),
            .in3(N__73041),
            .lcout(\c0.data_in_frame_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97773),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1793_LC_10_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1793_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1793_LC_10_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1793_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__47536),
            .in2(_gnd_net_),
            .in3(N__47360),
            .lcout(\c0.n19199 ),
            .ltout(\c0.n19199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1817_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1817_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1817_LC_10_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1817_LC_10_25_2  (
            .in0(N__53311),
            .in1(N__47589),
            .in2(N__42009),
            .in3(N__53241),
            .lcout(\c0.n22_adj_4723 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i68_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i68_LC_10_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i68_LC_10_25_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i68_LC_10_25_3  (
            .in0(N__78962),
            .in1(N__58405),
            .in2(N__81203),
            .in3(N__50126),
            .lcout(\c0.data_in_frame_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97773),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_10_25_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i27_LC_10_25_4  (
            .in0(N__78209),
            .in1(N__83959),
            .in2(N__46868),
            .in3(N__80664),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97773),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1875_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1875_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1875_LC_10_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1875_LC_10_25_5  (
            .in0(N__42006),
            .in1(N__50313),
            .in2(N__41976),
            .in3(N__53494),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i155_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i155_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i155_LC_10_25_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i155_LC_10_25_6  (
            .in0(N__78207),
            .in1(N__73040),
            .in2(N__65521),
            .in3(N__80663),
            .lcout(\c0.data_in_frame_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97773),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadB_I_0_91_2_lut_LC_11_5_0 .C_ON=1'b0;
    defparam \quad_counter1.quadB_I_0_91_2_lut_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.quadB_I_0_91_2_lut_LC_11_5_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \quad_counter1.quadB_I_0_91_2_lut_LC_11_5_0  (
            .in0(N__42147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42118),
            .lcout(\quad_counter1.b_delay_counter_15__N_4237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.quadA_delayed_70_LC_11_5_4 .C_ON=1'b0;
    defparam \quad_counter1.quadA_delayed_70_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.quadA_delayed_70_LC_11_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter1.quadA_delayed_70_LC_11_5_4  (
            .in0(N__44597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(quadA_delayed_adj_4812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97541),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_2060_LC_11_5_5.C_ON=1'b0;
    defparam i1_3_lut_adj_2060_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_2060_LC_11_5_5.LUT_INIT=16'b1111111101100110;
    LogicCell40 i1_3_lut_adj_2060_LC_11_5_5 (
            .in0(N__42119),
            .in1(N__42145),
            .in2(_gnd_net_),
            .in3(N__42101),
            .lcout(n19463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_74_LC_11_5_6 .C_ON=1'b0;
    defparam \quad_counter1.B_74_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_74_LC_11_5_6 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \quad_counter1.B_74_LC_11_5_6  (
            .in0(N__42146),
            .in1(N__42120),
            .in2(N__42105),
            .in3(N__59386),
            .lcout(B_filtered_adj_4810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97541),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1273_LC_11_6_0 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1273_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1273_LC_11_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1273_LC_11_6_0  (
            .in0(N__42525),
            .in1(N__42543),
            .in2(N__42186),
            .in3(N__42218),
            .lcout(),
            .ltout(\quad_counter1.n26_adj_4447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_adj_1276_LC_11_6_1 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_adj_1276_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_adj_1276_LC_11_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_adj_1276_LC_11_6_1  (
            .in0(N__42081),
            .in1(N__42093),
            .in2(N__42108),
            .in3(N__42087),
            .lcout(n17983),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1274_LC_11_6_2 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1274_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1274_LC_11_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1274_LC_11_6_2  (
            .in0(N__42471),
            .in1(N__42507),
            .in2(N__42204),
            .in3(N__42450),
            .lcout(\quad_counter1.n27_adj_4448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1275_LC_11_6_3 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1275_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1275_LC_11_6_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1275_LC_11_6_3  (
            .in0(N__42263),
            .in1(N__42165),
            .in2(N__42075),
            .in3(N__42248),
            .lcout(\quad_counter1.n25_adj_4449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1272_LC_11_6_4 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1272_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1272_LC_11_6_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1272_LC_11_6_4  (
            .in0(N__42278),
            .in1(N__42489),
            .in2(N__42057),
            .in3(N__42233),
            .lcout(\quad_counter1.n28_adj_4446 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.b_delay_counter__i0_LC_11_7_0 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i0_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i0_LC_11_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__42074),
            .in2(_gnd_net_),
            .in3(N__42060),
            .lcout(\quad_counter1.b_delay_counter_0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\quad_counter1.n30031 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i1_LC_11_7_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i1_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i1_LC_11_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i1_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__42056),
            .in2(_gnd_net_),
            .in3(N__42042),
            .lcout(\quad_counter1.b_delay_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n30031 ),
            .carryout(\quad_counter1.n30032 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i2_LC_11_7_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i2_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i2_LC_11_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__42279),
            .in2(_gnd_net_),
            .in3(N__42267),
            .lcout(\quad_counter1.b_delay_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n30032 ),
            .carryout(\quad_counter1.n30033 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i3_LC_11_7_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i3_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i3_LC_11_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i3_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__42264),
            .in2(_gnd_net_),
            .in3(N__42252),
            .lcout(\quad_counter1.b_delay_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n30033 ),
            .carryout(\quad_counter1.n30034 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i4_LC_11_7_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i4_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i4_LC_11_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i4_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__42249),
            .in2(_gnd_net_),
            .in3(N__42237),
            .lcout(\quad_counter1.b_delay_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n30034 ),
            .carryout(\quad_counter1.n30035 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i5_LC_11_7_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i5_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i5_LC_11_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i5_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__42234),
            .in2(_gnd_net_),
            .in3(N__42222),
            .lcout(\quad_counter1.b_delay_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n30035 ),
            .carryout(\quad_counter1.n30036 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i6_LC_11_7_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i6_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i6_LC_11_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i6_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__42219),
            .in2(_gnd_net_),
            .in3(N__42207),
            .lcout(\quad_counter1.b_delay_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n30036 ),
            .carryout(\quad_counter1.n30037 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i7_LC_11_7_7 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i7_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i7_LC_11_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i7_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__42203),
            .in2(_gnd_net_),
            .in3(N__42189),
            .lcout(\quad_counter1.b_delay_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n30037 ),
            .carryout(\quad_counter1.n30038 ),
            .clk(N__97547),
            .ce(N__42431),
            .sr(N__42410));
    defparam \quad_counter1.b_delay_counter__i8_LC_11_8_0 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i8_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i8_LC_11_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i8_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__42182),
            .in2(_gnd_net_),
            .in3(N__42168),
            .lcout(\quad_counter1.b_delay_counter_8 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\quad_counter1.n30039 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i9_LC_11_8_1 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i9_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i9_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i9_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__42164),
            .in2(_gnd_net_),
            .in3(N__42150),
            .lcout(\quad_counter1.b_delay_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n30039 ),
            .carryout(\quad_counter1.n30040 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i10_LC_11_8_2 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i10_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i10_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i10_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__42542),
            .in2(_gnd_net_),
            .in3(N__42528),
            .lcout(\quad_counter1.b_delay_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n30040 ),
            .carryout(\quad_counter1.n30041 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i11_LC_11_8_3 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i11_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i11_LC_11_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i11_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__42524),
            .in2(_gnd_net_),
            .in3(N__42510),
            .lcout(\quad_counter1.b_delay_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n30041 ),
            .carryout(\quad_counter1.n30042 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i12_LC_11_8_4 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i12_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i12_LC_11_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i12_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__42506),
            .in2(_gnd_net_),
            .in3(N__42492),
            .lcout(\quad_counter1.b_delay_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n30042 ),
            .carryout(\quad_counter1.n30043 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i13_LC_11_8_5 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i13_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i13_LC_11_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i13_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__42488),
            .in2(_gnd_net_),
            .in3(N__42474),
            .lcout(\quad_counter1.b_delay_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n30043 ),
            .carryout(\quad_counter1.n30044 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i14_LC_11_8_6 .C_ON=1'b1;
    defparam \quad_counter1.b_delay_counter__i14_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i14_LC_11_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i14_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__42470),
            .in2(_gnd_net_),
            .in3(N__42456),
            .lcout(\quad_counter1.b_delay_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n30044 ),
            .carryout(\quad_counter1.n30045 ),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter1.b_delay_counter__i15_LC_11_8_7 .C_ON=1'b0;
    defparam \quad_counter1.b_delay_counter__i15_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.b_delay_counter__i15_LC_11_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.b_delay_counter__i15_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__42449),
            .in2(_gnd_net_),
            .in3(N__42453),
            .lcout(\quad_counter1.b_delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97553),
            .ce(N__42435),
            .sr(N__42414));
    defparam \quad_counter0.i23581_2_lut_LC_11_9_1 .C_ON=1'b0;
    defparam \quad_counter0.i23581_2_lut_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23581_2_lut_LC_11_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23581_2_lut_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__59881),
            .in2(_gnd_net_),
            .in3(N__42388),
            .lcout(),
            .ltout(\quad_counter0.n28297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1171_LC_11_9_2 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1171_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1171_LC_11_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1171_LC_11_9_2  (
            .in0(N__42364),
            .in1(N__42340),
            .in2(N__42318),
            .in3(N__42313),
            .lcout(\quad_counter0.n10_adj_4357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23591_2_lut_LC_11_9_3 .C_ON=1'b0;
    defparam \quad_counter0.i23591_2_lut_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23591_2_lut_LC_11_9_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23591_2_lut_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__59795),
            .in2(_gnd_net_),
            .in3(N__42843),
            .lcout(\quad_counter0.n28307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1193_LC_11_9_4 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1193_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1193_LC_11_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1193_LC_11_9_4  (
            .in0(N__60391),
            .in1(N__60349),
            .in2(N__60435),
            .in3(N__60475),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1194_LC_11_9_5 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1194_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1194_LC_11_9_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1194_LC_11_9_5  (
            .in0(N__60307),
            .in1(N__60025),
            .in2(N__42816),
            .in3(N__60511),
            .lcout(\quad_counter0.n1847 ),
            .ltout(\quad_counter0.n1847_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30731_1_lut_LC_11_9_6 .C_ON=1'b0;
    defparam \quad_counter0.i30731_1_lut_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30731_1_lut_LC_11_9_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30731_1_lut_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42813),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30713_1_lut_LC_11_10_5 .C_ON=1'b0;
    defparam \quad_counter0.i30713_1_lut_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30713_1_lut_LC_11_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30713_1_lut_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45121),
            .lcout(\quad_counter0.n36140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.r_Bit_Index_1__bdd_4_lut_LC_11_11_5 .C_ON=1'b0;
    defparam \c0.r_Bit_Index_1__bdd_4_lut_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.r_Bit_Index_1__bdd_4_lut_LC_11_11_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.r_Bit_Index_1__bdd_4_lut_LC_11_11_5  (
            .in0(N__71616),
            .in1(N__42742),
            .in2(N__55050),
            .in3(N__42807),
            .lcout(\c0.n36167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36167_bdd_4_lut_LC_11_12_0 .C_ON=1'b0;
    defparam \c0.n36167_bdd_4_lut_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \c0.n36167_bdd_4_lut_LC_11_12_0 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \c0.n36167_bdd_4_lut_LC_11_12_0  (
            .in0(N__51252),
            .in1(N__42771),
            .in2(N__42747),
            .in3(N__42678),
            .lcout(\c0.n36170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1536_LC_11_12_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1536_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1536_LC_11_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_1536_LC_11_12_5  (
            .in0(N__45082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42658),
            .lcout(\c0.n32730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1163_LC_11_12_6 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1163_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1163_LC_11_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1163_LC_11_12_6  (
            .in0(N__42637),
            .in1(N__42613),
            .in2(N__42591),
            .in3(N__42564),
            .lcout(\quad_counter0.n10_adj_4349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_11_12_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_11_12_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_11_12_7  (
            .in0(N__71666),
            .in1(N__71154),
            .in2(N__42965),
            .in3(N__55023),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97578),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_11_13_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_11_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i30_LC_11_13_0  (
            .in0(N__75084),
            .in1(N__57870),
            .in2(_gnd_net_),
            .in3(N__42933),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97584),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_11_13_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_11_13_1 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_11_13_1  (
            .in0(N__42899),
            .in1(N__51396),
            .in2(N__71159),
            .in3(N__71651),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97584),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1733_LC_11_13_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1733_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1733_LC_11_13_5 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1733_LC_11_13_5  (
            .in0(N__92600),
            .in1(N__51377),
            .in2(_gnd_net_),
            .in3(N__49278),
            .lcout(\c0.n11057 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_2_lut_LC_11_14_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_2_lut_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_2_lut_LC_11_14_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1951_2_lut_LC_11_14_0  (
            .in0(N__59721),
            .in1(N__59720),
            .in2(N__43279),
            .in3(N__42858),
            .lcout(\quad_counter0.n2919 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\quad_counter0.n30314 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_3_lut_LC_11_14_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_3_lut_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_3_lut_LC_11_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_3_lut_LC_11_14_1  (
            .in0(N__45473),
            .in1(N__45472),
            .in2(N__45560),
            .in3(N__42855),
            .lcout(\quad_counter0.n2918 ),
            .ltout(),
            .carryin(\quad_counter0.n30314 ),
            .carryout(\quad_counter0.n30315 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_4_lut_LC_11_14_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_4_lut_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_4_lut_LC_11_14_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1951_4_lut_LC_11_14_2  (
            .in0(N__45431),
            .in1(N__45430),
            .in2(N__43280),
            .in3(N__42852),
            .lcout(\quad_counter0.n2917 ),
            .ltout(),
            .carryin(\quad_counter0.n30315 ),
            .carryout(\quad_counter0.n30316 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_5_lut_LC_11_14_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_5_lut_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_5_lut_LC_11_14_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1951_5_lut_LC_11_14_3  (
            .in0(N__45452),
            .in1(N__45451),
            .in2(N__43283),
            .in3(N__42849),
            .lcout(\quad_counter0.n2916 ),
            .ltout(),
            .carryin(\quad_counter0.n30316 ),
            .carryout(\quad_counter0.n30317 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_6_lut_LC_11_14_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_6_lut_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_6_lut_LC_11_14_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1951_6_lut_LC_11_14_4  (
            .in0(N__45386),
            .in1(N__45385),
            .in2(N__43281),
            .in3(N__42846),
            .lcout(\quad_counter0.n2915 ),
            .ltout(),
            .carryin(\quad_counter0.n30317 ),
            .carryout(\quad_counter0.n30318 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_7_lut_LC_11_14_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_7_lut_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_7_lut_LC_11_14_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1951_7_lut_LC_11_14_5  (
            .in0(N__45365),
            .in1(N__45364),
            .in2(N__43284),
            .in3(N__42993),
            .lcout(\quad_counter0.n2914 ),
            .ltout(),
            .carryin(\quad_counter0.n30318 ),
            .carryout(\quad_counter0.n30319 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_8_lut_LC_11_14_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_8_lut_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_8_lut_LC_11_14_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1951_8_lut_LC_11_14_6  (
            .in0(N__45407),
            .in1(N__45406),
            .in2(N__43282),
            .in3(N__42990),
            .lcout(\quad_counter0.n2913 ),
            .ltout(),
            .carryin(\quad_counter0.n30319 ),
            .carryout(\quad_counter0.n30320 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_9_lut_LC_11_14_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_9_lut_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_9_lut_LC_11_14_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_9_lut_LC_11_14_7  (
            .in0(N__45758),
            .in1(N__45757),
            .in2(N__45561),
            .in3(N__42987),
            .lcout(\quad_counter0.n2912 ),
            .ltout(),
            .carryin(\quad_counter0.n30320 ),
            .carryout(\quad_counter0.n30321 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_10_lut_LC_11_15_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_10_lut_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_10_lut_LC_11_15_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_10_lut_LC_11_15_0  (
            .in0(N__45663),
            .in1(N__45659),
            .in2(N__45552),
            .in3(N__42984),
            .lcout(\quad_counter0.n2911 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\quad_counter0.n30322 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_11_lut_LC_11_15_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_11_lut_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_11_lut_LC_11_15_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_11_lut_LC_11_15_1  (
            .in0(N__45738),
            .in1(N__45737),
            .in2(N__45556),
            .in3(N__42981),
            .lcout(\quad_counter0.n2910 ),
            .ltout(),
            .carryin(\quad_counter0.n30322 ),
            .carryout(\quad_counter0.n30323 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_12_lut_LC_11_15_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_12_lut_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_12_lut_LC_11_15_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_12_lut_LC_11_15_2  (
            .in0(N__45719),
            .in1(N__45718),
            .in2(N__45553),
            .in3(N__42978),
            .lcout(\quad_counter0.n2909 ),
            .ltout(),
            .carryin(\quad_counter0.n30323 ),
            .carryout(\quad_counter0.n30324 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_13_lut_LC_11_15_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_13_lut_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_13_lut_LC_11_15_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_13_lut_LC_11_15_3  (
            .in0(N__45342),
            .in1(N__45341),
            .in2(N__45557),
            .in3(N__42975),
            .lcout(\quad_counter0.n2908 ),
            .ltout(),
            .carryin(\quad_counter0.n30324 ),
            .carryout(\quad_counter0.n30325 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_14_lut_LC_11_15_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_14_lut_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_14_lut_LC_11_15_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_14_lut_LC_11_15_4  (
            .in0(N__45681),
            .in1(N__45680),
            .in2(N__45554),
            .in3(N__42972),
            .lcout(\quad_counter0.n2907 ),
            .ltout(),
            .carryin(\quad_counter0.n30325 ),
            .carryout(\quad_counter0.n30326 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_15_lut_LC_11_15_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_15_lut_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_15_lut_LC_11_15_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_15_lut_LC_11_15_5  (
            .in0(N__45699),
            .in1(N__45698),
            .in2(N__45558),
            .in3(N__42969),
            .lcout(\quad_counter0.n2906 ),
            .ltout(),
            .carryin(\quad_counter0.n30326 ),
            .carryout(\quad_counter0.n30327 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_16_lut_LC_11_15_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_16_lut_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_16_lut_LC_11_15_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_16_lut_LC_11_15_6  (
            .in0(N__45588),
            .in1(N__45587),
            .in2(N__45555),
            .in3(N__43293),
            .lcout(\quad_counter0.n2905 ),
            .ltout(),
            .carryin(\quad_counter0.n30327 ),
            .carryout(\quad_counter0.n30328 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_17_lut_LC_11_15_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1951_17_lut_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_17_lut_LC_11_15_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_17_lut_LC_11_15_7  (
            .in0(N__45631),
            .in1(N__45632),
            .in2(N__45559),
            .in3(N__43290),
            .lcout(\quad_counter0.n2904 ),
            .ltout(),
            .carryin(\quad_counter0.n30328 ),
            .carryout(\quad_counter0.n30329 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1951_18_lut_LC_11_16_0 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1951_18_lut_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1951_18_lut_LC_11_16_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1951_18_lut_LC_11_16_0  (
            .in0(N__45612),
            .in1(N__45611),
            .in2(N__45545),
            .in3(N__43287),
            .lcout(\quad_counter0.n2903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30720_1_lut_LC_11_16_1 .C_ON=1'b0;
    defparam \quad_counter0.i30720_1_lut_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30720_1_lut_LC_11_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30720_1_lut_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45512),
            .lcout(\quad_counter0.n36147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i6_2_lut_LC_11_16_4 .C_ON=1'b0;
    defparam \quad_counter0.i6_2_lut_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i6_2_lut_LC_11_16_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i6_2_lut_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43239),
            .in3(N__43207),
            .lcout(\quad_counter0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_LC_11_16_5 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_LC_11_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_LC_11_16_5  (
            .in0(N__43189),
            .in1(N__43173),
            .in2(N__43152),
            .in3(N__43129),
            .lcout(\quad_counter0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23599_2_lut_LC_11_16_6 .C_ON=1'b0;
    defparam \quad_counter0.i23599_2_lut_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23599_2_lut_LC_11_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23599_2_lut_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__59769),
            .in2(_gnd_net_),
            .in3(N__43113),
            .lcout(\quad_counter0.n28315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30718_1_lut_LC_11_16_7 .C_ON=1'b0;
    defparam \quad_counter0.i30718_1_lut_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30718_1_lut_LC_11_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30718_1_lut_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43543),
            .lcout(\quad_counter0.n36145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_LC_11_17_0 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_LC_11_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_LC_11_17_0  (
            .in0(N__43045),
            .in1(N__43018),
            .in2(N__43002),
            .in3(N__43362),
            .lcout(),
            .ltout(\quad_counter0.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_LC_11_17_1 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_LC_11_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_LC_11_17_1  (
            .in0(N__43647),
            .in1(N__43626),
            .in2(N__43605),
            .in3(N__43602),
            .lcout(\quad_counter0.n2936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1162_LC_11_17_3 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1162_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1162_LC_11_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1162_LC_11_17_3  (
            .in0(N__43500),
            .in1(N__43479),
            .in2(N__43458),
            .in3(N__43434),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_4_lut_LC_11_17_4 .C_ON=1'b0;
    defparam \quad_counter0.i1_4_lut_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_4_lut_LC_11_17_4 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i1_4_lut_LC_11_17_4  (
            .in0(N__43428),
            .in1(N__43407),
            .in2(N__43386),
            .in3(N__43383),
            .lcout(\quad_counter0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i61_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i61_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i61_LC_11_17_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i61_LC_11_17_5  (
            .in0(N__83968),
            .in1(N__62149),
            .in2(N__49656),
            .in3(N__84180),
            .lcout(\c0.data_in_frame_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97628),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30377_4_lut_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.i30377_4_lut_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i30377_4_lut_LC_11_18_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i30377_4_lut_LC_11_18_0  (
            .in0(N__49429),
            .in1(N__52064),
            .in2(N__43851),
            .in3(N__52106),
            .lcout(\c0.n35804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1971_LC_11_18_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1971_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1971_LC_11_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1971_LC_11_18_1  (
            .in0(N__43352),
            .in1(N__43329),
            .in2(N__46557),
            .in3(N__43315),
            .lcout(\c0.n30_adj_4765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2001_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2001_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2001_LC_11_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i6_4_lut_adj_2001_LC_11_18_2  (
            .in0(N__43846),
            .in1(N__61453),
            .in2(N__49438),
            .in3(N__46742),
            .lcout(\c0.n14_adj_4771 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_2002_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_2002_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_2002_LC_11_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_2002_LC_11_18_3  (
            .in0(N__46743),
            .in1(N__49428),
            .in2(N__61458),
            .in3(N__43847),
            .lcout(),
            .ltout(\c0.n14_adj_4772_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23003_4_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.i23003_4_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i23003_4_lut_LC_11_18_4 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \c0.i23003_4_lut_LC_11_18_4  (
            .in0(N__43746),
            .in1(N__43740),
            .in2(N__43734),
            .in3(N__43731),
            .lcout(\c0.n27708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_11_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_11_18_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i31_LC_11_18_5  (
            .in0(N__73594),
            .in1(N__78326),
            .in2(N__52396),
            .in3(N__83956),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97643),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_11_18_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i7_LC_11_18_6  (
            .in0(N__81241),
            .in1(N__73595),
            .in2(N__49439),
            .in3(N__83893),
            .lcout(\c0.data_in_frame_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97643),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_11_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_11_18_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i4_LC_11_18_7  (
            .in0(N__78914),
            .in1(N__83955),
            .in2(N__52119),
            .in3(N__81242),
            .lcout(\c0.data_in_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97643),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_11_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_LC_11_19_0  (
            .in0(N__43676),
            .in1(N__49883),
            .in2(N__44269),
            .in3(N__43725),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i90_LC_11_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i90_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i90_LC_11_19_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i90_LC_11_19_2  (
            .in0(N__75343),
            .in1(N__78333),
            .in2(N__43680),
            .in3(N__58302),
            .lcout(\c0.data_in_frame_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_2006_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_2006_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_2006_LC_11_19_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i12_4_lut_adj_2006_LC_11_19_3  (
            .in0(N__48904),
            .in1(N__52354),
            .in2(N__44286),
            .in3(N__44061),
            .lcout(\c0.n29_adj_4776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1867_LC_11_19_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1867_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1867_LC_11_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1867_LC_11_19_4  (
            .in0(N__43675),
            .in1(N__46644),
            .in2(_gnd_net_),
            .in3(N__43664),
            .lcout(\c0.n19102 ),
            .ltout(\c0.n19102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1869_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1869_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1869_LC_11_19_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1869_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43650),
            .in3(N__53226),
            .lcout(\c0.n33954 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i94_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i94_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i94_LC_11_19_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i94_LC_11_19_6  (
            .in0(N__75054),
            .in1(N__58301),
            .in2(N__43934),
            .in3(N__78334),
            .lcout(\c0.data_in_frame_11_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1968_LC_11_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1968_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1968_LC_11_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1968_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__55775),
            .in2(_gnd_net_),
            .in3(N__49310),
            .lcout(\c0.n33582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_1365_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1365_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1365_LC_11_20_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1365_LC_11_20_0  (
            .in0(N__46918),
            .in1(N__43901),
            .in2(N__55407),
            .in3(N__49824),
            .lcout(\c0.n20_adj_4534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1862_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1862_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1862_LC_11_20_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1862_LC_11_20_1  (
            .in0(N__43776),
            .in1(N__46986),
            .in2(_gnd_net_),
            .in3(N__43876),
            .lcout(\c0.n33650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1417_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1417_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1417_LC_11_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1417_LC_11_20_2  (
            .in0(N__43877),
            .in1(N__52605),
            .in2(N__46994),
            .in3(N__43777),
            .lcout(\c0.n15998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1337_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1337_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1337_LC_11_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1337_LC_11_20_4  (
            .in0(N__61438),
            .in1(N__46720),
            .in2(_gnd_net_),
            .in3(N__49434),
            .lcout(\c0.n33311 ),
            .ltout(\c0.n33311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1972_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1972_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1972_LC_11_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1972_LC_11_20_5  (
            .in0(N__46812),
            .in1(N__52389),
            .in2(N__43854),
            .in3(N__43845),
            .lcout(\c0.n31_adj_4766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i96_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i96_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i96_LC_11_20_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i96_LC_11_20_6  (
            .in0(N__58287),
            .in1(N__43778),
            .in2(N__78325),
            .in3(N__80099),
            .lcout(\c0.data_in_frame_11_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i126_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i126_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i126_LC_11_21_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_in_frame_0__i126_LC_11_21_0  (
            .in0(N__58367),
            .in1(N__43987),
            .in2(N__62239),
            .in3(N__74949),
            .lcout(\c0.data_in_frame_15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1856_LC_11_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1856_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1856_LC_11_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1856_LC_11_21_1  (
            .in0(N__44047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49647),
            .lcout(\c0.n33523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i62_LC_11_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i62_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i62_LC_11_21_2 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \c0.data_in_frame_0__i62_LC_11_21_2  (
            .in0(N__74946),
            .in1(N__44049),
            .in2(N__62240),
            .in3(N__83937),
            .lcout(\c0.data_in_frame_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_11_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_11_21_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i6_LC_11_21_3  (
            .in0(N__83936),
            .in1(N__81225),
            .in2(N__46744),
            .in3(N__74947),
            .lcout(\c0.data_in_frame_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1859_LC_11_21_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1859_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1859_LC_11_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1859_LC_11_21_4  (
            .in0(N__49686),
            .in1(N__44060),
            .in2(N__49452),
            .in3(N__44048),
            .lcout(\c0.n31439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1871_LC_11_21_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1871_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1871_LC_11_21_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1871_LC_11_21_5  (
            .in0(N__44153),
            .in1(N__52443),
            .in2(N__43989),
            .in3(N__52976),
            .lcout(\c0.n34003 ),
            .ltout(\c0.n34003_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1874_LC_11_21_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1874_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1874_LC_11_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1874_LC_11_21_6  (
            .in0(N__44037),
            .in1(N__52863),
            .in2(N__44019),
            .in3(N__44016),
            .lcout(\c0.n32_adj_4739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1798_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1798_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1798_LC_11_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1798_LC_11_22_0  (
            .in0(N__43969),
            .in1(N__44186),
            .in2(N__44238),
            .in3(N__52880),
            .lcout(\c0.n12_adj_4714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1761_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1761_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1761_LC_11_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1761_LC_11_22_2  (
            .in0(N__43941),
            .in1(N__43988),
            .in2(N__44208),
            .in3(N__50037),
            .lcout(\c0.n33601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1506_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1506_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1506_LC_11_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1506_LC_11_22_3  (
            .in0(N__44270),
            .in1(N__43970),
            .in2(_gnd_net_),
            .in3(N__46423),
            .lcout(\c0.n18847 ),
            .ltout(\c0.n18847_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1759_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1759_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1759_LC_11_22_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i2_2_lut_adj_1759_LC_11_22_4  (
            .in0(N__47237),
            .in1(_gnd_net_),
            .in2(N__43944),
            .in3(_gnd_net_),
            .lcout(\c0.n10_adj_4708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1505_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1505_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1505_LC_11_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1505_LC_11_22_5  (
            .in0(N__44271),
            .in1(N__44237),
            .in2(_gnd_net_),
            .in3(N__46424),
            .lcout(\c0.n33729 ),
            .ltout(\c0.n33729_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_3_lut_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_3_lut_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_3_lut_LC_11_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i6_4_lut_3_lut_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__68523),
            .in2(N__44211),
            .in3(N__44187),
            .lcout(\c0.n14_adj_4582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_11_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_11_22_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i24_LC_11_22_7  (
            .in0(N__80098),
            .in1(N__83960),
            .in2(N__80366),
            .in3(N__46785),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97705),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1872_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1872_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1872_LC_11_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1872_LC_11_23_0  (
            .in0(N__44199),
            .in1(N__52772),
            .in2(N__56075),
            .in3(N__44180),
            .lcout(\c0.n30_adj_4737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1472_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1472_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1472_LC_11_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1472_LC_11_23_2  (
            .in0(N__50082),
            .in1(N__55733),
            .in2(N__56076),
            .in3(N__59220),
            .lcout(\c0.n33554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1812_LC_11_23_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1812_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1812_LC_11_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1812_LC_11_23_3  (
            .in0(N__53625),
            .in1(N__53550),
            .in2(N__62451),
            .in3(N__56329),
            .lcout(\c0.n35_adj_4721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1863_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1863_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1863_LC_11_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1863_LC_11_23_4  (
            .in0(N__62007),
            .in1(N__52482),
            .in2(_gnd_net_),
            .in3(N__44157),
            .lcout(\c0.n33647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1850_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1850_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1850_LC_11_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1850_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__44142),
            .in2(_gnd_net_),
            .in3(N__61185),
            .lcout(),
            .ltout(\c0.n33908_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1873_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1873_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1873_LC_11_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_1873_LC_11_23_6  (
            .in0(N__52652),
            .in1(N__44111),
            .in2(N__44070),
            .in3(N__44067),
            .lcout(\c0.n34_adj_4738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i67_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i67_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i67_LC_11_24_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i67_LC_11_24_0  (
            .in0(N__80712),
            .in1(N__81221),
            .in2(N__49739),
            .in3(N__58377),
            .lcout(\c0.data_in_frame_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97741),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i121_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i121_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i121_LC_11_24_1 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \c0.data_in_frame_0__i121_LC_11_24_1  (
            .in0(N__44358),
            .in1(N__58368),
            .in2(N__62254),
            .in3(N__80906),
            .lcout(\c0.data_in_frame_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97741),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1413_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1413_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1413_LC_11_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1413_LC_11_24_2  (
            .in0(N__44357),
            .in1(N__44345),
            .in2(_gnd_net_),
            .in3(N__44449),
            .lcout(\c0.n34012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1888_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1888_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1888_LC_11_24_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1888_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__50301),
            .in2(_gnd_net_),
            .in3(N__49732),
            .lcout(\c0.n33871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1388_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1388_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1388_LC_11_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1388_LC_11_24_6  (
            .in0(N__52823),
            .in1(N__44346),
            .in2(_gnd_net_),
            .in3(N__53055),
            .lcout(\c0.n33886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i138_LC_11_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i138_LC_11_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i138_LC_11_24_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i138_LC_11_24_7  (
            .in0(N__73027),
            .in1(N__87139),
            .in2(N__50388),
            .in3(N__75370),
            .lcout(\c0.data_in_frame_17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97741),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1996_LC_11_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1996_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1996_LC_11_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1996_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__52524),
            .in2(_gnd_net_),
            .in3(N__44319),
            .lcout(\c0.n18511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i137_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i137_LC_11_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i137_LC_11_25_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i137_LC_11_25_2  (
            .in0(N__73028),
            .in1(N__53431),
            .in2(N__87199),
            .in3(N__80933),
            .lcout(\c0.data_in_frame_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97759),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1814_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1814_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1814_LC_11_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1814_LC_11_25_3  (
            .in0(N__53548),
            .in1(N__53510),
            .in2(_gnd_net_),
            .in3(N__53455),
            .lcout(),
            .ltout(\c0.n33824_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1816_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1816_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1816_LC_11_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1816_LC_11_25_4  (
            .in0(N__47069),
            .in1(N__44412),
            .in2(N__44403),
            .in3(N__50541),
            .lcout(),
            .ltout(\c0.n24_adj_4722_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1818_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1818_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1818_LC_11_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1818_LC_11_25_5  (
            .in0(N__50612),
            .in1(N__50448),
            .in2(N__44400),
            .in3(N__47561),
            .lcout(),
            .ltout(\c0.n26_adj_4724_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1819_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1819_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1819_LC_11_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1819_LC_11_25_6  (
            .in0(N__46995),
            .in1(N__53430),
            .in2(N__44397),
            .in3(N__44394),
            .lcout(\c0.n31940 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i141_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i141_LC_11_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i141_LC_11_26_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i141_LC_11_26_0  (
            .in0(N__44476),
            .in1(N__84221),
            .in2(N__87169),
            .in3(N__73025),
            .lcout(\c0.data_in_frame_17_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i161_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i161_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i161_LC_11_26_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i161_LC_11_26_1  (
            .in0(N__73022),
            .in1(N__80931),
            .in2(N__47478),
            .in3(N__73941),
            .lcout(\c0.data_in_frame_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i142_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i142_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i142_LC_11_26_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i142_LC_11_26_2  (
            .in0(N__87105),
            .in1(N__73024),
            .in2(N__47543),
            .in3(N__75079),
            .lcout(\c0.data_in_frame_17_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1454_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1454_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1454_LC_11_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1454_LC_11_26_3  (
            .in0(N__44496),
            .in1(N__50375),
            .in2(_gnd_net_),
            .in3(N__44475),
            .lcout(\c0.n33356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i139_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i139_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i139_LC_11_26_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i139_LC_11_26_4  (
            .in0(N__80693),
            .in1(N__73023),
            .in2(N__87168),
            .in3(N__44498),
            .lcout(\c0.data_in_frame_17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1877_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1877_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1877_LC_11_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_1877_LC_11_26_5  (
            .in0(N__44385),
            .in1(N__52581),
            .in2(N__44379),
            .in3(N__44367),
            .lcout(\c0.n17545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1823_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1823_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1823_LC_11_26_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1823_LC_11_26_6  (
            .in0(N__50376),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44497),
            .lcout(\c0.n19060 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i153_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i153_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i153_LC_11_26_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i153_LC_11_26_7  (
            .in0(N__73021),
            .in1(N__78219),
            .in2(N__47493),
            .in3(N__80932),
            .lcout(\c0.data_in_frame_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97774),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i132_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i132_LC_11_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i132_LC_11_27_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i132_LC_11_27_0  (
            .in0(N__73018),
            .in1(N__81279),
            .in2(N__53606),
            .in3(N__78964),
            .lcout(\c0.data_in_frame_16_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97788),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1878_LC_11_27_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1878_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1878_LC_11_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1878_LC_11_27_3  (
            .in0(N__47277),
            .in1(N__62320),
            .in2(_gnd_net_),
            .in3(N__47330),
            .lcout(\c0.n33735 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i160_LC_11_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i160_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i160_LC_11_27_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i160_LC_11_27_4  (
            .in0(N__73019),
            .in1(N__78220),
            .in2(N__80137),
            .in3(N__47644),
            .lcout(\c0.data_in_frame_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97788),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1784_LC_11_27_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1784_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1784_LC_11_27_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1784_LC_11_27_6  (
            .in0(_gnd_net_),
            .in1(N__44477),
            .in2(_gnd_net_),
            .in3(N__44457),
            .lcout(\c0.n33833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i152_LC_11_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i152_LC_11_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i152_LC_11_27_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i152_LC_11_27_7  (
            .in0(N__80386),
            .in1(N__73020),
            .in2(N__50613),
            .in3(N__80127),
            .lcout(\c0.data_in_frame_18_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97788),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23674_2_lut_LC_12_6_2 .C_ON=1'b0;
    defparam \quad_counter0.i23674_2_lut_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23674_2_lut_LC_12_6_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23674_2_lut_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__60061),
            .in2(_gnd_net_),
            .in3(N__54043),
            .lcout(),
            .ltout(\quad_counter0.n28397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1195_LC_12_6_3 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1195_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1195_LC_12_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1195_LC_12_6_3  (
            .in0(N__50707),
            .in1(N__47932),
            .in2(N__44418),
            .in3(N__47866),
            .lcout(\quad_counter0.n10_adj_4377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_2_lut_LC_12_7_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1281_2_lut_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_2_lut_LC_12_7_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1281_2_lut_LC_12_7_0  (
            .in0(N__60027),
            .in1(N__60026),
            .in2(N__44644),
            .in3(N__44415),
            .lcout(\quad_counter0.n1919 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\quad_counter0.n30209 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_3_lut_LC_12_7_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1281_3_lut_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_3_lut_LC_12_7_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1281_3_lut_LC_12_7_1  (
            .in0(N__60519),
            .in1(N__60518),
            .in2(N__44676),
            .in3(N__44664),
            .lcout(\quad_counter0.n1918 ),
            .ltout(),
            .carryin(\quad_counter0.n30209 ),
            .carryout(\quad_counter0.n30210 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_4_lut_LC_12_7_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1281_4_lut_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_4_lut_LC_12_7_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1281_4_lut_LC_12_7_2  (
            .in0(N__60477),
            .in1(N__60476),
            .in2(N__44645),
            .in3(N__44661),
            .lcout(\quad_counter0.n1917 ),
            .ltout(),
            .carryin(\quad_counter0.n30210 ),
            .carryout(\quad_counter0.n30211 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_5_lut_LC_12_7_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1281_5_lut_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_5_lut_LC_12_7_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1281_5_lut_LC_12_7_3  (
            .in0(N__60434),
            .in1(N__60433),
            .in2(N__44648),
            .in3(N__44658),
            .lcout(\quad_counter0.n1916 ),
            .ltout(),
            .carryin(\quad_counter0.n30211 ),
            .carryout(\quad_counter0.n30212 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_6_lut_LC_12_7_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1281_6_lut_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_6_lut_LC_12_7_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1281_6_lut_LC_12_7_4  (
            .in0(N__60393),
            .in1(N__60392),
            .in2(N__44646),
            .in3(N__44655),
            .lcout(\quad_counter0.n1915 ),
            .ltout(),
            .carryin(\quad_counter0.n30212 ),
            .carryout(\quad_counter0.n30213 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_7_lut_LC_12_7_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1281_7_lut_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_7_lut_LC_12_7_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1281_7_lut_LC_12_7_5  (
            .in0(N__60350),
            .in1(N__60351),
            .in2(N__44649),
            .in3(N__44652),
            .lcout(\quad_counter0.n1914 ),
            .ltout(),
            .carryin(\quad_counter0.n30213 ),
            .carryout(\quad_counter0.n30214 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1281_8_lut_LC_12_7_6 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1281_8_lut_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1281_8_lut_LC_12_7_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1281_8_lut_LC_12_7_6  (
            .in0(N__60308),
            .in1(N__60309),
            .in2(N__44647),
            .in3(N__44604),
            .lcout(\quad_counter0.n1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_72_LC_12_8_5 .C_ON=1'b0;
    defparam \quad_counter1.A_72_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_72_LC_12_8_5 .LUT_INIT=16'b1111111000100000;
    LogicCell40 \quad_counter1.A_72_LC_12_8_5  (
            .in0(N__44596),
            .in1(N__44547),
            .in2(N__44538),
            .in3(N__59419),
            .lcout(A_filtered_adj_4809),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97548),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_2_lut_LC_12_9_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_2_lut_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_2_lut_LC_12_9_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2286_2_lut_LC_12_9_0  (
            .in0(N__59916),
            .in1(N__59915),
            .in2(N__44824),
            .in3(N__44511),
            .lcout(\quad_counter0.n3419 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\quad_counter0.n30404 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_3_lut_LC_12_9_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_3_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_3_lut_LC_12_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_3_lut_LC_12_9_1  (
            .in0(N__48015),
            .in1(N__48014),
            .in2(N__45207),
            .in3(N__44508),
            .lcout(\quad_counter0.n3418 ),
            .ltout(),
            .carryin(\quad_counter0.n30404 ),
            .carryout(\quad_counter0.n30405 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_4_lut_LC_12_9_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_4_lut_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_4_lut_LC_12_9_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2286_4_lut_LC_12_9_2  (
            .in0(N__47991),
            .in1(N__47990),
            .in2(N__44825),
            .in3(N__44841),
            .lcout(\quad_counter0.n3417 ),
            .ltout(),
            .carryin(\quad_counter0.n30405 ),
            .carryout(\quad_counter0.n30406 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_5_lut_LC_12_9_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_5_lut_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_5_lut_LC_12_9_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2286_5_lut_LC_12_9_3  (
            .in0(N__47769),
            .in1(N__47768),
            .in2(N__44828),
            .in3(N__44838),
            .lcout(\quad_counter0.n3416 ),
            .ltout(),
            .carryin(\quad_counter0.n30406 ),
            .carryout(\quad_counter0.n30407 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_6_lut_LC_12_9_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_6_lut_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_6_lut_LC_12_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2286_6_lut_LC_12_9_4  (
            .in0(N__47826),
            .in1(N__47825),
            .in2(N__44826),
            .in3(N__44835),
            .lcout(\quad_counter0.n3415 ),
            .ltout(),
            .carryin(\quad_counter0.n30407 ),
            .carryout(\quad_counter0.n30408 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_7_lut_LC_12_9_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_7_lut_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_7_lut_LC_12_9_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2286_7_lut_LC_12_9_5  (
            .in0(N__47804),
            .in1(N__47803),
            .in2(N__44829),
            .in3(N__44832),
            .lcout(\quad_counter0.n3414 ),
            .ltout(),
            .carryin(\quad_counter0.n30408 ),
            .carryout(\quad_counter0.n30409 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_8_lut_LC_12_9_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_8_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_8_lut_LC_12_9_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2286_8_lut_LC_12_9_6  (
            .in0(N__47748),
            .in1(N__47747),
            .in2(N__44827),
            .in3(N__44787),
            .lcout(\quad_counter0.n3413 ),
            .ltout(),
            .carryin(\quad_counter0.n30409 ),
            .carryout(\quad_counter0.n30410 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_9_lut_LC_12_9_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_9_lut_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_9_lut_LC_12_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_9_lut_LC_12_9_7  (
            .in0(N__44784),
            .in1(N__44783),
            .in2(N__45208),
            .in3(N__44757),
            .lcout(\quad_counter0.n3412 ),
            .ltout(),
            .carryin(\quad_counter0.n30410 ),
            .carryout(\quad_counter0.n30411 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_10_lut_LC_12_10_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_10_lut_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_10_lut_LC_12_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_10_lut_LC_12_10_0  (
            .in0(N__44754),
            .in1(N__44753),
            .in2(N__45209),
            .in3(N__44730),
            .lcout(\quad_counter0.n3411 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\quad_counter0.n30412 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_11_lut_LC_12_10_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_11_lut_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_11_lut_LC_12_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_11_lut_LC_12_10_1  (
            .in0(N__44727),
            .in1(N__44726),
            .in2(N__45213),
            .in3(N__44706),
            .lcout(\quad_counter0.n3410 ),
            .ltout(),
            .carryin(\quad_counter0.n30412 ),
            .carryout(\quad_counter0.n30413 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_12_lut_LC_12_10_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_12_lut_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_12_lut_LC_12_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_12_lut_LC_12_10_2  (
            .in0(N__44703),
            .in1(N__44702),
            .in2(N__45210),
            .in3(N__44679),
            .lcout(\quad_counter0.n3409 ),
            .ltout(),
            .carryin(\quad_counter0.n30413 ),
            .carryout(\quad_counter0.n30414 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_13_lut_LC_12_10_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_13_lut_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_13_lut_LC_12_10_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_13_lut_LC_12_10_3  (
            .in0(N__45042),
            .in1(N__45041),
            .in2(N__45214),
            .in3(N__45018),
            .lcout(\quad_counter0.n3408 ),
            .ltout(),
            .carryin(\quad_counter0.n30414 ),
            .carryout(\quad_counter0.n30415 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_14_lut_LC_12_10_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_14_lut_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_14_lut_LC_12_10_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_14_lut_LC_12_10_4  (
            .in0(N__45015),
            .in1(N__45014),
            .in2(N__45211),
            .in3(N__44994),
            .lcout(\quad_counter0.n3407 ),
            .ltout(),
            .carryin(\quad_counter0.n30415 ),
            .carryout(\quad_counter0.n30416 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_15_lut_LC_12_10_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_15_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_15_lut_LC_12_10_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_15_lut_LC_12_10_5  (
            .in0(N__44991),
            .in1(N__44990),
            .in2(N__45215),
            .in3(N__44970),
            .lcout(\quad_counter0.n3406 ),
            .ltout(),
            .carryin(\quad_counter0.n30416 ),
            .carryout(\quad_counter0.n30417 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_16_lut_LC_12_10_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_16_lut_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_16_lut_LC_12_10_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_16_lut_LC_12_10_6  (
            .in0(N__44967),
            .in1(N__44966),
            .in2(N__45212),
            .in3(N__44946),
            .lcout(\quad_counter0.n3405 ),
            .ltout(),
            .carryin(\quad_counter0.n30417 ),
            .carryout(\quad_counter0.n30418 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_17_lut_LC_12_10_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_17_lut_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_17_lut_LC_12_10_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_17_lut_LC_12_10_7  (
            .in0(N__44943),
            .in1(N__44942),
            .in2(N__45216),
            .in3(N__44922),
            .lcout(\quad_counter0.n3404 ),
            .ltout(),
            .carryin(\quad_counter0.n30418 ),
            .carryout(\quad_counter0.n30419 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_18_lut_LC_12_11_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_18_lut_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_18_lut_LC_12_11_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_18_lut_LC_12_11_0  (
            .in0(N__44919),
            .in1(N__44918),
            .in2(N__45217),
            .in3(N__44895),
            .lcout(\quad_counter0.n3403 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\quad_counter0.n30420 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_19_lut_LC_12_11_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_19_lut_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_19_lut_LC_12_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_19_lut_LC_12_11_1  (
            .in0(N__44892),
            .in1(N__44891),
            .in2(N__45220),
            .in3(N__44871),
            .lcout(\quad_counter0.n3402 ),
            .ltout(),
            .carryin(\quad_counter0.n30420 ),
            .carryout(\quad_counter0.n30421 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_20_lut_LC_12_11_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_20_lut_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_20_lut_LC_12_11_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_20_lut_LC_12_11_2  (
            .in0(N__44868),
            .in1(N__44867),
            .in2(N__45218),
            .in3(N__44844),
            .lcout(\quad_counter0.n3401 ),
            .ltout(),
            .carryin(\quad_counter0.n30421 ),
            .carryout(\quad_counter0.n30422 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_21_lut_LC_12_11_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_21_lut_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_21_lut_LC_12_11_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_21_lut_LC_12_11_3  (
            .in0(N__45291),
            .in1(N__45290),
            .in2(N__45221),
            .in3(N__45270),
            .lcout(\quad_counter0.n3400 ),
            .ltout(),
            .carryin(\quad_counter0.n30422 ),
            .carryout(\quad_counter0.n30423 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_22_lut_LC_12_11_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2286_22_lut_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_22_lut_LC_12_11_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_22_lut_LC_12_11_4  (
            .in0(N__45267),
            .in1(N__45266),
            .in2(N__45219),
            .in3(N__45246),
            .lcout(\quad_counter0.n3399 ),
            .ltout(),
            .carryin(\quad_counter0.n30423 ),
            .carryout(\quad_counter0.n30424 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2286_23_lut_LC_12_11_5 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_2286_23_lut_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2286_23_lut_LC_12_11_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2286_23_lut_LC_12_11_5  (
            .in0(N__45242),
            .in1(N__45243),
            .in2(N__45222),
            .in3(N__45093),
            .lcout(\quad_counter0.n3398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i5_LC_12_12_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_12_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_12_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__45083),
            .in2(_gnd_net_),
            .in3(N__71322),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97569),
            .ce(),
            .sr(N__45063));
    defparam \quad_counter0.mod_61_add_1884_2_lut_LC_12_13_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_2_lut_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_2_lut_LC_12_13_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1884_2_lut_LC_12_13_0  (
            .in0(N__59670),
            .in1(N__59669),
            .in2(N__48055),
            .in3(N__45057),
            .lcout(\quad_counter0.n2819 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\quad_counter0.n30299 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_3_lut_LC_12_13_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_3_lut_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_3_lut_LC_12_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_3_lut_LC_12_13_1  (
            .in0(N__50946),
            .in1(N__50945),
            .in2(N__48123),
            .in3(N__45054),
            .lcout(\quad_counter0.n2818 ),
            .ltout(),
            .carryin(\quad_counter0.n30299 ),
            .carryout(\quad_counter0.n30300 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_4_lut_LC_12_13_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_4_lut_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_4_lut_LC_12_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1884_4_lut_LC_12_13_2  (
            .in0(N__50919),
            .in1(N__50918),
            .in2(N__48056),
            .in3(N__45051),
            .lcout(\quad_counter0.n2817 ),
            .ltout(),
            .carryin(\quad_counter0.n30300 ),
            .carryout(\quad_counter0.n30301 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_5_lut_LC_12_13_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_5_lut_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_5_lut_LC_12_13_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1884_5_lut_LC_12_13_3  (
            .in0(N__50892),
            .in1(N__50891),
            .in2(N__48059),
            .in3(N__45048),
            .lcout(\quad_counter0.n2816 ),
            .ltout(),
            .carryin(\quad_counter0.n30301 ),
            .carryout(\quad_counter0.n30302 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_6_lut_LC_12_13_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_6_lut_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_6_lut_LC_12_13_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1884_6_lut_LC_12_13_4  (
            .in0(N__50865),
            .in1(N__50864),
            .in2(N__48057),
            .in3(N__45045),
            .lcout(\quad_counter0.n2815 ),
            .ltout(),
            .carryin(\quad_counter0.n30302 ),
            .carryout(\quad_counter0.n30303 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_7_lut_LC_12_13_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_7_lut_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_7_lut_LC_12_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1884_7_lut_LC_12_13_5  (
            .in0(N__51204),
            .in1(N__51203),
            .in2(N__48060),
            .in3(N__45318),
            .lcout(\quad_counter0.n2814 ),
            .ltout(),
            .carryin(\quad_counter0.n30303 ),
            .carryout(\quad_counter0.n30304 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_8_lut_LC_12_13_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_8_lut_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_8_lut_LC_12_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1884_8_lut_LC_12_13_6  (
            .in0(N__51177),
            .in1(N__51176),
            .in2(N__48058),
            .in3(N__45315),
            .lcout(\quad_counter0.n2813 ),
            .ltout(),
            .carryin(\quad_counter0.n30304 ),
            .carryout(\quad_counter0.n30305 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_9_lut_LC_12_13_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_9_lut_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_9_lut_LC_12_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_9_lut_LC_12_13_7  (
            .in0(N__51150),
            .in1(N__51149),
            .in2(N__48124),
            .in3(N__45312),
            .lcout(\quad_counter0.n2812 ),
            .ltout(),
            .carryin(\quad_counter0.n30305 ),
            .carryout(\quad_counter0.n30306 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_10_lut_LC_12_14_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_10_lut_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_10_lut_LC_12_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_10_lut_LC_12_14_0  (
            .in0(N__51123),
            .in1(N__51122),
            .in2(N__48125),
            .in3(N__45309),
            .lcout(\quad_counter0.n2811 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\quad_counter0.n30307 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_11_lut_LC_12_14_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_11_lut_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_11_lut_LC_12_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_11_lut_LC_12_14_1  (
            .in0(N__51096),
            .in1(N__51095),
            .in2(N__48129),
            .in3(N__45306),
            .lcout(\quad_counter0.n2810 ),
            .ltout(),
            .carryin(\quad_counter0.n30307 ),
            .carryout(\quad_counter0.n30308 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_12_lut_LC_12_14_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_12_lut_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_12_lut_LC_12_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_12_lut_LC_12_14_2  (
            .in0(N__51066),
            .in1(N__51065),
            .in2(N__48126),
            .in3(N__45303),
            .lcout(\quad_counter0.n2809 ),
            .ltout(),
            .carryin(\quad_counter0.n30308 ),
            .carryout(\quad_counter0.n30309 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_13_lut_LC_12_14_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_13_lut_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_13_lut_LC_12_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_13_lut_LC_12_14_3  (
            .in0(N__51039),
            .in1(N__51038),
            .in2(N__48130),
            .in3(N__45300),
            .lcout(\quad_counter0.n2808 ),
            .ltout(),
            .carryin(\quad_counter0.n30309 ),
            .carryout(\quad_counter0.n30310 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_14_lut_LC_12_14_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_14_lut_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_14_lut_LC_12_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_14_lut_LC_12_14_4  (
            .in0(N__51012),
            .in1(N__51011),
            .in2(N__48127),
            .in3(N__45297),
            .lcout(\quad_counter0.n2807 ),
            .ltout(),
            .carryin(\quad_counter0.n30310 ),
            .carryout(\quad_counter0.n30311 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_15_lut_LC_12_14_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_15_lut_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_15_lut_LC_12_14_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_15_lut_LC_12_14_5  (
            .in0(N__51348),
            .in1(N__51347),
            .in2(N__48131),
            .in3(N__45294),
            .lcout(\quad_counter0.n2806 ),
            .ltout(),
            .carryin(\quad_counter0.n30311 ),
            .carryout(\quad_counter0.n30312 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_16_lut_LC_12_14_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1884_16_lut_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_16_lut_LC_12_14_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_16_lut_LC_12_14_6  (
            .in0(N__51318),
            .in1(N__51317),
            .in2(N__48128),
            .in3(N__45765),
            .lcout(\quad_counter0.n2805 ),
            .ltout(),
            .carryin(\quad_counter0.n30312 ),
            .carryout(\quad_counter0.n30313 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1884_17_lut_LC_12_14_7 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1884_17_lut_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1884_17_lut_LC_12_14_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1884_17_lut_LC_12_14_7  (
            .in0(N__51287),
            .in1(N__51288),
            .in2(N__48132),
            .in3(N__45762),
            .lcout(\quad_counter0.n2804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i7_4_lut_adj_1227_LC_12_15_0 .C_ON=1'b0;
    defparam \quad_counter0.i7_4_lut_adj_1227_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i7_4_lut_adj_1227_LC_12_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i7_4_lut_adj_1227_LC_12_15_0  (
            .in0(N__45759),
            .in1(N__45736),
            .in2(N__45720),
            .in3(N__45697),
            .lcout(\quad_counter0.n18_adj_4408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_adj_1228_LC_12_15_1 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_adj_1228_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_adj_1228_LC_12_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_adj_1228_LC_12_15_1  (
            .in0(N__45679),
            .in1(N__45658),
            .in2(N__45633),
            .in3(N__45601),
            .lcout(),
            .ltout(\quad_counter0.n19_adj_4409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1229_LC_12_15_2 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1229_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1229_LC_12_15_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1229_LC_12_15_2  (
            .in0(N__45586),
            .in1(N__45324),
            .in2(N__45570),
            .in3(N__45567),
            .lcout(\quad_counter0.n2837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23607_2_lut_LC_12_15_3 .C_ON=1'b0;
    defparam \quad_counter0.i23607_2_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23607_2_lut_LC_12_15_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i23607_2_lut_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45477),
            .in3(N__59719),
            .lcout(),
            .ltout(\quad_counter0.n28323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1225_LC_12_15_4 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1225_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1225_LC_12_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1225_LC_12_15_4  (
            .in0(N__45453),
            .in1(N__45432),
            .in2(N__45411),
            .in3(N__45408),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_4_lut_adj_1226_LC_12_15_5 .C_ON=1'b0;
    defparam \quad_counter0.i1_4_lut_adj_1226_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_4_lut_adj_1226_LC_12_15_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i1_4_lut_adj_1226_LC_12_15_5  (
            .in0(N__45387),
            .in1(N__45366),
            .in2(N__45345),
            .in3(N__45340),
            .lcout(\quad_counter0.n12_adj_4407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1614_LC_12_16_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1614_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1614_LC_12_16_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1614_LC_12_16_0  (
            .in0(N__45903),
            .in1(N__46058),
            .in2(N__46331),
            .in3(N__46184),
            .lcout(\c0.n32740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i10_LC_12_16_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_12_16_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_12_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__71316),
            .in2(_gnd_net_),
            .in3(N__46327),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97602),
            .ce(),
            .sr(N__46344));
    defparam \c0.i2_3_lut_adj_1948_LC_12_16_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1948_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1948_LC_12_16_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1948_LC_12_16_2  (
            .in0(N__46323),
            .in1(N__46307),
            .in2(_gnd_net_),
            .in3(N__46265),
            .lcout(\c0.n19909 ),
            .ltout(\c0.n19909_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1949_LC_12_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1949_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1949_LC_12_16_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1949_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46248),
            .in3(N__71262),
            .lcout(),
            .ltout(\c0.n34017_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i97_4_lut_LC_12_16_4 .C_ON=1'b0;
    defparam \c0.i97_4_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i97_4_lut_LC_12_16_4 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \c0.i97_4_lut_LC_12_16_4  (
            .in0(N__46245),
            .in1(N__49095),
            .in2(N__46215),
            .in3(N__49272),
            .lcout(\c0.n29675 ),
            .ltout(\c0.n29675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1377_LC_12_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1377_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1377_LC_12_16_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1377_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__51850),
            .in2(N__46212),
            .in3(N__51552),
            .lcout(),
            .ltout(\c0.n81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1954_LC_12_16_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1954_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1954_LC_12_16_6 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \c0.i2_4_lut_adj_1954_LC_12_16_6  (
            .in0(N__51897),
            .in1(N__48633),
            .in2(N__46209),
            .in3(N__51522),
            .lcout(\c0.n1286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1621_LC_12_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1621_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1621_LC_12_16_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1621_LC_12_16_7  (
            .in0(N__46183),
            .in1(N__71263),
            .in2(N__46062),
            .in3(N__45902),
            .lcout(\c0.n32750 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_2008_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_2008_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_2008_LC_12_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_2008_LC_12_17_1  (
            .in0(N__46950),
            .in1(N__46479),
            .in2(N__46470),
            .in3(N__46566),
            .lcout(\c0.n32_adj_4778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i35_3_lut_4_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.i35_3_lut_4_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i35_3_lut_4_lut_LC_12_17_3 .LUT_INIT=16'b1011010110110000;
    LogicCell40 \c0.i35_3_lut_4_lut_LC_12_17_3  (
            .in0(N__51898),
            .in1(N__51953),
            .in2(N__51695),
            .in3(N__84822),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_2007_LC_12_17_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_2007_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_2007_LC_12_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i11_4_lut_adj_2007_LC_12_17_4  (
            .in0(N__46428),
            .in1(N__49761),
            .in2(N__48958),
            .in3(N__61177),
            .lcout(),
            .ltout(\c0.n28_adj_4777_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_2010_LC_12_17_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_2010_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_2010_LC_12_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_2010_LC_12_17_5  (
            .in0(N__46539),
            .in1(N__46392),
            .in2(N__46383),
            .in3(N__46380),
            .lcout(\c0.n27710 ),
            .ltout(\c0.n27710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30605_4_lut_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.i30605_4_lut_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30605_4_lut_LC_12_17_6 .LUT_INIT=16'b1000101100000000;
    LogicCell40 \c0.i30605_4_lut_LC_12_17_6  (
            .in0(N__51234),
            .in1(N__51899),
            .in2(N__46374),
            .in3(N__51851),
            .lcout(),
            .ltout(\c0.n35947_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_5282_LC_12_17_7 .C_ON=1'b0;
    defparam \c0.tx_transmit_5282_LC_12_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_5282_LC_12_17_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \c0.tx_transmit_5282_LC_12_17_7  (
            .in0(N__51750),
            .in1(N__84823),
            .in2(N__46371),
            .in3(N__51686),
            .lcout(r_SM_Main_2_N_3755_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97614),
            .ce(),
            .sr(N__51942));
    defparam \c0.i14_4_lut_adj_2011_LC_12_18_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_2011_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_2011_LC_12_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14_4_lut_adj_2011_LC_12_18_0  (
            .in0(N__76145),
            .in1(N__64828),
            .in2(N__64739),
            .in3(N__58689),
            .lcout(),
            .ltout(\c0.n38_adj_4780_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_2014_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_2014_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_2014_LC_12_18_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.i22_4_lut_adj_2014_LC_12_18_1  (
            .in0(N__46368),
            .in1(N__46758),
            .in2(N__46356),
            .in3(N__46752),
            .lcout(),
            .ltout(\c0.n46_adj_4783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_3_lut_LC_12_18_2 .C_ON=1'b0;
    defparam \c0.i23_3_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i23_3_lut_LC_12_18_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \c0.i23_3_lut_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__46353),
            .in2(N__46347),
            .in3(N__48771),
            .lcout(FRAME_MATCHER_state_31_N_2976_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_2012_LC_12_18_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_2012_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_2012_LC_12_18_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i15_4_lut_adj_2012_LC_12_18_3  (
            .in0(N__46528),
            .in1(N__46794),
            .in2(N__77214),
            .in3(N__61457),
            .lcout(\c0.n39_adj_4781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_2013_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_2013_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_2013_LC_12_18_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.i13_4_lut_adj_2013_LC_12_18_4  (
            .in0(N__72425),
            .in1(N__46741),
            .in2(N__57648),
            .in3(N__83619),
            .lcout(\c0.n37_adj_4782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1979_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1979_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1979_LC_12_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1979_LC_12_18_7  (
            .in0(N__46740),
            .in1(N__46689),
            .in2(_gnd_net_),
            .in3(N__76144),
            .lcout(\c0.n33500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_12_19_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_12_19_0  (
            .in0(N__52569),
            .in1(N__80807),
            .in2(N__55929),
            .in3(N__46677),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97644),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_2005_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_2005_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_2005_LC_12_19_1 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \c0.i9_4_lut_adj_2005_LC_12_19_1  (
            .in0(N__55646),
            .in1(N__46647),
            .in2(N__46578),
            .in3(N__49688),
            .lcout(\c0.n26_adj_4775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1959_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1959_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1959_LC_12_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1959_LC_12_19_3  (
            .in0(N__46556),
            .in1(N__58681),
            .in2(N__46491),
            .in3(N__83618),
            .lcout(\c0.n33291 ),
            .ltout(\c0.n33291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_2009_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_2009_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_2009_LC_12_19_4 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \c0.i2_2_lut_adj_2009_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46542),
            .in3(N__49568),
            .lcout(\c0.n19_adj_4779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_12_19_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i23_LC_12_19_5  (
            .in0(N__83913),
            .in1(N__80422),
            .in2(N__46529),
            .in3(N__73593),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97644),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_12_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_12_19_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i47_LC_12_19_6  (
            .in0(N__78619),
            .in1(N__68307),
            .in2(N__73633),
            .in3(N__46490),
            .lcout(\c0.data_in_frame_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97644),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_12_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_12_19_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i46_LC_12_19_7  (
            .in0(N__68306),
            .in1(N__78620),
            .in2(N__46839),
            .in3(N__75051),
            .lcout(\c0.data_in_frame_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97644),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_12_20_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i56_LC_12_20_0  (
            .in0(N__80111),
            .in1(N__83920),
            .in2(N__89826),
            .in3(N__46928),
            .lcout(\c0.data_in_frame_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1336_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1336_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1336_LC_12_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1336_LC_12_20_1  (
            .in0(N__46814),
            .in1(N__61440),
            .in2(_gnd_net_),
            .in3(N__58688),
            .lcout(),
            .ltout(\c0.n6_adj_4501_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1999_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1999_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1999_LC_12_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1999_LC_12_20_2  (
            .in0(N__49386),
            .in1(N__68217),
            .in2(N__46875),
            .in3(N__46872),
            .lcout(\c0.n18709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_12_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_12_20_3  (
            .in0(N__46813),
            .in1(N__61439),
            .in2(_gnd_net_),
            .in3(N__68092),
            .lcout(),
            .ltout(\c0.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1958_LC_12_20_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1958_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1958_LC_12_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1958_LC_12_20_4  (
            .in0(N__46835),
            .in1(N__55776),
            .in2(N__46824),
            .in3(N__64712),
            .lcout(\c0.n18141 ),
            .ltout(\c0.n18141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1886_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1886_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1886_LC_12_20_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1886_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46821),
            .in3(N__49712),
            .lcout(\c0.n33877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_12_20_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i12_LC_12_20_6  (
            .in0(N__87290),
            .in1(N__83919),
            .in2(N__64738),
            .in3(N__78913),
            .lcout(data_in_frame_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_12_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_12_20_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i28_LC_12_20_7  (
            .in0(N__83918),
            .in1(N__46818),
            .in2(N__78961),
            .in3(N__78331),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1884_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1884_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1884_LC_12_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1884_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__49543),
            .in2(_gnd_net_),
            .in3(N__49682),
            .lcout(),
            .ltout(\c0.n33927_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1885_LC_12_21_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1885_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1885_LC_12_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1885_LC_12_21_1  (
            .in0(N__47123),
            .in1(N__47003),
            .in2(N__47010),
            .in3(N__49754),
            .lcout(\c0.n33708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i83_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i83_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i83_LC_12_21_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i83_LC_12_21_2  (
            .in0(N__58362),
            .in1(N__80408),
            .in2(N__47007),
            .in3(N__80633),
            .lcout(\c0.data_in_frame_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i66_LC_12_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i66_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i66_LC_12_21_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i66_LC_12_21_3  (
            .in0(N__75316),
            .in1(N__81248),
            .in2(N__47127),
            .in3(N__58364),
            .lcout(\c0.data_in_frame_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i82_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i82_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i82_LC_12_21_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i82_LC_12_21_4  (
            .in0(N__58361),
            .in1(N__80407),
            .in2(N__49485),
            .in3(N__75317),
            .lcout(\c0.data_in_frame_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i85_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i85_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i85_LC_12_21_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i85_LC_12_21_5  (
            .in0(N__80406),
            .in1(N__58363),
            .in2(N__49884),
            .in3(N__84171),
            .lcout(\c0.data_in_frame_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1853_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1853_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1853_LC_12_21_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_adj_1853_LC_12_21_6  (
            .in0(N__46990),
            .in1(N__52805),
            .in2(N__47062),
            .in3(N__52743),
            .lcout(\c0.n33417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_12_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_12_21_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i30_LC_12_21_7  (
            .in0(N__74948),
            .in1(N__83953),
            .in2(N__78336),
            .in3(N__49309),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i114_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i114_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i114_LC_12_22_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i114_LC_12_22_0  (
            .in0(N__89823),
            .in1(N__58316),
            .in2(N__46968),
            .in3(N__75319),
            .lcout(\c0.data_in_frame_14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1960_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1960_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1960_LC_12_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1960_LC_12_22_1  (
            .in0(N__52681),
            .in1(N__64829),
            .in2(N__47036),
            .in3(N__49782),
            .lcout(\c0.n2_adj_4741 ),
            .ltout(\c0.n2_adj_4741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1887_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1887_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1887_LC_12_22_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i2_2_lut_adj_1887_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47145),
            .in3(N__49793),
            .lcout(\c0.n33283 ),
            .ltout(\c0.n33283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1889_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1889_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1889_LC_12_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1889_LC_12_22_3  (
            .in0(N__49467),
            .in1(N__47122),
            .in2(N__47106),
            .in3(N__47102),
            .lcout(\c0.n18805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i148_LC_12_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i148_LC_12_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i148_LC_12_22_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i148_LC_12_22_4  (
            .in0(N__78948),
            .in1(N__80423),
            .in2(N__47082),
            .in3(N__73031),
            .lcout(\c0.data_in_frame_18_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1801_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1801_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1801_LC_12_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1801_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__47078),
            .in2(_gnd_net_),
            .in3(N__47168),
            .lcout(\c0.n6_adj_4715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i118_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i118_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i118_LC_12_22_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i118_LC_12_22_6  (
            .in0(N__89824),
            .in1(N__58317),
            .in2(N__47070),
            .in3(N__75052),
            .lcout(\c0.data_in_frame_14_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_12_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_12_22_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_12_22_7  (
            .in0(N__75318),
            .in1(N__89825),
            .in2(N__47037),
            .in3(N__83941),
            .lcout(\c0.data_in_frame_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1841_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1841_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1841_LC_12_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1841_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__47264),
            .in2(_gnd_net_),
            .in3(N__49522),
            .lcout(\c0.n4_adj_4734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1507_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1507_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1507_LC_12_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1507_LC_12_23_1  (
            .in0(N__52653),
            .in1(N__68515),
            .in2(_gnd_net_),
            .in3(N__47022),
            .lcout(\c0.n33880 ),
            .ltout(\c0.n33880_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1804_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1804_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1804_LC_12_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1804_LC_12_23_2  (
            .in0(N__56368),
            .in1(N__50088),
            .in2(N__47013),
            .in3(N__51627),
            .lcout(),
            .ltout(\c0.n12_adj_4716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1805_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1805_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1805_LC_12_23_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1805_LC_12_23_3  (
            .in0(N__49523),
            .in1(N__47304),
            .in2(N__47280),
            .in3(N__47219),
            .lcout(\c0.n33532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1824_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1824_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1824_LC_12_23_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1824_LC_12_23_4  (
            .in0(N__49976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47233),
            .lcout(\c0.n33741 ),
            .ltout(\c0.n33741_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1683_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1683_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1683_LC_12_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1683_LC_12_23_5  (
            .in0(N__47265),
            .in1(N__47374),
            .in2(N__47247),
            .in3(N__47244),
            .lcout(\c0.n10_adj_4697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1807_LC_12_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1807_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1807_LC_12_23_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1807_LC_12_23_6  (
            .in0(N__47164),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55987),
            .lcout(\c0.n33711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i144_LC_12_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i144_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i144_LC_12_23_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i144_LC_12_23_7  (
            .in0(N__80128),
            .in1(N__87305),
            .in2(N__47238),
            .in3(N__73032),
            .lcout(\c0.data_in_frame_17_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97706),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1808_LC_12_24_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1808_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1808_LC_12_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1808_LC_12_24_0  (
            .in0(N__47220),
            .in1(N__47207),
            .in2(N__47379),
            .in3(N__52910),
            .lcout(),
            .ltout(\c0.n34_adj_4718_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1809_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1809_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1809_LC_12_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1809_LC_12_24_1  (
            .in0(N__65522),
            .in1(N__56007),
            .in2(N__47193),
            .in3(N__47385),
            .lcout(),
            .ltout(\c0.n38_adj_4719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_adj_1813_LC_12_24_2 .C_ON=1'b0;
    defparam \c0.i20_4_lut_adj_1813_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_adj_1813_LC_12_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_adj_1813_LC_12_24_2  (
            .in0(N__47190),
            .in1(N__47178),
            .in2(N__47172),
            .in3(N__47661),
            .lcout(\c0.n33972 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i130_LC_12_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i130_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i130_LC_12_24_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i130_LC_12_24_3  (
            .in0(N__75371),
            .in1(N__73029),
            .in2(N__47169),
            .in3(N__81222),
            .lcout(\c0.data_in_frame_16_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97724),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_12_24_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__52722),
            .in2(_gnd_net_),
            .in3(N__47394),
            .lcout(\c0.n24_adj_4717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i145_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i145_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i145_LC_12_24_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i145_LC_12_24_5  (
            .in0(N__80332),
            .in1(N__73030),
            .in2(N__80924),
            .in3(N__47378),
            .lcout(\c0.data_in_frame_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97724),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1762_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1762_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1762_LC_12_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1762_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__47652),
            .in2(_gnd_net_),
            .in3(N__56350),
            .lcout(\c0.n19226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1879_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1879_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1879_LC_12_25_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_adj_1879_LC_12_25_2  (
            .in0(N__56730),
            .in1(N__56114),
            .in2(_gnd_net_),
            .in3(N__47447),
            .lcout(\c0.n33717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1684_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1684_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1684_LC_12_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1684_LC_12_25_3  (
            .in0(N__47361),
            .in1(N__47340),
            .in2(_gnd_net_),
            .in3(N__53031),
            .lcout(\c0.n18588 ),
            .ltout(\c0.n18588_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1678_LC_12_25_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1678_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1678_LC_12_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1678_LC_12_25_4  (
            .in0(N__47331),
            .in1(N__56567),
            .in2(N__47319),
            .in3(N__47316),
            .lcout(\c0.n12_adj_4696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1415_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1415_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1415_LC_12_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1415_LC_12_25_5  (
            .in0(N__53607),
            .in1(N__50511),
            .in2(N__53362),
            .in3(N__53406),
            .lcout(\c0.n33789 ),
            .ltout(\c0.n33789_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1865_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1865_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1865_LC_12_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1865_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__56729),
            .in2(N__47310),
            .in3(N__56113),
            .lcout(\c0.n19108 ),
            .ltout(\c0.n19108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1406_LC_12_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1406_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1406_LC_12_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1406_LC_12_25_7  (
            .in0(_gnd_net_),
            .in1(N__47531),
            .in2(N__47307),
            .in3(N__47684),
            .lcout(\c0.n31589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_12_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_12_26_0  (
            .in0(N__47691),
            .in1(N__47571),
            .in2(_gnd_net_),
            .in3(N__47562),
            .lcout(\c0.n8_adj_4745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1880_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1880_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1880_LC_12_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1880_LC_12_26_1  (
            .in0(_gnd_net_),
            .in1(N__47532),
            .in2(_gnd_net_),
            .in3(N__47683),
            .lcout(),
            .ltout(\c0.n6242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1903_LC_12_26_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1903_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1903_LC_12_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1903_LC_12_26_2  (
            .in0(N__47409),
            .in1(N__47505),
            .in2(N__47499),
            .in3(N__47417),
            .lcout(\c0.n33665 ),
            .ltout(\c0.n33665_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1815_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1815_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1815_LC_12_26_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1815_LC_12_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47496),
            .in3(N__47489),
            .lcout(\c0.n33942 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1763_LC_12_26_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1763_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1763_LC_12_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1763_LC_12_26_4  (
            .in0(N__47432),
            .in1(N__47474),
            .in2(N__47463),
            .in3(N__47448),
            .lcout(\c0.n33514 ),
            .ltout(\c0.n33514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1770_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1770_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1770_LC_12_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1770_LC_12_26_5  (
            .in0(N__50393),
            .in1(N__59352),
            .in2(N__47436),
            .in3(N__50418),
            .lcout(\c0.n10_adj_4709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1679_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1679_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1679_LC_12_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1679_LC_12_26_6  (
            .in0(N__47433),
            .in1(N__47424),
            .in2(N__47610),
            .in3(N__47418),
            .lcout(\c0.n32341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i154_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i154_LC_12_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i154_LC_12_27_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i154_LC_12_27_0  (
            .in0(N__75358),
            .in1(N__73016),
            .in2(N__78327),
            .in3(N__47408),
            .lcout(\c0.data_in_frame_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1386_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1386_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1386_LC_12_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1386_LC_12_27_1  (
            .in0(N__50598),
            .in1(N__47582),
            .in2(_gnd_net_),
            .in3(N__53715),
            .lcout(\c0.n33308 ),
            .ltout(\c0.n33308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1810_LC_12_27_2 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1810_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1810_LC_12_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_1810_LC_12_27_2  (
            .in0(N__47685),
            .in1(N__50481),
            .in2(N__47664),
            .in3(N__56456),
            .lcout(\c0.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i136_LC_12_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i136_LC_12_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i136_LC_12_27_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i136_LC_12_27_3  (
            .in0(N__73013),
            .in1(N__80102),
            .in2(N__53361),
            .in3(N__81202),
            .lcout(\c0.data_in_frame_16_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i168_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i168_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i168_LC_12_27_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i168_LC_12_27_4  (
            .in0(N__80101),
            .in1(N__53803),
            .in2(N__73949),
            .in3(N__73017),
            .lcout(\c0.data_in_frame_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1495_LC_12_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1495_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1495_LC_12_27_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1495_LC_12_27_5  (
            .in0(N__47645),
            .in1(N__53436),
            .in2(_gnd_net_),
            .in3(N__53153),
            .lcout(\c0.n22_adj_4574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i134_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i134_LC_12_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i134_LC_12_27_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i134_LC_12_27_6  (
            .in0(N__74992),
            .in1(N__73015),
            .in2(N__59151),
            .in3(N__81201),
            .lcout(\c0.data_in_frame_16_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i162_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i162_LC_12_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i162_LC_12_27_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i162_LC_12_27_7  (
            .in0(N__73014),
            .in1(N__73937),
            .in2(N__47609),
            .in3(N__75359),
            .lcout(\c0.data_in_frame_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1389_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1389_LC_12_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1389_LC_12_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1389_LC_12_28_0  (
            .in0(N__59137),
            .in1(N__53594),
            .in2(_gnd_net_),
            .in3(N__61999),
            .lcout(\c0.n33945 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1864_LC_12_28_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1864_LC_12_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1864_LC_12_28_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1864_LC_12_28_3  (
            .in0(N__53595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50521),
            .lcout(\c0.n18166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i185_LC_12_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i185_LC_12_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i185_LC_12_28_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_in_frame_0__i185_LC_12_28_6  (
            .in0(N__62241),
            .in1(N__73026),
            .in2(N__50649),
            .in3(N__80968),
            .lcout(\c0.data_in_frame_23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97789),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23806_4_lut_LC_13_6_0 .C_ON=1'b0;
    defparam \quad_counter0.i23806_4_lut_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23806_4_lut_LC_13_6_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter0.i23806_4_lut_LC_13_6_0  (
            .in0(N__50665),
            .in1(N__47840),
            .in2(N__47906),
            .in3(N__47721),
            .lcout(\quad_counter0.n1946 ),
            .ltout(\quad_counter0.n1946_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1354_3_lut_LC_13_6_1 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1354_3_lut_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1354_3_lut_LC_13_6_1 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \quad_counter0.mod_61_i1354_3_lut_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__47916),
            .in2(N__47715),
            .in3(N__47936),
            .lcout(\quad_counter0.n2016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1357_3_lut_LC_13_6_2 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1357_3_lut_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1357_3_lut_LC_13_6_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter0.mod_61_i1357_3_lut_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__60063),
            .in2(N__47709),
            .in3(N__53994),
            .lcout(\quad_counter0.n2019 ),
            .ltout(\quad_counter0.n2019_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23653_2_lut_LC_13_6_3 .C_ON=1'b0;
    defparam \quad_counter0.i23653_2_lut_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23653_2_lut_LC_13_6_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i23653_2_lut_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47712),
            .in3(N__60106),
            .lcout(\quad_counter0.n28371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1351_3_lut_LC_13_6_4 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1351_3_lut_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1351_3_lut_LC_13_6_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \quad_counter0.mod_61_i1351_3_lut_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__47850),
            .in2(N__47874),
            .in3(N__53998),
            .lcout(\quad_counter0.n2013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1353_3_lut_LC_13_6_7 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1353_3_lut_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1353_3_lut_LC_13_6_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter0.mod_61_i1353_3_lut_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__47902),
            .in2(N__54009),
            .in3(N__47886),
            .lcout(\quad_counter0.n2015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_2_lut_LC_13_7_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_2_lut_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_2_lut_LC_13_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_2_lut_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__60062),
            .in2(_gnd_net_),
            .in3(N__47700),
            .lcout(\quad_counter0.n1987 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\quad_counter0.n30215 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_3_lut_LC_13_7_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_3_lut_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_3_lut_LC_13_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_3_lut_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__54044),
            .in2(N__99331),
            .in3(N__47697),
            .lcout(\quad_counter0.n1986 ),
            .ltout(),
            .carryin(\quad_counter0.n30215 ),
            .carryout(\quad_counter0.n30216 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_4_lut_LC_13_7_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_4_lut_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_4_lut_LC_13_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_4_lut_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50714),
            .in3(N__47694),
            .lcout(\quad_counter0.n1985 ),
            .ltout(),
            .carryin(\quad_counter0.n30216 ),
            .carryout(\quad_counter0.n30217 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_5_lut_LC_13_7_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_5_lut_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_5_lut_LC_13_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_5_lut_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47937),
            .in3(N__47910),
            .lcout(\quad_counter0.n1984 ),
            .ltout(),
            .carryin(\quad_counter0.n30217 ),
            .carryout(\quad_counter0.n30218 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_6_lut_LC_13_7_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_6_lut_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_6_lut_LC_13_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_6_lut_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47907),
            .in3(N__47880),
            .lcout(\quad_counter0.n1983 ),
            .ltout(),
            .carryin(\quad_counter0.n30218 ),
            .carryout(\quad_counter0.n30219 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_7_lut_LC_13_7_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_7_lut_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_7_lut_LC_13_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_7_lut_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50672),
            .in3(N__47877),
            .lcout(\quad_counter0.n1982 ),
            .ltout(),
            .carryin(\quad_counter0.n30219 ),
            .carryout(\quad_counter0.n30220 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_8_lut_LC_13_7_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1348_8_lut_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_8_lut_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1348_8_lut_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47873),
            .in3(N__47844),
            .lcout(\quad_counter0.n1981 ),
            .ltout(),
            .carryin(\quad_counter0.n30220 ),
            .carryout(\quad_counter0.n30221 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1348_9_lut_LC_13_7_7 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1348_9_lut_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1348_9_lut_LC_13_7_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \quad_counter0.mod_61_add_1348_9_lut_LC_13_7_7  (
            .in0(N__99161),
            .in1(N__47841),
            .in2(N__54012),
            .in3(N__47829),
            .lcout(\quad_counter0.n2012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1178_LC_13_9_0 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1178_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1178_LC_13_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1178_LC_13_9_0  (
            .in0(N__47824),
            .in1(N__47967),
            .in2(N__47805),
            .in3(N__47727),
            .lcout(\quad_counter0.n35311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_2_lut_adj_1176_LC_13_9_1 .C_ON=1'b0;
    defparam \quad_counter0.i2_2_lut_adj_1176_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_2_lut_adj_1176_LC_13_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \quad_counter0.i2_2_lut_adj_1176_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__47767),
            .in2(_gnd_net_),
            .in3(N__47746),
            .lcout(\quad_counter0.n8_adj_4362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_2_lut_adj_1185_LC_13_9_2 .C_ON=1'b0;
    defparam \quad_counter0.i2_2_lut_adj_1185_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_2_lut_adj_1185_LC_13_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter0.i2_2_lut_adj_1185_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54295),
            .in3(N__54214),
            .lcout(),
            .ltout(\quad_counter0.n8_adj_4369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1187_LC_13_9_3 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1187_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1187_LC_13_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1187_LC_13_9_3  (
            .in0(N__54262),
            .in1(N__54238),
            .in2(N__48018),
            .in3(N__47961),
            .lcout(\quad_counter0.n34805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_3_lut_adj_1177_LC_13_9_4 .C_ON=1'b0;
    defparam \quad_counter0.i1_3_lut_adj_1177_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_3_lut_adj_1177_LC_13_9_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \quad_counter0.i1_3_lut_adj_1177_LC_13_9_4  (
            .in0(N__59914),
            .in1(N__48013),
            .in2(_gnd_net_),
            .in3(N__47989),
            .lcout(\quad_counter0.n7_adj_4363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_3_lut_adj_1186_LC_13_9_5 .C_ON=1'b0;
    defparam \quad_counter0.i1_3_lut_adj_1186_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_3_lut_adj_1186_LC_13_9_5 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \quad_counter0.i1_3_lut_adj_1186_LC_13_9_5  (
            .in0(N__59947),
            .in1(_gnd_net_),
            .in2(N__54346),
            .in3(N__54313),
            .lcout(\quad_counter0.n7_adj_4370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1211_LC_13_9_6 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1211_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1211_LC_13_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1211_LC_13_9_6  (
            .in0(N__63591),
            .in1(N__47946),
            .in2(N__63558),
            .in3(N__70578),
            .lcout(\quad_counter0.n34759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1191_LC_13_10_0 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1191_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1191_LC_13_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1191_LC_13_10_0  (
            .in0(N__54119),
            .in1(N__54973),
            .in2(N__54508),
            .in3(N__54850),
            .lcout(\quad_counter0.n27_adj_4374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_2_lut_adj_1184_LC_13_10_2 .C_ON=1'b0;
    defparam \quad_counter0.i1_2_lut_adj_1184_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_2_lut_adj_1184_LC_13_10_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i1_2_lut_adj_1184_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54541),
            .in3(N__54421),
            .lcout(),
            .ltout(\quad_counter0.n18_adj_4368_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i13_4_lut_adj_1188_LC_13_10_3 .C_ON=1'b0;
    defparam \quad_counter0.i13_4_lut_adj_1188_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i13_4_lut_adj_1188_LC_13_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i13_4_lut_adj_1188_LC_13_10_3  (
            .in0(N__54475),
            .in1(N__54362),
            .in2(N__47955),
            .in3(N__54949),
            .lcout(\quad_counter0.n30_adj_4371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i11_4_lut_adj_1189_LC_13_10_4 .C_ON=1'b0;
    defparam \quad_counter0.i11_4_lut_adj_1189_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i11_4_lut_adj_1189_LC_13_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i11_4_lut_adj_1189_LC_13_10_4  (
            .in0(N__47952),
            .in1(N__54898),
            .in2(N__54931),
            .in3(N__54874),
            .lcout(\quad_counter0.n28_adj_4372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_adj_1190_LC_13_10_5 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_adj_1190_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_adj_1190_LC_13_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i12_4_lut_adj_1190_LC_13_10_5  (
            .in0(N__54148),
            .in1(N__54451),
            .in2(N__54574),
            .in3(N__54391),
            .lcout(\quad_counter0.n29_adj_4373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_3_lut_adj_1210_LC_13_11_5 .C_ON=1'b0;
    defparam \quad_counter0.i1_3_lut_adj_1210_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_3_lut_adj_1210_LC_13_11_5 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \quad_counter0.i1_3_lut_adj_1210_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__63697),
            .in2(N__63663),
            .in3(N__63622),
            .lcout(\quad_counter0.n7_adj_4395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i6_4_lut_adj_1222_LC_13_12_1 .C_ON=1'b0;
    defparam \quad_counter0.i6_4_lut_adj_1222_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i6_4_lut_adj_1222_LC_13_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i6_4_lut_adj_1222_LC_13_12_1  (
            .in0(N__51137),
            .in1(N__51026),
            .in2(N__51340),
            .in3(N__51275),
            .lcout(\quad_counter0.n16_adj_4403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23615_2_lut_LC_13_12_4 .C_ON=1'b0;
    defparam \quad_counter0.i23615_2_lut_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23615_2_lut_LC_13_12_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23615_2_lut_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__59662),
            .in2(_gnd_net_),
            .in3(N__50933),
            .lcout(),
            .ltout(\quad_counter0.n28331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1221_LC_13_12_5 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1221_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1221_LC_13_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1221_LC_13_12_5  (
            .in0(N__51164),
            .in1(N__50906),
            .in2(N__48153),
            .in3(N__50879),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1223_LC_13_12_6 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1223_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1223_LC_13_12_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1223_LC_13_12_6  (
            .in0(N__50852),
            .in1(N__51110),
            .in2(N__48150),
            .in3(N__51191),
            .lcout(\quad_counter0.n14_adj_4404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_3_lut_LC_13_13_3 .C_ON=1'b0;
    defparam \quad_counter0.i8_3_lut_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_3_lut_LC_13_13_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter0.i8_3_lut_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__50999),
            .in2(N__51088),
            .in3(N__48147),
            .lcout(),
            .ltout(\quad_counter0.n18_adj_4405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i9_4_lut_adj_1224_LC_13_13_4 .C_ON=1'b0;
    defparam \quad_counter0.i9_4_lut_adj_1224_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i9_4_lut_adj_1224_LC_13_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i9_4_lut_adj_1224_LC_13_13_4  (
            .in0(N__48141),
            .in1(N__51053),
            .in2(N__48135),
            .in3(N__51305),
            .lcout(\quad_counter0.n2738 ),
            .ltout(\quad_counter0.n2738_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30722_1_lut_LC_13_13_5 .C_ON=1'b0;
    defparam \quad_counter0.i30722_1_lut_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30722_1_lut_LC_13_13_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30722_1_lut_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48063),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1737_LC_13_13_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1737_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1737_LC_13_13_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1737_LC_13_13_6  (
            .in0(N__91240),
            .in1(N__91071),
            .in2(_gnd_net_),
            .in3(N__93185),
            .lcout(\c0.n18011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1565_LC_13_14_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1565_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1565_LC_13_14_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.i3_4_lut_adj_1565_LC_13_14_0  (
            .in0(N__92679),
            .in1(N__84351),
            .in2(N__48344),
            .in3(N__55687),
            .lcout(\c0.n33170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1669_LC_13_14_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1669_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1669_LC_13_14_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1669_LC_13_14_1  (
            .in0(N__48359),
            .in1(N__48608),
            .in2(N__51747),
            .in3(N__48662),
            .lcout(\c0.n31012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1668_LC_13_14_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1668_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1668_LC_13_14_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1668_LC_13_14_2  (
            .in0(N__48661),
            .in1(N__48324),
            .in2(N__48612),
            .in3(N__48358),
            .lcout(\c0.data_out_frame_0__7__N_2569 ),
            .ltout(\c0.data_out_frame_0__7__N_2569_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i60_4_lut_LC_13_14_3 .C_ON=1'b0;
    defparam \c0.i60_4_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.i60_4_lut_LC_13_14_3 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \c0.i60_4_lut_LC_13_14_3  (
            .in0(N__48283),
            .in1(N__48207),
            .in2(N__48315),
            .in3(N__48308),
            .lcout(\c0.n58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30686_3_lut_4_lut_LC_13_14_4 .C_ON=1'b0;
    defparam \c0.i30686_3_lut_4_lut_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i30686_3_lut_4_lut_LC_13_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.i30686_3_lut_4_lut_LC_13_14_4  (
            .in0(N__48282),
            .in1(N__57492),
            .in2(N__55068),
            .in3(N__48239),
            .lcout(\c0.tx_transmit_N_3651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i286_2_lut_3_lut_4_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \c0.i286_2_lut_3_lut_4_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.i286_2_lut_3_lut_4_lut_LC_13_14_5 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \c0.i286_2_lut_3_lut_4_lut_LC_13_14_5  (
            .in0(N__57490),
            .in1(N__55063),
            .in2(N__48240),
            .in3(N__48281),
            .lcout(\c0.n688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30632_2_lut_3_lut_LC_13_14_6 .C_ON=1'b0;
    defparam \c0.i30632_2_lut_3_lut_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30632_2_lut_3_lut_LC_13_14_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \c0.i30632_2_lut_3_lut_LC_13_14_6  (
            .in0(N__55064),
            .in1(N__57491),
            .in2(_gnd_net_),
            .in3(N__48238),
            .lcout(\c0.n35938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1592_LC_13_14_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1592_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1592_LC_13_14_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i4_4_lut_adj_1592_LC_13_14_7  (
            .in0(N__84350),
            .in1(N__48201),
            .in2(N__55691),
            .in3(N__92678),
            .lcout(\c0.n35339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i114_4_lut_LC_13_15_0 .C_ON=1'b0;
    defparam \c0.i114_4_lut_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i114_4_lut_LC_13_15_0 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \c0.i114_4_lut_LC_13_15_0  (
            .in0(N__48408),
            .in1(N__48508),
            .in2(N__55371),
            .in3(N__51510),
            .lcout(\c0.n4_adj_4623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2045_LC_13_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2045_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2045_LC_13_15_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_2045_LC_13_15_1  (
            .in0(N__49111),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49268),
            .lcout(\c0.n14779 ),
            .ltout(\c0.n14779_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1951_LC_13_15_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1951_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1951_LC_13_15_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \c0.i1_4_lut_adj_1951_LC_13_15_2  (
            .in0(N__48557),
            .in1(N__48599),
            .in2(N__48627),
            .in3(N__48401),
            .lcout(\c0.n78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_403_Select_2_i6_3_lut_4_lut_LC_13_15_3 .C_ON=1'b0;
    defparam \c0.select_403_Select_2_i6_3_lut_4_lut_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_403_Select_2_i6_3_lut_4_lut_LC_13_15_3 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.select_403_Select_2_i6_3_lut_4_lut_LC_13_15_3  (
            .in0(N__51509),
            .in1(N__65363),
            .in2(N__92617),
            .in3(N__51694),
            .lcout(\c0.n6_adj_4617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1769_LC_13_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1769_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1769_LC_13_15_4 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1769_LC_13_15_4  (
            .in0(N__49270),
            .in1(N__49160),
            .in2(N__51861),
            .in3(N__49115),
            .lcout(\c0.n3315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23018_2_lut_3_lut_LC_13_15_5 .C_ON=1'b0;
    defparam \c0.i23018_2_lut_3_lut_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i23018_2_lut_3_lut_LC_13_15_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.i23018_2_lut_3_lut_LC_13_15_5  (
            .in0(N__48402),
            .in1(_gnd_net_),
            .in2(N__49121),
            .in3(N__49269),
            .lcout(\c0.n18115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23002_3_lut_4_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \c0.i23002_3_lut_4_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.i23002_3_lut_4_lut_LC_13_15_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.i23002_3_lut_4_lut_LC_13_15_6  (
            .in0(N__48600),
            .in1(N__48680),
            .in2(N__48561),
            .in3(N__48507),
            .lcout(\c0.n18045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i124_3_lut_4_lut_LC_13_15_7 .C_ON=1'b0;
    defparam \c0.i124_3_lut_4_lut_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i124_3_lut_4_lut_LC_13_15_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i124_3_lut_4_lut_LC_13_15_7  (
            .in0(N__49116),
            .in1(N__48473),
            .in2(N__48436),
            .in3(N__49271),
            .lcout(\c0.n118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1571_LC_13_16_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1571_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1571_LC_13_16_1 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1571_LC_13_16_1  (
            .in0(N__49094),
            .in1(N__48400),
            .in2(N__49173),
            .in3(N__49274),
            .lcout(\c0.n18100 ),
            .ltout(\c0.n18100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1676_LC_13_16_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1676_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1676_LC_13_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1676_LC_13_16_2  (
            .in0(N__48660),
            .in1(N__51858),
            .in2(N__48363),
            .in3(N__48360),
            .lcout(\c0.n63_adj_4633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1383_LC_13_16_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1383_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1383_LC_13_16_3 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1383_LC_13_16_3  (
            .in0(N__49093),
            .in1(N__51693),
            .in2(N__71271),
            .in3(N__49273),
            .lcout(\c0.n4_adj_4537 ),
            .ltout(\c0.n4_adj_4537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1947_LC_13_16_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1947_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1947_LC_13_16_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1947_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48765),
            .in3(N__51859),
            .lcout(),
            .ltout(\c0.n18020_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1508_LC_13_16_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1508_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1508_LC_13_16_5 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \c0.i2_4_lut_adj_1508_LC_13_16_5  (
            .in0(N__51370),
            .in1(N__92613),
            .in2(N__48762),
            .in3(N__48669),
            .lcout(),
            .ltout(\c0.n35757_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1509_LC_13_16_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1509_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1509_LC_13_16_6 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \c0.i1_4_lut_adj_1509_LC_13_16_6  (
            .in0(N__92614),
            .in1(N__55235),
            .in2(N__48759),
            .in3(N__48756),
            .lcout(),
            .ltout(\c0.n47_adj_4611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_13_16_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_13_16_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i0_LC_13_16_7 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_13_16_7  (
            .in0(N__51905),
            .in1(N__48720),
            .in2(N__48732),
            .in3(N__51559),
            .lcout(\c0.FRAME_MATCHER_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97594),
            .ce(),
            .sr(N__96914));
    defparam \c0.i1_4_lut_adj_1510_LC_13_17_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1510_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1510_LC_13_17_1 .LUT_INIT=16'b1111111110100010;
    LogicCell40 \c0.i1_4_lut_adj_1510_LC_13_17_1  (
            .in0(N__51521),
            .in1(N__65364),
            .in2(N__92615),
            .in3(N__48729),
            .lcout(\c0.n4_adj_4612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23419_2_lut_3_lut_LC_13_17_2 .C_ON=1'b0;
    defparam \c0.i23419_2_lut_3_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i23419_2_lut_3_lut_LC_13_17_2 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \c0.i23419_2_lut_3_lut_LC_13_17_2  (
            .in0(N__49070),
            .in1(_gnd_net_),
            .in2(N__49167),
            .in3(N__49275),
            .lcout(\c0.data_out_frame_29_7_N_1483_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_13_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_13_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i26_LC_13_17_4  (
            .in0(N__75325),
            .in1(N__57838),
            .in2(_gnd_net_),
            .in3(N__48703),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97603),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1946_LC_13_17_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1946_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1946_LC_13_17_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i2_3_lut_adj_1946_LC_13_17_5  (
            .in0(N__49276),
            .in1(N__48681),
            .in2(_gnd_net_),
            .in3(N__49071),
            .lcout(\c0.n30862 ),
            .ltout(\c0.n30862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1378_LC_13_17_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1378_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1378_LC_13_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1378_LC_13_17_6  (
            .in0(N__48663),
            .in1(N__51857),
            .in2(N__48636),
            .in3(N__51560),
            .lcout(\c0.n72 ),
            .ltout(\c0.n72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1538_LC_13_17_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1538_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1538_LC_13_17_7 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1538_LC_13_17_7  (
            .in0(N__49277),
            .in1(N__49156),
            .in2(N__49125),
            .in3(N__49072),
            .lcout(\c0.data_out_frame_0__7__N_2570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1965_LC_13_18_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1965_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1965_LC_13_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1965_LC_13_18_0  (
            .in0(N__48838),
            .in1(N__48796),
            .in2(_gnd_net_),
            .in3(N__52052),
            .lcout(),
            .ltout(\c0.n18675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1981_LC_13_18_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1981_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1981_LC_13_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1981_LC_13_18_1  (
            .in0(N__61341),
            .in1(N__49284),
            .in2(N__48978),
            .in3(N__48936),
            .lcout(\c0.n5_adj_4545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1991_LC_13_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1991_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1991_LC_13_18_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1991_LC_13_18_2  (
            .in0(N__57641),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48834),
            .lcout(\c0.n33347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1992_LC_13_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1992_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1992_LC_13_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1992_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__77210),
            .in2(_gnd_net_),
            .in3(N__64827),
            .lcout(\c0.n18667 ),
            .ltout(\c0.n18667_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1993_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1993_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1993_LC_13_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1993_LC_13_18_4  (
            .in0(N__51995),
            .in1(N__49379),
            .in2(N__48930),
            .in3(N__48917),
            .lcout(\c0.n18319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_13_18_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i1_LC_13_18_5  (
            .in0(N__81245),
            .in1(N__83914),
            .in2(N__48849),
            .in3(N__80808),
            .lcout(\c0.data_in_frame_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97615),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30379_4_lut_LC_13_18_7 .C_ON=1'b0;
    defparam \c0.i30379_4_lut_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30379_4_lut_LC_13_18_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i30379_4_lut_LC_13_18_7  (
            .in0(N__68079),
            .in1(N__52268),
            .in2(N__48801),
            .in3(N__61214),
            .lcout(\c0.n35806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1975_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1975_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1975_LC_13_19_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1975_LC_13_19_0  (
            .in0(N__72417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49320),
            .lcout(\c0.n33288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1366_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1366_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1366_LC_13_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1366_LC_13_19_1  (
            .in0(N__57668),
            .in1(N__72416),
            .in2(N__49938),
            .in3(N__52683),
            .lcout(\c0.n33326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1998_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1998_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1998_LC_13_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1998_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__49440),
            .in2(_gnd_net_),
            .in3(N__76142),
            .lcout(\c0.n18354 ),
            .ltout(\c0.n18354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1973_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1973_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1973_LC_13_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1973_LC_13_19_3  (
            .in0(N__49380),
            .in1(N__49364),
            .in2(N__49350),
            .in3(N__61226),
            .lcout(),
            .ltout(\c0.n29_adj_4767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1974_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1974_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1974_LC_13_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1974_LC_13_19_4  (
            .in0(N__49347),
            .in1(N__49335),
            .in2(N__49323),
            .in3(N__52005),
            .lcout(\c0.n33830 ),
            .ltout(\c0.n33830_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1961_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1961_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1961_LC_13_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1961_LC_13_19_5  (
            .in0(N__52214),
            .in1(N__49314),
            .in2(N__49287),
            .in3(N__64711),
            .lcout(\c0.data_out_frame_0__7__N_2580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1368_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1368_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1368_LC_13_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1368_LC_13_19_6  (
            .in0(N__49936),
            .in1(N__52261),
            .in2(_gnd_net_),
            .in3(N__52291),
            .lcout(\c0.n6_adj_4535 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_13_20_0 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_13_20_0  (
            .in0(N__65148),
            .in1(N__55623),
            .in2(_gnd_net_),
            .in3(N__55494),
            .lcout(\c0.rx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97645),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_13_20_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i17_LC_13_20_1  (
            .in0(N__80397),
            .in1(N__83911),
            .in2(N__52269),
            .in3(N__80955),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97645),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i64_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i64_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i64_LC_13_20_2 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_in_frame_0__i64_LC_13_20_2  (
            .in0(N__83910),
            .in1(N__49581),
            .in2(N__62178),
            .in3(N__80112),
            .lcout(\c0.data_in_frame_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97645),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_13_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_13_20_3  (
            .in0(N__49544),
            .in1(N__49500),
            .in2(_gnd_net_),
            .in3(N__49687),
            .lcout(),
            .ltout(\c0.n8_adj_4555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1851_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1851_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1851_LC_13_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1851_LC_13_20_4  (
            .in0(N__49655),
            .in1(N__49620),
            .in2(N__49596),
            .in3(N__49593),
            .lcout(\c0.n33441 ),
            .ltout(\c0.n33441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1836_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1836_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1836_LC_13_20_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1836_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49584),
            .in3(N__50197),
            .lcout(\c0.n6_adj_4733 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1395_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1395_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1395_LC_13_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1395_LC_13_20_6  (
            .in0(N__49580),
            .in1(N__49564),
            .in2(_gnd_net_),
            .in3(N__49711),
            .lcout(\c0.n33698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i63_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i63_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i63_LC_13_20_7 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i63_LC_13_20_7  (
            .in0(N__73518),
            .in1(N__62130),
            .in2(N__49548),
            .in3(N__83912),
            .lcout(\c0.data_in_frame_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97645),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1837_LC_13_21_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1837_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1837_LC_13_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1837_LC_13_21_0  (
            .in0(N__52622),
            .in1(N__49530),
            .in2(N__49911),
            .in3(N__49524),
            .lcout(\c0.n32302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i80_LC_13_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i80_LC_13_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i80_LC_13_21_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i80_LC_13_21_1  (
            .in0(N__58205),
            .in1(N__87259),
            .in2(N__80082),
            .in3(N__49499),
            .lcout(\c0.data_in_frame_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97659),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1858_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1858_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1858_LC_13_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1858_LC_13_21_2  (
            .in0(N__49498),
            .in1(N__49894),
            .in2(N__49484),
            .in3(N__49463),
            .lcout(\c0.n10_adj_4736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1890_LC_13_21_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1890_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1890_LC_13_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1890_LC_13_21_3  (
            .in0(N__49895),
            .in1(N__49958),
            .in2(N__49797),
            .in3(N__49944),
            .lcout(\c0.n18438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i35_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i35_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i35_LC_13_21_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i35_LC_13_21_5  (
            .in0(N__83863),
            .in1(N__73817),
            .in2(N__80640),
            .in3(N__49937),
            .lcout(\c0.data_in_frame_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97659),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i115_LC_13_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i115_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i115_LC_13_21_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i115_LC_13_21_6  (
            .in0(N__49910),
            .in1(N__80592),
            .in2(N__58365),
            .in3(N__89771),
            .lcout(\c0.data_in_frame_14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97659),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i65_LC_13_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i65_LC_13_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i65_LC_13_21_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i65_LC_13_21_7  (
            .in0(N__58204),
            .in1(N__80954),
            .in2(N__49899),
            .in3(N__81244),
            .lcout(\c0.data_in_frame_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97659),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1896_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1896_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1896_LC_13_22_0 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i5_3_lut_adj_1896_LC_13_22_0  (
            .in0(N__49879),
            .in1(N__49695),
            .in2(N__49823),
            .in3(_gnd_net_),
            .lcout(\c0.n33874 ),
            .ltout(\c0.n33874_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1401_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1401_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1401_LC_13_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1401_LC_13_22_1  (
            .in0(N__49860),
            .in1(N__50137),
            .in2(N__49827),
            .in3(N__52349),
            .lcout(\c0.n33422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1962_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1962_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1962_LC_13_22_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1962_LC_13_22_2  (
            .in0(N__49816),
            .in1(N__55399),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n5_adj_4742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1982_LC_13_22_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1982_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1982_LC_13_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1982_LC_13_22_3  (
            .in0(N__52218),
            .in1(N__52401),
            .in2(N__58710),
            .in3(N__49781),
            .lcout(\c0.n18705 ),
            .ltout(\c0.n18705_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1895_LC_13_22_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1895_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1895_LC_13_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1895_LC_13_22_4  (
            .in0(N__49743),
            .in1(N__55400),
            .in2(N__49719),
            .in3(N__49716),
            .lcout(\c0.n10_adj_4743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1899_LC_13_22_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1899_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1899_LC_13_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1899_LC_13_22_5  (
            .in0(N__50097),
            .in1(N__50166),
            .in2(N__52695),
            .in3(N__50138),
            .lcout(\c0.n10_adj_4744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1429_LC_13_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1429_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1429_LC_13_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1429_LC_13_22_6  (
            .in0(N__52350),
            .in1(N__50139),
            .in2(_gnd_net_),
            .in3(N__50096),
            .lcout(\c0.n18290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i98_LC_13_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i98_LC_13_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i98_LC_13_22_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i98_LC_13_22_7  (
            .in0(N__58321),
            .in1(N__73781),
            .in2(N__52626),
            .in3(N__75320),
            .lcout(\c0.data_in_frame_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1868_LC_13_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1868_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1868_LC_13_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1868_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__53023),
            .in2(_gnd_net_),
            .in3(N__53099),
            .lcout(\c0.n19064 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1835_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1835_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1835_LC_13_23_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1835_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__50081),
            .in2(_gnd_net_),
            .in3(N__55729),
            .lcout(\c0.n18373 ),
            .ltout(\c0.n18373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1843_LC_13_23_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1843_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1843_LC_13_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1843_LC_13_23_2  (
            .in0(N__68514),
            .in1(N__50036),
            .in2(N__49995),
            .in3(N__49992),
            .lcout(\c0.n33610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3286_2_lut_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.i3286_2_lut_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3286_2_lut_LC_13_23_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3286_2_lut_LC_13_23_3  (
            .in0(N__53098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55986),
            .lcout(\c0.n5965 ),
            .ltout(\c0.n5965_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1842_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1842_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1842_LC_13_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1842_LC_13_23_4  (
            .in0(N__49986),
            .in1(N__51623),
            .in2(N__49980),
            .in3(N__50469),
            .lcout(\c0.n33526 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i143_LC_13_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i143_LC_13_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i143_LC_13_23_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i143_LC_13_23_5  (
            .in0(N__73596),
            .in1(N__72902),
            .in2(N__49977),
            .in3(N__87296),
            .lcout(\c0.data_in_frame_17_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97690),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i84_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i84_LC_13_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i84_LC_13_23_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i84_LC_13_23_6  (
            .in0(N__58381),
            .in1(N__78981),
            .in2(N__80409),
            .in3(N__50297),
            .lcout(\c0.data_in_frame_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97690),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i151_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i151_LC_13_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i151_LC_13_23_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i151_LC_13_23_7  (
            .in0(N__73597),
            .in1(N__72903),
            .in2(N__50580),
            .in3(N__80385),
            .lcout(\c0.data_in_frame_18_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97690),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1787_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1787_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1787_LC_13_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1787_LC_13_24_0  (
            .in0(N__50337),
            .in1(N__53054),
            .in2(N__50283),
            .in3(N__53174),
            .lcout(\c0.n12_adj_4712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i100_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i100_LC_13_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i100_LC_13_24_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i100_LC_13_24_1  (
            .in0(N__78915),
            .in1(N__73878),
            .in2(N__58438),
            .in3(N__50338),
            .lcout(\c0.data_in_frame_12_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i228_LC_13_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i228_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i228_LC_13_24_2 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i228_LC_13_24_2  (
            .in0(N__79838),
            .in1(N__78916),
            .in2(N__73929),
            .in3(N__56165),
            .lcout(\c0.data_in_frame_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i33_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i33_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i33_LC_13_24_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i33_LC_13_24_3  (
            .in0(N__80969),
            .in1(N__73879),
            .in2(N__83975),
            .in3(N__52426),
            .lcout(\c0.data_in_frame_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1776_LC_13_24_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1776_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1776_LC_13_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1776_LC_13_24_4  (
            .in0(N__50268),
            .in1(N__52721),
            .in2(N__50259),
            .in3(N__50217),
            .lcout(\c0.n18971 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i129_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i129_LC_13_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i129_LC_13_24_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i129_LC_13_24_5  (
            .in0(N__81213),
            .in1(N__73007),
            .in2(N__80979),
            .in3(N__56372),
            .lcout(\c0.data_in_frame_16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i97_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i97_LC_13_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i97_LC_13_24_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i97_LC_13_24_7  (
            .in0(N__80970),
            .in1(N__73880),
            .in2(N__58439),
            .in3(N__50190),
            .lcout(\c0.data_in_frame_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97707),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_4_lut_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.i4_2_lut_4_lut_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_4_lut_LC_13_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_2_lut_4_lut_LC_13_25_0  (
            .in0(N__58956),
            .in1(N__59346),
            .in2(N__50438),
            .in3(N__53360),
            .lcout(\c0.n18_adj_4563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1516_LC_13_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1516_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1516_LC_13_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1516_LC_13_25_1  (
            .in0(N__59347),
            .in1(N__50434),
            .in2(_gnd_net_),
            .in3(N__58957),
            .lcout(\c0.n33994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i157_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i157_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i157_LC_13_25_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i157_LC_13_25_2  (
            .in0(N__84142),
            .in1(N__78166),
            .in2(N__50439),
            .in3(N__72975),
            .lcout(\c0.data_in_frame_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1504_LC_13_25_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1504_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1504_LC_13_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1504_LC_13_25_3  (
            .in0(N__59307),
            .in1(N__53405),
            .in2(N__50394),
            .in3(N__56414),
            .lcout(\c0.n14_adj_4578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1902_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1902_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1902_LC_13_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1902_LC_13_25_4  (
            .in0(N__50430),
            .in1(N__62324),
            .in2(_gnd_net_),
            .in3(N__50417),
            .lcout(\c0.n33551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1503_LC_13_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1503_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1503_LC_13_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1503_LC_13_25_5  (
            .in0(N__50389),
            .in1(N__74315),
            .in2(_gnd_net_),
            .in3(N__53404),
            .lcout(\c0.n6215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i159_LC_13_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i159_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i159_LC_13_25_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i159_LC_13_25_6  (
            .in0(N__73634),
            .in1(N__59348),
            .in2(N__73006),
            .in3(N__78167),
            .lcout(\c0.data_in_frame_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i213_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i213_LC_13_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i213_LC_13_26_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i213_LC_13_26_2  (
            .in0(N__69044),
            .in1(N__84232),
            .in2(N__80427),
            .in3(N__79880),
            .lcout(\c0.data_in_frame_26_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97742),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1617_LC_13_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1617_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1617_LC_13_26_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1617_LC_13_26_3  (
            .in0(N__50523),
            .in1(N__50529),
            .in2(N__65559),
            .in3(N__50483),
            .lcout(\c0.n32433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1849_LC_13_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1849_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1849_LC_13_26_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1849_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__53237),
            .in2(_gnd_net_),
            .in3(N__50342),
            .lcout(\c0.n33545 ),
            .ltout(\c0.n33545_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_13_26_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_13_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_13_26_5  (
            .in0(N__59121),
            .in1(N__50482),
            .in2(N__50619),
            .in3(N__52757),
            .lcout(),
            .ltout(\c0.n35505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1488_LC_13_26_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1488_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1488_LC_13_26_6 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \c0.i2_3_lut_adj_1488_LC_13_26_6  (
            .in0(N__50578),
            .in1(N__59091),
            .in2(N__50616),
            .in3(_gnd_net_),
            .lcout(\c0.n33653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1908_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1908_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1908_LC_13_26_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1908_LC_13_26_7  (
            .in0(N__69034),
            .in1(N__53636),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n33350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1892_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1892_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1892_LC_13_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1892_LC_13_27_1  (
            .in0(_gnd_net_),
            .in1(N__50608),
            .in2(_gnd_net_),
            .in3(N__53706),
            .lcout(),
            .ltout(\c0.n33852_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1496_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1496_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1496_LC_13_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1496_LC_13_27_2  (
            .in0(N__53154),
            .in1(N__50579),
            .in2(N__50544),
            .in3(N__50540),
            .lcout(\c0.n10_adj_4575 ),
            .ltout(\c0.n10_adj_4575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1618_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1618_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1618_LC_13_27_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1618_LC_13_27_3  (
            .in0(N__53846),
            .in1(N__50522),
            .in2(N__50487),
            .in3(N__50484),
            .lcout(\c0.n32390 ),
            .ltout(\c0.n32390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_13_27_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_13_27_4  (
            .in0(N__59362),
            .in1(N__59308),
            .in2(N__50451),
            .in3(N__56610),
            .lcout(\c0.n20_adj_4627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i183_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i183_LC_13_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i183_LC_13_27_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i183_LC_13_27_5  (
            .in0(N__73038),
            .in1(N__89752),
            .in2(N__74123),
            .in3(N__73636),
            .lcout(\c0.data_in_frame_22_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i167_LC_13_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i167_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i167_LC_13_27_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i167_LC_13_27_7  (
            .in0(N__73037),
            .in1(N__73928),
            .in2(N__53787),
            .in3(N__73635),
            .lcout(\c0.data_in_frame_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97760),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i150_LC_13_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i150_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i150_LC_13_28_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i150_LC_13_28_0  (
            .in0(N__80336),
            .in1(N__72984),
            .in2(N__53549),
            .in3(N__75087),
            .lcout(\c0.data_in_frame_18_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i166_LC_13_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i166_LC_13_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i166_LC_13_28_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i166_LC_13_28_2  (
            .in0(N__73927),
            .in1(N__75086),
            .in2(N__56492),
            .in3(N__72983),
            .lcout(\c0.data_in_frame_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97776),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1677_LC_13_28_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1677_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1677_LC_13_28_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1677_LC_13_28_5  (
            .in0(N__65679),
            .in1(N__50645),
            .in2(N__74119),
            .in3(N__53726),
            .lcout(\c0.n33939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i219_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i219_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i219_LC_13_28_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i219_LC_13_28_6  (
            .in0(N__78321),
            .in1(N__80709),
            .in2(N__79881),
            .in3(N__68807),
            .lcout(\c0.data_in_frame_27_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97776),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_2_lut_LC_14_5_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_2_lut_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_2_lut_LC_14_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_2_lut_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60108),
            .in3(N__50634),
            .lcout(\quad_counter0.n2087 ),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\quad_counter0.n30222 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_3_lut_LC_14_5_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_3_lut_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_3_lut_LC_14_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_3_lut_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__99150),
            .in2(N__50796),
            .in3(N__50631),
            .lcout(\quad_counter0.n2086 ),
            .ltout(),
            .carryin(\quad_counter0.n30222 ),
            .carryout(\quad_counter0.n30223 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_4_lut_LC_14_5_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_4_lut_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_4_lut_LC_14_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_4_lut_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53967),
            .in3(N__50628),
            .lcout(\quad_counter0.n2085 ),
            .ltout(),
            .carryin(\quad_counter0.n30223 ),
            .carryout(\quad_counter0.n30224 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_5_lut_LC_14_5_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_5_lut_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_5_lut_LC_14_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_5_lut_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53679),
            .in3(N__50625),
            .lcout(\quad_counter0.n2084 ),
            .ltout(),
            .carryin(\quad_counter0.n30224 ),
            .carryout(\quad_counter0.n30225 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_6_lut_LC_14_5_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_6_lut_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_6_lut_LC_14_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_6_lut_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53942),
            .in3(N__50622),
            .lcout(\quad_counter0.n2083 ),
            .ltout(),
            .carryin(\quad_counter0.n30225 ),
            .carryout(\quad_counter0.n30226 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_7_lut_LC_14_5_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_7_lut_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_7_lut_LC_14_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_7_lut_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54080),
            .in3(N__50748),
            .lcout(\quad_counter0.n2082 ),
            .ltout(),
            .carryin(\quad_counter0.n30226 ),
            .carryout(\quad_counter0.n30227 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_8_lut_LC_14_5_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_8_lut_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_8_lut_LC_14_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_8_lut_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54102),
            .in3(N__50745),
            .lcout(\quad_counter0.n2081 ),
            .ltout(),
            .carryin(\quad_counter0.n30227 ),
            .carryout(\quad_counter0.n30228 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_9_lut_LC_14_5_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1415_9_lut_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_9_lut_LC_14_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.mod_61_add_1415_9_lut_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__99151),
            .in2(N__50820),
            .in3(N__50742),
            .lcout(\quad_counter0.n2080 ),
            .ltout(),
            .carryin(\quad_counter0.n30228 ),
            .carryout(\quad_counter0.n30229 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1415_10_lut_LC_14_6_0 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1415_10_lut_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1415_10_lut_LC_14_6_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \quad_counter0.mod_61_add_1415_10_lut_LC_14_6_0  (
            .in0(N__99149),
            .in1(N__50832),
            .in2(N__53907),
            .in3(N__50739),
            .lcout(\quad_counter0.n2111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1425_3_lut_LC_14_6_1 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1425_3_lut_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1425_3_lut_LC_14_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.mod_61_i1425_3_lut_LC_14_6_1  (
            .in0(N__60107),
            .in1(N__50736),
            .in2(_gnd_net_),
            .in3(N__53900),
            .lcout(\quad_counter0.n2119 ),
            .ltout(\quad_counter0.n2119_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_3_lut_adj_1198_LC_14_6_2 .C_ON=1'b0;
    defparam \quad_counter0.i1_3_lut_adj_1198_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_3_lut_adj_1198_LC_14_6_2 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \quad_counter0.i1_3_lut_adj_1198_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__60145),
            .in2(N__50730),
            .in3(N__56879),
            .lcout(\quad_counter0.n7_adj_4381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1355_3_lut_LC_14_6_3 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1355_3_lut_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1355_3_lut_LC_14_6_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \quad_counter0.mod_61_i1355_3_lut_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__50727),
            .in2(N__50721),
            .in3(N__54011),
            .lcout(\quad_counter0.n2017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1418_3_lut_LC_14_7_1 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1418_3_lut_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1418_3_lut_LC_14_7_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \quad_counter0.mod_61_i1418_3_lut_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__50691),
            .in2(N__50819),
            .in3(N__53904),
            .lcout(\quad_counter0.n2112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1352_3_lut_LC_14_7_2 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1352_3_lut_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1352_3_lut_LC_14_7_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \quad_counter0.mod_61_i1352_3_lut_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__50682),
            .in2(N__50676),
            .in3(N__54005),
            .lcout(\quad_counter0.n2014 ),
            .ltout(\quad_counter0.n2014_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1196_LC_14_7_3 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1196_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1196_LC_14_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1196_LC_14_7_3  (
            .in0(N__53966),
            .in1(N__53677),
            .in2(N__50841),
            .in3(N__50838),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4378_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_4_lut_LC_14_7_4 .C_ON=1'b0;
    defparam \quad_counter0.i2_4_lut_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_4_lut_LC_14_7_4 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \quad_counter0.i2_4_lut_LC_14_7_4  (
            .in0(N__50831),
            .in1(N__50812),
            .in2(N__50799),
            .in3(N__50769),
            .lcout(\quad_counter0.n2045 ),
            .ltout(\quad_counter0.n2045_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1424_3_lut_LC_14_7_5 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1424_3_lut_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1424_3_lut_LC_14_7_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter0.mod_61_i1424_3_lut_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__50795),
            .in2(N__50781),
            .in3(N__50778),
            .lcout(\quad_counter0.n2118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_2_lut_LC_14_7_6 .C_ON=1'b0;
    defparam \quad_counter0.i3_2_lut_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_2_lut_LC_14_7_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter0.i3_2_lut_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53941),
            .in3(N__54073),
            .lcout(\quad_counter0.n9_adj_4379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12_4_lut_LC_14_9_0 .C_ON=1'b0;
    defparam \quad_counter0.i12_4_lut_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12_4_lut_LC_14_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i12_4_lut_LC_14_9_0  (
            .in0(N__54585),
            .in1(N__54408),
            .in2(N__54711),
            .in3(N__54438),
            .lcout(),
            .ltout(\quad_counter0.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i15_4_lut_LC_14_9_1 .C_ON=1'b0;
    defparam \quad_counter0.i15_4_lut_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i15_4_lut_LC_14_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i15_4_lut_LC_14_9_1  (
            .in0(N__54552),
            .in1(N__54993),
            .in2(N__50763),
            .in3(N__50754),
            .lcout(\quad_counter0.n33_adj_4346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23575_2_lut_LC_14_9_2 .C_ON=1'b0;
    defparam \quad_counter0.i23575_2_lut_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23575_2_lut_LC_14_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23575_2_lut_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__59983),
            .in2(_gnd_net_),
            .in3(N__57154),
            .lcout(),
            .ltout(\quad_counter0.n28291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_LC_14_9_3 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_LC_14_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_LC_14_9_3  (
            .in0(N__57094),
            .in1(N__57127),
            .in2(N__50760),
            .in3(N__57316),
            .lcout(),
            .ltout(\quad_counter0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_LC_14_9_4 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_LC_14_9_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \quad_counter0.i3_4_lut_LC_14_9_4  (
            .in0(N__54519),
            .in1(N__57355),
            .in2(N__50757),
            .in3(N__57388),
            .lcout(\quad_counter0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30610_4_lut_LC_14_9_5 .C_ON=1'b0;
    defparam \quad_counter0.i30610_4_lut_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30610_4_lut_LC_14_9_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i30610_4_lut_LC_14_9_5  (
            .in0(N__57356),
            .in1(N__59984),
            .in2(N__57161),
            .in3(N__50979),
            .lcout(\quad_counter0.n35976 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30712_1_lut_LC_14_9_6 .C_ON=1'b0;
    defparam \quad_counter0.i30712_1_lut_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30712_1_lut_LC_14_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30712_1_lut_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54769),
            .lcout(\quad_counter0.n36139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1212_LC_14_10_0 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1212_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1212_LC_14_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1212_LC_14_10_0  (
            .in0(N__64020),
            .in1(N__64050),
            .in2(N__64113),
            .in3(N__50985),
            .lcout(\quad_counter0.n12_adj_4396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_LC_14_10_5 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_LC_14_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i5_4_lut_LC_14_10_5  (
            .in0(N__57128),
            .in1(N__57095),
            .in2(N__57392),
            .in3(N__57317),
            .lcout(\quad_counter0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i16_4_lut_adj_1192_LC_14_10_6 .C_ON=1'b0;
    defparam \quad_counter0.i16_4_lut_adj_1192_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i16_4_lut_adj_1192_LC_14_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i16_4_lut_adj_1192_LC_14_10_6  (
            .in0(N__50973),
            .in1(N__50967),
            .in2(N__50961),
            .in3(N__50952),
            .lcout(\quad_counter0.n3431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_2_lut_LC_14_11_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_2_lut_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_2_lut_LC_14_11_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1817_2_lut_LC_14_11_0  (
            .in0(N__60204),
            .in1(N__60203),
            .in2(N__54694),
            .in3(N__50922),
            .lcout(\quad_counter0.n2719 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\quad_counter0.n30285 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_3_lut_LC_14_11_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_3_lut_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_3_lut_LC_14_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_3_lut_LC_14_11_1  (
            .in0(N__60234),
            .in1(N__60233),
            .in2(N__54649),
            .in3(N__50895),
            .lcout(\quad_counter0.n2718 ),
            .ltout(),
            .carryin(\quad_counter0.n30285 ),
            .carryout(\quad_counter0.n30286 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_4_lut_LC_14_11_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_4_lut_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_4_lut_LC_14_11_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1817_4_lut_LC_14_11_2  (
            .in0(N__60753),
            .in1(N__60752),
            .in2(N__54695),
            .in3(N__50868),
            .lcout(\quad_counter0.n2717 ),
            .ltout(),
            .carryin(\quad_counter0.n30286 ),
            .carryout(\quad_counter0.n30287 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_5_lut_LC_14_11_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_5_lut_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_5_lut_LC_14_11_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1817_5_lut_LC_14_11_3  (
            .in0(N__60726),
            .in1(N__60725),
            .in2(N__54698),
            .in3(N__51207),
            .lcout(\quad_counter0.n2716 ),
            .ltout(),
            .carryin(\quad_counter0.n30287 ),
            .carryout(\quad_counter0.n30288 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_6_lut_LC_14_11_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_6_lut_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_6_lut_LC_14_11_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1817_6_lut_LC_14_11_4  (
            .in0(N__60696),
            .in1(N__60695),
            .in2(N__54696),
            .in3(N__51180),
            .lcout(\quad_counter0.n2715 ),
            .ltout(),
            .carryin(\quad_counter0.n30288 ),
            .carryout(\quad_counter0.n30289 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_7_lut_LC_14_11_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_7_lut_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_7_lut_LC_14_11_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1817_7_lut_LC_14_11_5  (
            .in0(N__60669),
            .in1(N__60668),
            .in2(N__54699),
            .in3(N__51153),
            .lcout(\quad_counter0.n2714 ),
            .ltout(),
            .carryin(\quad_counter0.n30289 ),
            .carryout(\quad_counter0.n30290 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_8_lut_LC_14_11_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_8_lut_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_8_lut_LC_14_11_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1817_8_lut_LC_14_11_6  (
            .in0(N__60639),
            .in1(N__60638),
            .in2(N__54697),
            .in3(N__51126),
            .lcout(\quad_counter0.n2713 ),
            .ltout(),
            .carryin(\quad_counter0.n30290 ),
            .carryout(\quad_counter0.n30291 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_9_lut_LC_14_11_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_9_lut_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_9_lut_LC_14_11_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_9_lut_LC_14_11_7  (
            .in0(N__60612),
            .in1(N__60611),
            .in2(N__54650),
            .in3(N__51099),
            .lcout(\quad_counter0.n2712 ),
            .ltout(),
            .carryin(\quad_counter0.n30291 ),
            .carryout(\quad_counter0.n30292 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_10_lut_LC_14_12_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_10_lut_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_10_lut_LC_14_12_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_10_lut_LC_14_12_0  (
            .in0(N__60579),
            .in1(N__60578),
            .in2(N__54651),
            .in3(N__51069),
            .lcout(\quad_counter0.n2711 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\quad_counter0.n30293 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_11_lut_LC_14_12_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_11_lut_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_11_lut_LC_14_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_11_lut_LC_14_12_1  (
            .in0(N__60549),
            .in1(N__60548),
            .in2(N__54655),
            .in3(N__51042),
            .lcout(\quad_counter0.n2710 ),
            .ltout(),
            .carryin(\quad_counter0.n30293 ),
            .carryout(\quad_counter0.n30294 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_12_lut_LC_14_12_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_12_lut_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_12_lut_LC_14_12_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_12_lut_LC_14_12_2  (
            .in0(N__60912),
            .in1(N__60911),
            .in2(N__54652),
            .in3(N__51015),
            .lcout(\quad_counter0.n2709 ),
            .ltout(),
            .carryin(\quad_counter0.n30294 ),
            .carryout(\quad_counter0.n30295 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_13_lut_LC_14_12_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_13_lut_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_13_lut_LC_14_12_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_13_lut_LC_14_12_3  (
            .in0(N__60882),
            .in1(N__60881),
            .in2(N__54656),
            .in3(N__50988),
            .lcout(\quad_counter0.n2708 ),
            .ltout(),
            .carryin(\quad_counter0.n30295 ),
            .carryout(\quad_counter0.n30296 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_14_lut_LC_14_12_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_14_lut_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_14_lut_LC_14_12_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_14_lut_LC_14_12_4  (
            .in0(N__60855),
            .in1(N__60854),
            .in2(N__54653),
            .in3(N__51321),
            .lcout(\quad_counter0.n2707 ),
            .ltout(),
            .carryin(\quad_counter0.n30296 ),
            .carryout(\quad_counter0.n30297 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_15_lut_LC_14_12_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1817_15_lut_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_15_lut_LC_14_12_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_15_lut_LC_14_12_5  (
            .in0(N__60828),
            .in1(N__60827),
            .in2(N__54657),
            .in3(N__51294),
            .lcout(\quad_counter0.n2706 ),
            .ltout(),
            .carryin(\quad_counter0.n30297 ),
            .carryout(\quad_counter0.n30298 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1817_16_lut_LC_14_12_6 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1817_16_lut_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1817_16_lut_LC_14_12_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1817_16_lut_LC_14_12_6  (
            .in0(N__60797),
            .in1(N__60798),
            .in2(N__54654),
            .in3(N__51291),
            .lcout(\quad_counter0.n2705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i6_4_lut_LC_14_13_1 .C_ON=1'b0;
    defparam \quad_counter0.i6_4_lut_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i6_4_lut_LC_14_13_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i6_4_lut_LC_14_13_1  (
            .in0(N__64175),
            .in1(N__64080),
            .in2(N__64146),
            .in3(N__51264),
            .lcout(\quad_counter0.n2441 ),
            .ltout(\quad_counter0.n2441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30726_1_lut_LC_14_13_2 .C_ON=1'b0;
    defparam \quad_counter0.i30726_1_lut_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30726_1_lut_LC_14_13_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30726_1_lut_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51255),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_14_13_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_14_13_3 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_14_13_3  (
            .in0(N__58617),
            .in1(N__51248),
            .in2(N__71147),
            .in3(N__71676),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97562),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1427__i0_LC_14_14_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i0_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i0_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i0_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__95913),
            .in2(N__51230),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\c0.n30202 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i1_LC_14_14_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i1_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i1_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i1_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__90193),
            .in2(_gnd_net_),
            .in3(N__51213),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n30202 ),
            .carryout(\c0.n30203 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i2_LC_14_14_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i2_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i2_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i2_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__89949),
            .in2(_gnd_net_),
            .in3(N__51210),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(\c0.n30203 ),
            .carryout(\c0.n30204 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i3_LC_14_14_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i3_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i3_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i3_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__95734),
            .in2(_gnd_net_),
            .in3(N__51456),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(\c0.n30204 ),
            .carryout(\c0.n30205 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i4_LC_14_14_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i4_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i4_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i4_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__90693),
            .in2(_gnd_net_),
            .in3(N__51453),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(\c0.n30205 ),
            .carryout(\c0.n30206 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i5_LC_14_14_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i5_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i5_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i5_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__71124),
            .in2(_gnd_net_),
            .in3(N__51450),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(\c0.n30206 ),
            .carryout(\c0.n30207 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i6_LC_14_14_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter_1427__i6_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i6_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i6_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__55080),
            .in2(_gnd_net_),
            .in3(N__51447),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(\c0.n30207 ),
            .carryout(\c0.n30208 ),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.byte_transmit_counter_1427__i7_LC_14_14_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1427__i7_LC_14_14_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter_1427__i7_LC_14_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter_1427__i7_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__55092),
            .in2(_gnd_net_),
            .in3(N__51444),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97570),
            .ce(N__51441),
            .sr(N__51414));
    defparam \c0.i2_3_lut_4_lut_adj_1345_LC_14_15_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1345_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1345_LC_14_15_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1345_LC_14_15_0  (
            .in0(N__51551),
            .in1(N__51856),
            .in2(N__51906),
            .in3(N__51586),
            .lcout(data_out_frame_29__7__N_1482),
            .ltout(data_out_frame_29__7__N_1482_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__2__5451_LC_14_15_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__2__5451_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__2__5451_LC_14_15_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_9__2__5451_LC_14_15_1  (
            .in0(N__57477),
            .in1(N__85161),
            .in2(N__51399),
            .in3(N__83331),
            .lcout(data_out_frame_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97579),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_LC_14_15_3.C_ON=1'b0;
    defparam i24_3_lut_4_lut_LC_14_15_3.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_LC_14_15_3.LUT_INIT=16'b1111001011010000;
    LogicCell40 i24_3_lut_4_lut_LC_14_15_3 (
            .in0(N__95732),
            .in1(N__90692),
            .in2(N__71523),
            .in3(N__55278),
            .lcout(n10_adj_4805),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1734_LC_14_15_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1734_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1734_LC_14_15_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1734_LC_14_15_4  (
            .in0(N__91456),
            .in1(N__62071),
            .in2(N__91329),
            .in3(N__90493),
            .lcout(\c0.n17961 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__5__5448_LC_14_15_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__5__5448_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__5__5448_LC_14_15_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_9__5__5448_LC_14_15_5  (
            .in0(N__84422),
            .in1(N__85162),
            .in2(N__96642),
            .in3(N__67715),
            .lcout(data_out_frame_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__0__5429_LC_14_15_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__0__5429_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__0__5429_LC_14_15_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_12__0__5429_LC_14_15_6  (
            .in0(N__85160),
            .in1(N__84423),
            .in2(N__75885),
            .in3(N__55118),
            .lcout(data_out_frame_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1952_LC_14_15_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1952_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1952_LC_14_15_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1952_LC_14_15_7  (
            .in0(N__51855),
            .in1(N__51901),
            .in2(N__51590),
            .in3(N__51550),
            .lcout(\c0.data_out_frame_0__7__N_2571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30570_2_lut_LC_14_16_0 .C_ON=1'b0;
    defparam \c0.i30570_2_lut_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i30570_2_lut_LC_14_16_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i30570_2_lut_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__90206),
            .in2(_gnd_net_),
            .in3(N__51464),
            .lcout(\c0.n35963 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__2__5523_LC_14_16_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__2__5523_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__2__5523_LC_14_16_2 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \c0.data_out_frame_0__2__5523_LC_14_16_2  (
            .in0(N__51758),
            .in1(N__51745),
            .in2(N__51483),
            .in3(N__51707),
            .lcout(\c0.data_out_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97585),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30604_2_lut_LC_14_16_3 .C_ON=1'b0;
    defparam \c0.i30604_2_lut_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i30604_2_lut_LC_14_16_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i30604_2_lut_LC_14_16_3  (
            .in0(N__90207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51479),
            .lcout(),
            .ltout(\c0.n35960_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_14_16_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_14_16_4 .LUT_INIT=16'b1000100000110000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_14_16_4  (
            .in0(N__51983),
            .in1(N__90017),
            .in2(N__51471),
            .in3(N__96068),
            .lcout(),
            .ltout(\c0.n6_adj_4510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30406_4_lut_LC_14_16_5 .C_ON=1'b0;
    defparam \c0.i30406_4_lut_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30406_4_lut_LC_14_16_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.i30406_4_lut_LC_14_16_5  (
            .in0(N__90208),
            .in1(N__90018),
            .in2(N__51468),
            .in3(N__55305),
            .lcout(\c0.n35833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__3__5522_LC_14_16_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__3__5522_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__3__5522_LC_14_16_6 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \c0.data_out_frame_0__3__5522_LC_14_16_6  (
            .in0(N__51759),
            .in1(N__51746),
            .in2(N__51708),
            .in3(N__51465),
            .lcout(\c0.data_out_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97585),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__2__5483_LC_14_16_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__2__5483_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__2__5483_LC_14_16_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__2__5483_LC_14_16_7  (
            .in0(N__85146),
            .in1(N__84426),
            .in2(N__72207),
            .in3(N__51984),
            .lcout(data_out_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97585),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_14_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_14_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_14_17_0  (
            .in0(N__51965),
            .in1(N__51974),
            .in2(_gnd_net_),
            .in3(N__96067),
            .lcout(\c0.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__0__5477_LC_14_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__0__5477_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__0__5477_LC_14_17_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_6__0__5477_LC_14_17_1  (
            .in0(N__51975),
            .in1(N__84475),
            .in2(N__78048),
            .in3(N__85096),
            .lcout(data_out_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97595),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__0__5469_LC_14_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__0__5469_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__0__5469_LC_14_17_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_7__0__5469_LC_14_17_3  (
            .in0(N__85076),
            .in1(N__84476),
            .in2(N__86430),
            .in3(N__51966),
            .lcout(data_out_frame_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97595),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1335_LC_14_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1335_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1335_LC_14_17_5 .LUT_INIT=16'b1101110111111100;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1335_LC_14_17_5  (
            .in0(N__51957),
            .in1(N__51748),
            .in2(N__85178),
            .in3(N__51696),
            .lcout(),
            .ltout(\c0.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_2048_LC_14_17_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_2048_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_2048_LC_14_17_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \c0.i3_4_lut_adj_2048_LC_14_17_6  (
            .in0(N__51938),
            .in1(N__51900),
            .in2(N__51864),
            .in3(N__51860),
            .lcout(\c0.n19297 ),
            .ltout(\c0.n19297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_0__4__5521_LC_14_17_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_0__4__5521_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_0__4__5521_LC_14_17_7 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \c0.data_out_frame_0__4__5521_LC_14_17_7  (
            .in0(N__65168),
            .in1(N__51749),
            .in2(N__51711),
            .in3(N__51697),
            .lcout(\c0.data_out_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97595),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i113_LC_14_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i113_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i113_LC_14_18_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i113_LC_14_18_0  (
            .in0(N__58298),
            .in1(N__89735),
            .in2(N__51622),
            .in3(N__80922),
            .lcout(\c0.data_in_frame_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1367_LC_14_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1367_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1367_LC_14_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1367_LC_14_18_1  (
            .in0(N__77203),
            .in1(N__64826),
            .in2(_gnd_net_),
            .in3(N__83616),
            .lcout(\c0.n18663 ),
            .ltout(\c0.n18663_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1969_LC_14_18_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1969_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1969_LC_14_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1969_LC_14_18_2  (
            .in0(N__68072),
            .in1(N__64731),
            .in2(N__52224),
            .in3(N__58680),
            .lcout(),
            .ltout(\c0.n33397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1970_LC_14_18_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1970_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1970_LC_14_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1970_LC_14_18_3  (
            .in0(N__61210),
            .in1(N__57640),
            .in2(N__52221),
            .in3(N__52236),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_14_18_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i10_LC_14_18_4  (
            .in0(N__68073),
            .in1(N__75269),
            .in2(N__87299),
            .in3(N__83811),
            .lcout(data_in_frame_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1976_LC_14_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1976_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1976_LC_14_18_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1976_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__52433),
            .in2(_gnd_net_),
            .in3(N__83617),
            .lcout(\c0.n33604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_14_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_14_18_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i2_LC_14_18_6  (
            .in0(N__81243),
            .in1(N__83810),
            .in2(N__52065),
            .in3(N__75270),
            .lcout(\c0.data_in_frame_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i73_LC_14_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i73_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i73_LC_14_18_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i73_LC_14_18_7  (
            .in0(N__80921),
            .in1(N__58299),
            .in2(N__52192),
            .in3(N__87270),
            .lcout(\c0.data_in_frame_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_LC_14_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_3_lut_4_lut_LC_14_19_0  (
            .in0(N__52170),
            .in1(N__52121),
            .in2(N__52063),
            .in3(N__52011),
            .lcout(\c0.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_14_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_14_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_14_19_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i52_LC_14_19_1  (
            .in0(N__83808),
            .in1(N__78947),
            .in2(N__51999),
            .in3(N__89773),
            .lcout(\c0.data_in_frame_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1990_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1990_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1990_LC_14_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1990_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__57669),
            .in2(_gnd_net_),
            .in3(N__72418),
            .lcout(),
            .ltout(\c0.n33344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1994_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1994_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1994_LC_14_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1994_LC_14_19_3  (
            .in0(N__52434),
            .in1(N__52410),
            .in2(N__52404),
            .in3(N__52260),
            .lcout(),
            .ltout(\c0.n10_adj_4770_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1995_LC_14_19_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1995_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1995_LC_14_19_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_3_lut_adj_1995_LC_14_19_4  (
            .in0(N__52397),
            .in1(_gnd_net_),
            .in2(N__52362),
            .in3(N__52310),
            .lcout(\c0.n18314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_14_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_14_19_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i51_LC_14_19_5  (
            .in0(N__83807),
            .in1(N__80601),
            .in2(N__52314),
            .in3(N__89772),
            .lcout(\c0.data_in_frame_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i36_LC_14_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i36_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i36_LC_14_19_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i36_LC_14_19_6  (
            .in0(N__78946),
            .in1(N__73848),
            .in2(N__52295),
            .in3(N__83809),
            .lcout(\c0.data_in_frame_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1977_LC_14_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1977_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1977_LC_14_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1977_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__52287),
            .in2(_gnd_net_),
            .in3(N__52259),
            .lcout(\c0.n33692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_14_20_1 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_14_20_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.rx.i2_2_lut_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__65076),
            .in2(_gnd_net_),
            .in3(N__55801),
            .lcout(),
            .ltout(\c0.rx.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30689_4_lut_LC_14_20_2 .C_ON=1'b0;
    defparam \c0.rx.i30689_4_lut_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30689_4_lut_LC_14_20_2 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \c0.rx.i30689_4_lut_LC_14_20_2  (
            .in0(N__76991),
            .in1(N__65138),
            .in2(N__52230),
            .in3(N__55930),
            .lcout(n19327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30592_4_lut_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.rx.i30592_4_lut_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30592_4_lut_LC_14_20_3 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \c0.rx.i30592_4_lut_LC_14_20_3  (
            .in0(N__58533),
            .in1(N__65075),
            .in2(N__58566),
            .in3(N__55782),
            .lcout(),
            .ltout(\c0.rx.n35949_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_1326_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_1326_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_1326_LC_14_20_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \c0.rx.i1_4_lut_adj_1326_LC_14_20_4  (
            .in0(N__76990),
            .in1(N__65137),
            .in2(N__52227),
            .in3(N__55740),
            .lcout(n19940),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_107_i4_2_lut_LC_14_20_5 .C_ON=1'b0;
    defparam \c0.rx.equal_107_i4_2_lut_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_107_i4_2_lut_LC_14_20_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.equal_107_i4_2_lut_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__55436),
            .in2(_gnd_net_),
            .in3(N__55549),
            .lcout(n4_adj_4807),
            .ltout(n4_adj_4807_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_14_20_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_14_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_14_20_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_14_20_6  (
            .in0(N__75202),
            .in1(N__55931),
            .in2(N__52557),
            .in3(N__52554),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97629),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1353_LC_14_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1353_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1353_LC_14_20_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1353_LC_14_20_7  (
            .in0(N__58016),
            .in1(N__68581),
            .in2(N__57829),
            .in3(N__92837),
            .lcout(\c0.n33241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_14_21_0 .C_ON=1'b0;
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.equal_87_i9_2_lut_3_lut_LC_14_21_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.equal_87_i9_2_lut_3_lut_LC_14_21_0  (
            .in0(N__93202),
            .in1(N__91263),
            .in2(_gnd_net_),
            .in3(N__91111),
            .lcout(\c0.n9_adj_4631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1343_LC_14_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1343_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1343_LC_14_21_1 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1343_LC_14_21_1  (
            .in0(N__91470),
            .in1(N__91560),
            .in2(N__91371),
            .in3(N__91653),
            .lcout(\c0.n12_adj_4518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_14_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_14_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_14_21_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i43_LC_14_21_2  (
            .in0(N__80720),
            .in1(N__68304),
            .in2(N__78639),
            .in3(N__52509),
            .lcout(\c0.data_in_frame_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1407_LC_14_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1407_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1407_LC_14_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1407_LC_14_21_3  (
            .in0(N__52705),
            .in1(N__52947),
            .in2(_gnd_net_),
            .in3(N__52481),
            .lcout(\c0.n6_adj_4546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i111_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i111_LC_14_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i111_LC_14_21_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i111_LC_14_21_4  (
            .in0(N__73617),
            .in1(N__53097),
            .in2(N__78638),
            .in3(N__68590),
            .lcout(\c0.data_in_frame_13_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i123_LC_14_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i123_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i123_LC_14_21_5 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.data_in_frame_0__i123_LC_14_21_5  (
            .in0(N__52707),
            .in1(N__80721),
            .in2(N__62225),
            .in3(N__58206),
            .lcout(\c0.data_in_frame_15_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i105_LC_14_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i105_LC_14_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i105_LC_14_21_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i105_LC_14_21_6  (
            .in0(N__80956),
            .in1(N__68589),
            .in2(N__52955),
            .in3(N__78628),
            .lcout(\c0.data_in_frame_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97646),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1897_LC_14_21_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1897_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1897_LC_14_21_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1897_LC_14_21_7  (
            .in0(N__52706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52948),
            .lcout(\c0.n33321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_14_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_14_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_14_22_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i32_LC_14_22_1  (
            .in0(N__78335),
            .in1(N__83812),
            .in2(N__52682),
            .in3(N__80123),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i127_LC_14_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i127_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i127_LC_14_22_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i127_LC_14_22_2  (
            .in0(N__58318),
            .in1(N__62173),
            .in2(N__52651),
            .in3(N__73621),
            .lcout(\c0.data_in_frame_15_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i124_LC_14_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i124_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i124_LC_14_22_3 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.data_in_frame_0__i124_LC_14_22_3  (
            .in0(N__78982),
            .in1(N__58319),
            .in2(N__56068),
            .in3(N__62177),
            .lcout(\c0.data_in_frame_15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1411_LC_14_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1411_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1411_LC_14_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1411_LC_14_22_4  (
            .in0(N__53017),
            .in1(N__53121),
            .in2(_gnd_net_),
            .in3(N__53096),
            .lcout(\c0.n33591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i128_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i128_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i128_LC_14_22_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_in_frame_0__i128_LC_14_22_5  (
            .in0(N__62172),
            .in1(N__80122),
            .in2(N__53129),
            .in3(N__58320),
            .lcout(\c0.data_in_frame_15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i110_LC_14_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i110_LC_14_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i110_LC_14_22_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i110_LC_14_22_6  (
            .in0(N__68594),
            .in1(N__75053),
            .in2(N__53027),
            .in3(N__78575),
            .lcout(\c0.data_in_frame_13_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1861_LC_14_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1861_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1861_LC_14_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1861_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__56253),
            .in2(_gnd_net_),
            .in3(N__52621),
            .lcout(\c0.n33843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1876_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1876_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1876_LC_14_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1876_LC_14_23_0  (
            .in0(N__52831),
            .in1(N__56227),
            .in2(N__52992),
            .in3(N__53561),
            .lcout(\c0.n31_adj_4740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2052_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2052_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_2052_LC_14_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_2052_LC_14_23_1  (
            .in0(N__53125),
            .in1(N__53022),
            .in2(N__53103),
            .in3(N__52841),
            .lcout(),
            .ltout(\c0.n31480_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1802_LC_14_23_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1802_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1802_LC_14_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1802_LC_14_23_2  (
            .in0(N__53070),
            .in1(N__53503),
            .in2(N__53058),
            .in3(N__56670),
            .lcout(\c0.n32357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1893_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1893_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1893_LC_14_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1893_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__53044),
            .in2(_gnd_net_),
            .in3(N__52830),
            .lcout(\c0.n18881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1797_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1797_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1797_LC_14_23_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1797_LC_14_23_4  (
            .in0(N__53021),
            .in1(N__52988),
            .in2(_gnd_net_),
            .in3(N__52977),
            .lcout(\c0.n33913 ),
            .ltout(\c0.n33913_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1799_LC_14_23_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1799_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1799_LC_14_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1799_LC_14_23_5  (
            .in0(N__52956),
            .in1(N__52932),
            .in2(N__52920),
            .in3(N__52917),
            .lcout(\c0.n16010 ),
            .ltout(\c0.n16010_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1796_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1796_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1796_LC_14_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1796_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__52911),
            .in2(N__52890),
            .in3(N__52887),
            .lcout(\c0.n32241 ),
            .ltout(\c0.n32241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1492_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1492_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1492_LC_14_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1492_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__52859),
            .in2(N__52845),
            .in3(N__52842),
            .lcout(\c0.n33827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1473_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1473_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1473_LC_14_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1473_LC_14_24_0  (
            .in0(N__53211),
            .in1(N__52833),
            .in2(N__52779),
            .in3(N__52756),
            .lcout(\c0.n33629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i101_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i101_LC_14_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i101_LC_14_24_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i101_LC_14_24_1  (
            .in0(N__84246),
            .in1(N__58426),
            .in2(N__53221),
            .in3(N__73847),
            .lcout(\c0.data_in_frame_12_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97691),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i229_LC_14_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i229_LC_14_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i229_LC_14_24_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i229_LC_14_24_2  (
            .in0(N__53274),
            .in1(N__84247),
            .in2(N__73910),
            .in3(N__79846),
            .lcout(\c0.data_in_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97691),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1911_LC_14_24_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1911_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1911_LC_14_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1911_LC_14_24_3  (
            .in0(N__68474),
            .in1(N__53273),
            .in2(N__58797),
            .in3(N__53262),
            .lcout(),
            .ltout(\c0.n12_adj_4748_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1913_LC_14_24_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1913_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1913_LC_14_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1913_LC_14_24_4  (
            .in0(N__79508),
            .in1(N__61631),
            .in2(N__53265),
            .in3(N__65640),
            .lcout(\c0.n34566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1530_LC_14_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1530_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1530_LC_14_24_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1530_LC_14_24_5  (
            .in0(N__66018),
            .in1(N__69083),
            .in2(_gnd_net_),
            .in3(N__68895),
            .lcout(\c0.n33517 ),
            .ltout(\c0.n33517_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1932_LC_14_24_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1932_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1932_LC_14_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1932_LC_14_24_6  (
            .in0(N__58821),
            .in1(N__59022),
            .in2(N__53256),
            .in3(N__68871),
            .lcout(\c0.n35633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1630_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1630_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1630_LC_14_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1630_LC_14_25_0  (
            .in0(N__56609),
            .in1(N__59280),
            .in2(N__73173),
            .in3(N__56178),
            .lcout(\c0.n33662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1852_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1852_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1852_LC_14_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1852_LC_14_25_1  (
            .in0(N__56516),
            .in1(N__56248),
            .in2(_gnd_net_),
            .in3(N__53253),
            .lcout(\c0.n33768 ),
            .ltout(\c0.n33768_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1854_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1854_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1854_LC_14_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1854_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__53207),
            .in2(N__53178),
            .in3(N__53175),
            .lcout(\c0.n6023 ),
            .ltout(\c0.n6023_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1500_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1500_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1500_LC_14_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1500_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__53710),
            .in2(N__53439),
            .in3(N__53432),
            .lcout(\c0.n33458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1514_LC_14_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1514_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1514_LC_14_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1514_LC_14_25_5  (
            .in0(N__56028),
            .in1(N__56608),
            .in2(_gnd_net_),
            .in3(N__79453),
            .lcout(\c0.n33889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1771_LC_14_25_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1771_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1771_LC_14_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1771_LC_14_25_6  (
            .in0(N__56568),
            .in1(N__53388),
            .in2(_gnd_net_),
            .in3(N__53379),
            .lcout(\c0.n32339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1773_LC_14_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1773_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1773_LC_14_25_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1773_LC_14_25_7  (
            .in0(N__56027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79452),
            .lcout(\c0.n33979 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1907_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1907_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1907_LC_14_26_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1907_LC_14_26_0  (
            .in0(N__73321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56192),
            .lcout(\c0.n32366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1795_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1795_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1795_LC_14_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1795_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__53363),
            .in2(_gnd_net_),
            .in3(N__56220),
            .lcout(\c0.n33966 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1499_LC_14_26_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1499_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1499_LC_14_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1499_LC_14_26_2  (
            .in0(N__56687),
            .in1(N__59224),
            .in2(N__56228),
            .in3(N__59177),
            .lcout(\c0.n33621 ),
            .ltout(\c0.n33621_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1786_LC_14_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1786_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1786_LC_14_26_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1786_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53367),
            .in3(N__53364),
            .lcout(),
            .ltout(\c0.n8_adj_4711_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1788_LC_14_26_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1788_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1788_LC_14_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1788_LC_14_26_4  (
            .in0(N__53319),
            .in1(N__53295),
            .in2(N__53286),
            .in3(N__53283),
            .lcout(\c0.n18578 ),
            .ltout(\c0.n18578_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1904_LC_14_26_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1904_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1904_LC_14_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1904_LC_14_26_5  (
            .in0(N__53817),
            .in1(N__59042),
            .in2(N__53652),
            .in3(N__53472),
            .lcout(),
            .ltout(\c0.n15_adj_4746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1905_LC_14_26_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1905_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1905_LC_14_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1905_LC_14_26_6  (
            .in0(N__74246),
            .in1(N__65584),
            .in2(N__53649),
            .in3(N__53646),
            .lcout(\c0.n32087 ),
            .ltout(\c0.n32087_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_14_26_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_14_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_14_26_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_14_26_7  (
            .in0(N__65942),
            .in1(N__73322),
            .in2(N__53640),
            .in3(N__65879),
            .lcout(\c0.n14_adj_4538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i187_LC_14_27_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i187_LC_14_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i187_LC_14_27_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i187_LC_14_27_1  (
            .in0(N__80680),
            .in1(N__62224),
            .in2(N__53764),
            .in3(N__73039),
            .lcout(\c0.data_in_frame_23_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97743),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i214_LC_14_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i214_LC_14_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i214_LC_14_27_2 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i214_LC_14_27_2  (
            .in0(N__75049),
            .in1(N__53637),
            .in2(N__80395),
            .in3(N__79843),
            .lcout(\c0.data_in_frame_26_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97743),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i206_LC_14_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i206_LC_14_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i206_LC_14_27_4 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i206_LC_14_27_4  (
            .in0(N__75048),
            .in1(N__65937),
            .in2(N__87301),
            .in3(N__79842),
            .lcout(\c0.data_in_frame_25_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97743),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1693_LC_14_27_5 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1693_LC_14_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1693_LC_14_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1693_LC_14_27_5  (
            .in0(N__65880),
            .in1(N__53621),
            .in2(N__53763),
            .in3(N__53471),
            .lcout(\c0.n38_adj_4701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1650_LC_14_27_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1650_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1650_LC_14_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1650_LC_14_27_6  (
            .in0(N__56717),
            .in1(N__53605),
            .in2(N__62447),
            .in3(N__53568),
            .lcout(\c0.n18559 ),
            .ltout(\c0.n18559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_4_lut_LC_14_27_7 .C_ON=1'b0;
    defparam \c0.i3_2_lut_4_lut_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_4_lut_LC_14_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_2_lut_4_lut_LC_14_27_7  (
            .in0(N__53535),
            .in1(N__53514),
            .in2(N__53475),
            .in3(N__53470),
            .lcout(\c0.n16_adj_4667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1634_LC_14_28_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1634_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1634_LC_14_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1634_LC_14_28_0  (
            .in0(N__74060),
            .in1(N__66401),
            .in2(N__53769),
            .in3(N__53826),
            .lcout(),
            .ltout(\c0.n15_adj_4664_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1635_LC_14_28_1 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1635_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1635_LC_14_28_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1635_LC_14_28_1  (
            .in0(N__53853),
            .in1(N__53832),
            .in2(N__53835),
            .in3(N__66371),
            .lcout(\c0.n16118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1647_LC_14_28_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1647_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1647_LC_14_28_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1647_LC_14_28_2  (
            .in0(N__56481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53738),
            .lcout(\c0.n33563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1633_LC_14_28_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1633_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1633_LC_14_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1633_LC_14_28_3  (
            .in0(N__69213),
            .in1(N__61740),
            .in2(_gnd_net_),
            .in3(N__74093),
            .lcout(\c0.n14_adj_4663 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1569_LC_14_28_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1569_LC_14_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1569_LC_14_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1569_LC_14_28_4  (
            .in0(N__53782),
            .in1(N__53812),
            .in2(N__56488),
            .in3(N__53825),
            .lcout(\c0.n33858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3725_2_lut_LC_14_28_5 .C_ON=1'b0;
    defparam \c0.i3725_2_lut_LC_14_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3725_2_lut_LC_14_28_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i3725_2_lut_LC_14_28_5  (
            .in0(N__53813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53783),
            .lcout(),
            .ltout(\c0.n6404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1636_LC_14_28_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1636_LC_14_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1636_LC_14_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1636_LC_14_28_6  (
            .in0(N__53765),
            .in1(N__53739),
            .in2(N__53730),
            .in3(N__53727),
            .lcout(\c0.n33638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i135_LC_14_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i135_LC_14_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i135_LC_14_28_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i135_LC_14_28_7  (
            .in0(N__81220),
            .in1(N__72985),
            .in2(N__53714),
            .in3(N__73622),
            .lcout(\c0.data_in_frame_16_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97761),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1422_3_lut_LC_15_6_0 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1422_3_lut_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1422_3_lut_LC_15_6_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter0.mod_61_i1422_3_lut_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(N__53678),
            .in2(N__53905),
            .in3(N__53658),
            .lcout(\quad_counter0.n2116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1419_3_lut_LC_15_6_2 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1419_3_lut_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1419_3_lut_LC_15_6_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \quad_counter0.mod_61_i1419_3_lut_LC_15_6_2  (
            .in0(N__54108),
            .in1(N__54098),
            .in2(N__53906),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n2113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1420_3_lut_LC_15_6_3 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1420_3_lut_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1420_3_lut_LC_15_6_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \quad_counter0.mod_61_i1420_3_lut_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__53892),
            .in2(N__54084),
            .in3(N__54057),
            .lcout(\quad_counter0.n2114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1356_3_lut_LC_15_6_4 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1356_3_lut_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1356_3_lut_LC_15_6_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter0.mod_61_i1356_3_lut_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(N__54051),
            .in2(N__54027),
            .in3(N__54010),
            .lcout(\quad_counter0.n2018 ),
            .ltout(\quad_counter0.n2018_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1423_3_lut_LC_15_6_5 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1423_3_lut_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1423_3_lut_LC_15_6_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \quad_counter0.mod_61_i1423_3_lut_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(N__53952),
            .in2(N__53946),
            .in3(N__53891),
            .lcout(\quad_counter0.n2117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_i1421_3_lut_LC_15_6_7 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_i1421_3_lut_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_i1421_3_lut_LC_15_6_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter0.mod_61_i1421_3_lut_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(N__53943),
            .in2(N__53916),
            .in3(N__53896),
            .lcout(\quad_counter0.n2115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_2_lut_adj_1197_LC_15_7_0 .C_ON=1'b0;
    defparam \quad_counter0.i2_2_lut_adj_1197_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_2_lut_adj_1197_LC_15_7_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter0.i2_2_lut_adj_1197_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56865),
            .in3(N__56797),
            .lcout(),
            .ltout(\quad_counter0.n8_adj_4380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1199_LC_15_7_1 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1199_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1199_LC_15_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1199_LC_15_7_1  (
            .in0(N__56818),
            .in1(N__56839),
            .in2(N__53865),
            .in3(N__53862),
            .lcout(),
            .ltout(\quad_counter0.n35542_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i3_4_lut_adj_1200_LC_15_7_2 .C_ON=1'b0;
    defparam \quad_counter0.i3_4_lut_adj_1200_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i3_4_lut_adj_1200_LC_15_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i3_4_lut_adj_1200_LC_15_7_2  (
            .in0(N__56770),
            .in1(N__56746),
            .in2(N__53856),
            .in3(N__57053),
            .lcout(\quad_counter0.n2144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_2_lut_LC_15_9_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_2_lut_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_2_lut_LC_15_9_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2353_2_lut_LC_15_9_0  (
            .in0(N__59949),
            .in1(N__59948),
            .in2(N__54196),
            .in3(N__54351),
            .lcout(\quad_counter0.n3519 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\quad_counter0.n30425 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_3_lut_LC_15_9_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_3_lut_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_3_lut_LC_15_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_3_lut_LC_15_9_1  (
            .in0(N__54348),
            .in1(N__54347),
            .in2(N__54821),
            .in3(N__54324),
            .lcout(\quad_counter0.n3518 ),
            .ltout(),
            .carryin(\quad_counter0.n30425 ),
            .carryout(\quad_counter0.n30426 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_4_lut_LC_15_9_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_4_lut_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_4_lut_LC_15_9_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2353_4_lut_LC_15_9_2  (
            .in0(N__54321),
            .in1(N__54320),
            .in2(N__54197),
            .in3(N__54300),
            .lcout(\quad_counter0.n3517 ),
            .ltout(),
            .carryin(\quad_counter0.n30426 ),
            .carryout(\quad_counter0.n30427 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_5_lut_LC_15_9_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_5_lut_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_5_lut_LC_15_9_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2353_5_lut_LC_15_9_3  (
            .in0(N__54297),
            .in1(N__54296),
            .in2(N__54200),
            .in3(N__54273),
            .lcout(\quad_counter0.n3516 ),
            .ltout(),
            .carryin(\quad_counter0.n30427 ),
            .carryout(\quad_counter0.n30428 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_6_lut_LC_15_9_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_6_lut_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_6_lut_LC_15_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2353_6_lut_LC_15_9_4  (
            .in0(N__54270),
            .in1(N__54269),
            .in2(N__54198),
            .in3(N__54249),
            .lcout(\quad_counter0.n3515 ),
            .ltout(),
            .carryin(\quad_counter0.n30428 ),
            .carryout(\quad_counter0.n30429 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_7_lut_LC_15_9_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_7_lut_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_7_lut_LC_15_9_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2353_7_lut_LC_15_9_5  (
            .in0(N__54246),
            .in1(N__54245),
            .in2(N__54201),
            .in3(N__54225),
            .lcout(\quad_counter0.n3514 ),
            .ltout(),
            .carryin(\quad_counter0.n30429 ),
            .carryout(\quad_counter0.n30430 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_8_lut_LC_15_9_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_8_lut_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_8_lut_LC_15_9_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_2353_8_lut_LC_15_9_6  (
            .in0(N__54222),
            .in1(N__54221),
            .in2(N__54199),
            .in3(N__54159),
            .lcout(\quad_counter0.n3513 ),
            .ltout(),
            .carryin(\quad_counter0.n30430 ),
            .carryout(\quad_counter0.n30431 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_9_lut_LC_15_9_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_9_lut_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_9_lut_LC_15_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_9_lut_LC_15_9_7  (
            .in0(N__54156),
            .in1(N__54155),
            .in2(N__54822),
            .in3(N__54135),
            .lcout(\quad_counter0.n3512 ),
            .ltout(),
            .carryin(\quad_counter0.n30431 ),
            .carryout(\quad_counter0.n30432 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_10_lut_LC_15_10_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_10_lut_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_10_lut_LC_15_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_10_lut_LC_15_10_0  (
            .in0(N__54132),
            .in1(N__54131),
            .in2(N__54823),
            .in3(N__54579),
            .lcout(\quad_counter0.n3511 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\quad_counter0.n30433 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_11_lut_LC_15_10_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_11_lut_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_11_lut_LC_15_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_11_lut_LC_15_10_1  (
            .in0(N__54576),
            .in1(N__54575),
            .in2(N__54827),
            .in3(N__54546),
            .lcout(\quad_counter0.n3510 ),
            .ltout(),
            .carryin(\quad_counter0.n30433 ),
            .carryout(\quad_counter0.n30434 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_12_lut_LC_15_10_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_12_lut_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_12_lut_LC_15_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_12_lut_LC_15_10_2  (
            .in0(N__54543),
            .in1(N__54542),
            .in2(N__54824),
            .in3(N__54513),
            .lcout(\quad_counter0.n3509 ),
            .ltout(),
            .carryin(\quad_counter0.n30434 ),
            .carryout(\quad_counter0.n30435 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_13_lut_LC_15_10_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_13_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_13_lut_LC_15_10_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_13_lut_LC_15_10_3  (
            .in0(N__54510),
            .in1(N__54509),
            .in2(N__54828),
            .in3(N__54486),
            .lcout(\quad_counter0.n3508 ),
            .ltout(),
            .carryin(\quad_counter0.n30435 ),
            .carryout(\quad_counter0.n30436 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_14_lut_LC_15_10_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_14_lut_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_14_lut_LC_15_10_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_14_lut_LC_15_10_4  (
            .in0(N__54483),
            .in1(N__54482),
            .in2(N__54825),
            .in3(N__54462),
            .lcout(\quad_counter0.n3507 ),
            .ltout(),
            .carryin(\quad_counter0.n30436 ),
            .carryout(\quad_counter0.n30437 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_15_lut_LC_15_10_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_15_lut_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_15_lut_LC_15_10_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_15_lut_LC_15_10_5  (
            .in0(N__54459),
            .in1(N__54458),
            .in2(N__54829),
            .in3(N__54432),
            .lcout(\quad_counter0.n3506 ),
            .ltout(),
            .carryin(\quad_counter0.n30437 ),
            .carryout(\quad_counter0.n30438 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_16_lut_LC_15_10_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_16_lut_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_16_lut_LC_15_10_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_16_lut_LC_15_10_6  (
            .in0(N__54429),
            .in1(N__54428),
            .in2(N__54826),
            .in3(N__54402),
            .lcout(\quad_counter0.n3505 ),
            .ltout(),
            .carryin(\quad_counter0.n30438 ),
            .carryout(\quad_counter0.n30439 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_17_lut_LC_15_10_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_17_lut_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_17_lut_LC_15_10_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_17_lut_LC_15_10_7  (
            .in0(N__54399),
            .in1(N__54398),
            .in2(N__54830),
            .in3(N__54378),
            .lcout(\quad_counter0.n3504 ),
            .ltout(),
            .carryin(\quad_counter0.n30439 ),
            .carryout(\quad_counter0.n30440 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_18_lut_LC_15_11_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_18_lut_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_18_lut_LC_15_11_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_18_lut_LC_15_11_0  (
            .in0(N__54375),
            .in1(N__54374),
            .in2(N__54831),
            .in3(N__54984),
            .lcout(\quad_counter0.n3503 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\quad_counter0.n30441 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_19_lut_LC_15_11_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_19_lut_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_19_lut_LC_15_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_19_lut_LC_15_11_1  (
            .in0(N__54981),
            .in1(N__54980),
            .in2(N__54835),
            .in3(N__54960),
            .lcout(\quad_counter0.n3502 ),
            .ltout(),
            .carryin(\quad_counter0.n30441 ),
            .carryout(\quad_counter0.n30442 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_20_lut_LC_15_11_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_20_lut_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_20_lut_LC_15_11_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_20_lut_LC_15_11_2  (
            .in0(N__54957),
            .in1(N__54956),
            .in2(N__54832),
            .in3(N__54936),
            .lcout(\quad_counter0.n3501 ),
            .ltout(),
            .carryin(\quad_counter0.n30442 ),
            .carryout(\quad_counter0.n30443 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_21_lut_LC_15_11_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_21_lut_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_21_lut_LC_15_11_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_21_lut_LC_15_11_3  (
            .in0(N__54933),
            .in1(N__54932),
            .in2(N__54836),
            .in3(N__54909),
            .lcout(\quad_counter0.n3500 ),
            .ltout(),
            .carryin(\quad_counter0.n30443 ),
            .carryout(\quad_counter0.n30444 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_22_lut_LC_15_11_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_22_lut_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_22_lut_LC_15_11_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_22_lut_LC_15_11_4  (
            .in0(N__54906),
            .in1(N__54905),
            .in2(N__54833),
            .in3(N__54885),
            .lcout(\quad_counter0.n3499 ),
            .ltout(),
            .carryin(\quad_counter0.n30444 ),
            .carryout(\quad_counter0.n30445 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_23_lut_LC_15_11_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_2353_23_lut_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_23_lut_LC_15_11_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_23_lut_LC_15_11_5  (
            .in0(N__54882),
            .in1(N__54881),
            .in2(N__54837),
            .in3(N__54861),
            .lcout(\quad_counter0.n3498 ),
            .ltout(),
            .carryin(\quad_counter0.n30445 ),
            .carryout(\quad_counter0.n30446 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_2353_24_lut_LC_15_11_6 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_2353_24_lut_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_2353_24_lut_LC_15_11_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_2353_24_lut_LC_15_11_6  (
            .in0(N__54857),
            .in1(N__54858),
            .in2(N__54834),
            .in3(N__54714),
            .lcout(\quad_counter0.n3497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30723_1_lut_LC_15_11_7 .C_ON=1'b0;
    defparam \quad_counter0.i30723_1_lut_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30723_1_lut_LC_15_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30723_1_lut_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54648),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_adj_1220_LC_15_12_0 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_adj_1220_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_adj_1220_LC_15_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_adj_1220_LC_15_12_0  (
            .in0(N__60610),
            .in1(N__60826),
            .in2(N__57273),
            .in3(N__57291),
            .lcout(\quad_counter0.n2639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__0__5421_LC_15_13_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__0__5421_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__0__5421_LC_15_13_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_13__0__5421_LC_15_13_6  (
            .in0(N__85164),
            .in1(N__55104),
            .in2(N__101334),
            .in3(N__84497),
            .lcout(data_out_frame_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97557),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_15_14_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_15_14_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_15_14_2  (
            .in0(N__71113),
            .in1(N__71688),
            .in2(N__55139),
            .in3(N__57444),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_15_14_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_15_14_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_15_14_3  (
            .in0(N__55119),
            .in1(N__95989),
            .in2(_gnd_net_),
            .in3(N__55103),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1601_LC_15_14_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1601_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1601_LC_15_14_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1601_LC_15_14_4  (
            .in0(N__71112),
            .in1(N__55091),
            .in2(_gnd_net_),
            .in3(N__55079),
            .lcout(\c0.n4_adj_4646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_15_14_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_15_14_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_15_14_6  (
            .in0(N__71114),
            .in1(N__71689),
            .in2(N__55049),
            .in3(N__57438),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30656_4_lut_LC_15_15_0 .C_ON=1'b0;
    defparam \c0.i30656_4_lut_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \c0.i30656_4_lut_LC_15_15_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.i30656_4_lut_LC_15_15_0  (
            .in0(N__90192),
            .in1(N__57450),
            .in2(N__90074),
            .in3(N__89166),
            .lcout(),
            .ltout(n36084_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2063_LC_15_15_1.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2063_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2063_LC_15_15_1.LUT_INIT=16'b1011100010101010;
    LogicCell40 i24_3_lut_4_lut_adj_2063_LC_15_15_1 (
            .in0(N__55170),
            .in1(N__90694),
            .in2(N__55026),
            .in3(N__95733),
            .lcout(n10_adj_4804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_15_15_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_15_15_2 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_15_15_2  (
            .in0(N__55007),
            .in1(N__71690),
            .in2(N__71146),
            .in3(N__55257),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97571),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__1__5436_LC_15_15_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__1__5436_LC_15_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__1__5436_LC_15_15_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_11__1__5436_LC_15_15_3  (
            .in0(N__84424),
            .in1(N__85070),
            .in2(N__77877),
            .in3(N__55188),
            .lcout(data_out_frame_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97571),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__1__5444_LC_15_15_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__1__5444_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__1__5444_LC_15_15_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_10__1__5444_LC_15_15_4  (
            .in0(N__85069),
            .in1(N__84425),
            .in2(N__67815),
            .in3(N__55197),
            .lcout(data_out_frame_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97571),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_15_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_15_5 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_15_5  (
            .in0(N__55196),
            .in1(N__95912),
            .in2(N__90314),
            .in3(N__55187),
            .lcout(\c0.n36209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7838_2_lut_LC_15_16_0 .C_ON=1'b0;
    defparam \c0.i7838_2_lut_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7838_2_lut_LC_15_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i7838_2_lut_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__85028),
            .in2(_gnd_net_),
            .in3(N__84352),
            .lcout(\c0.n12483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__0__5453_LC_15_16_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__0__5453_LC_15_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__0__5453_LC_15_16_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_9__0__5453_LC_15_16_2  (
            .in0(N__55164),
            .in1(N__84353),
            .in2(N__85632),
            .in3(N__85029),
            .lcout(data_out_frame_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30408_4_lut_LC_15_16_3 .C_ON=1'b0;
    defparam \c0.i30408_4_lut_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i30408_4_lut_LC_15_16_3 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.i30408_4_lut_LC_15_16_3  (
            .in0(N__93888),
            .in1(N__55179),
            .in2(N__90885),
            .in3(N__90724),
            .lcout(n35835),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1586_LC_15_16_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1586_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1586_LC_15_16_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_1586_LC_15_16_4  (
            .in0(N__90498),
            .in1(N__91321),
            .in2(_gnd_net_),
            .in3(N__91452),
            .lcout(\c0.n17959 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36197_bdd_4_lut_LC_15_16_6 .C_ON=1'b0;
    defparam \c0.n36197_bdd_4_lut_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.n36197_bdd_4_lut_LC_15_16_6 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n36197_bdd_4_lut_LC_15_16_6  (
            .in0(N__55163),
            .in1(N__61047),
            .in2(N__90379),
            .in3(N__57587),
            .lcout(),
            .ltout(\c0.n36200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30659_4_lut_LC_15_16_7 .C_ON=1'b0;
    defparam \c0.i30659_4_lut_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30659_4_lut_LC_15_16_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.i30659_4_lut_LC_15_16_7  (
            .in0(N__55155),
            .in1(N__90005),
            .in2(N__55146),
            .in3(N__90335),
            .lcout(n36088),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__2__5475_LC_15_17_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__2__5475_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__2__5475_LC_15_17_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_6__2__5475_LC_15_17_0  (
            .in0(N__55314),
            .in1(N__84627),
            .in2(N__85165),
            .in3(N__85929),
            .lcout(data_out_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_15_17_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_15_17_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_15_17_1  (
            .in0(N__61095),
            .in1(N__55313),
            .in2(_gnd_net_),
            .in3(N__96015),
            .lcout(\c0.n5_adj_4511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__1__5460_LC_15_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__1__5460_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__1__5460_LC_15_17_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_8__1__5460_LC_15_17_3  (
            .in0(N__84626),
            .in1(N__85041),
            .in2(N__77460),
            .in3(N__55290),
            .lcout(data_out_frame_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__3__5466_LC_15_17_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__3__5466_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__3__5466_LC_15_17_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_7__3__5466_LC_15_17_4  (
            .in0(N__85040),
            .in1(N__84628),
            .in2(N__72077),
            .in3(N__57528),
            .lcout(data_out_frame_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36209_bdd_4_lut_LC_15_17_5 .C_ON=1'b0;
    defparam \c0.n36209_bdd_4_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.n36209_bdd_4_lut_LC_15_17_5 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n36209_bdd_4_lut_LC_15_17_5  (
            .in0(N__61251),
            .in1(N__55299),
            .in2(N__90394),
            .in3(N__55289),
            .lcout(),
            .ltout(\c0.n36212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30663_4_lut_LC_15_17_6 .C_ON=1'b0;
    defparam \c0.i30663_4_lut_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30663_4_lut_LC_15_17_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i30663_4_lut_LC_15_17_6  (
            .in0(N__90370),
            .in1(N__67494),
            .in2(N__55281),
            .in3(N__90004),
            .lcout(n36092),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i30393_3_lut_4_lut_LC_15_18_2.C_ON=1'b0;
    defparam i30393_3_lut_4_lut_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam i30393_3_lut_4_lut_LC_15_18_2.LUT_INIT=16'b1100101011001100;
    LogicCell40 i30393_3_lut_4_lut_LC_15_18_2 (
            .in0(N__55266),
            .in1(N__57675),
            .in2(N__90794),
            .in3(N__95762),
            .lcout(n35820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_LC_15_18_3 .C_ON=1'b0;
    defparam \c0.i14_2_lut_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_LC_15_18_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i14_2_lut_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__58009),
            .in2(_gnd_net_),
            .in3(N__57788),
            .lcout(\c0.n161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_15_18_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_15_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_15_18_4  (
            .in0(N__96014),
            .in1(N__57599),
            .in2(_gnd_net_),
            .in3(N__57506),
            .lcout(\c0.n11_adj_4626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1587_LC_15_18_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1587_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1587_LC_15_18_5 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \c0.i2_4_lut_adj_1587_LC_15_18_5  (
            .in0(N__91078),
            .in1(N__91259),
            .in2(N__93234),
            .in3(N__55248),
            .lcout(\c0.n30906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23139_2_lut_LC_15_18_7 .C_ON=1'b0;
    defparam \c0.i23139_2_lut_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i23139_2_lut_LC_15_18_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i23139_2_lut_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__92599),
            .in2(_gnd_net_),
            .in3(N__65356),
            .lcout(\c0.n5024 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30569_3_lut_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.rx.i30569_3_lut_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30569_3_lut_LC_15_19_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.rx.i30569_3_lut_LC_15_19_0  (
            .in0(N__55803),
            .in1(N__65080),
            .in2(_gnd_net_),
            .in3(N__55916),
            .lcout(),
            .ltout(n35991_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_15_19_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_15_19_1 .LUT_INIT=16'b0000000000100111;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_15_19_1  (
            .in0(N__65145),
            .in1(N__55635),
            .in2(N__55347),
            .in3(N__76995),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30667_4_lut_LC_15_19_2 .C_ON=1'b0;
    defparam \c0.i30667_4_lut_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i30667_4_lut_LC_15_19_2 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \c0.i30667_4_lut_LC_15_19_2  (
            .in0(N__60981),
            .in1(N__90045),
            .in2(N__90393),
            .in3(N__55344),
            .lcout(n36096),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_15_19_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_15_19_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_15_19_3  (
            .in0(N__65079),
            .in1(_gnd_net_),
            .in2(N__55932),
            .in3(N__55802),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_LC_15_19_4 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_15_19_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_3_lut_LC_15_19_4  (
            .in0(N__55548),
            .in1(N__55435),
            .in2(_gnd_net_),
            .in3(N__55613),
            .lcout(\c0.rx.n28401 ),
            .ltout(\c0.rx.n28401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_15_19_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_15_19_5 .LUT_INIT=16'b1010111101010101;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_LC_15_19_5  (
            .in0(N__65081),
            .in1(_gnd_net_),
            .in2(N__55338),
            .in3(N__58054),
            .lcout(),
            .ltout(n28381_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_15_19_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_15_19_6 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_15_19_6  (
            .in0(N__76994),
            .in1(N__65146),
            .in2(N__55335),
            .in3(N__55332),
            .lcout(\c0.rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__6__5463_LC_15_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__6__5463_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__6__5463_LC_15_19_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_7__6__5463_LC_15_19_7  (
            .in0(N__85199),
            .in1(N__84554),
            .in2(N__76750),
            .in3(N__55326),
            .lcout(data_out_frame_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_15_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_15_20_0  (
            .in0(N__55325),
            .in1(N__61287),
            .in2(_gnd_net_),
            .in3(N__96107),
            .lcout(\c0.n5_adj_4624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_1329_LC_15_20_1 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_1329_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_1329_LC_15_20_1 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.rx.i2_3_lut_adj_1329_LC_15_20_1  (
            .in0(N__77095),
            .in1(N__77046),
            .in2(_gnd_net_),
            .in3(N__77021),
            .lcout(\c0.rx.r_SM_Main_2_N_3687_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30640_2_lut_3_lut_4_lut_LC_15_20_2 .C_ON=1'b0;
    defparam \c0.rx.i30640_2_lut_3_lut_4_lut_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30640_2_lut_3_lut_4_lut_LC_15_20_2 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \c0.rx.i30640_2_lut_3_lut_4_lut_LC_15_20_2  (
            .in0(N__77048),
            .in1(N__65074),
            .in2(N__77030),
            .in3(N__77096),
            .lcout(n35992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i23489_2_lut_3_lut_LC_15_20_3 .C_ON=1'b0;
    defparam \c0.rx.i23489_2_lut_3_lut_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i23489_2_lut_3_lut_LC_15_20_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.rx.i23489_2_lut_3_lut_LC_15_20_3  (
            .in0(N__77094),
            .in1(N__77047),
            .in2(_gnd_net_),
            .in3(N__77020),
            .lcout(\c0.rx.r_SM_Main_2_N_3681_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_3681_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_15_20_4 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_15_20_4 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \c0.rx.i2_4_lut_LC_15_20_4  (
            .in0(N__76993),
            .in1(N__65135),
            .in2(N__55629),
            .in3(N__65073),
            .lcout(\c0.rx.n34091 ),
            .ltout(\c0.rx.n34091_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_15_20_5 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_15_20_5 .LUT_INIT=16'b1100011000000000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_15_20_5  (
            .in0(N__55606),
            .in1(N__55550),
            .in2(N__55566),
            .in3(N__55500),
            .lcout(\c0.rx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_LC_15_20_6 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_LC_15_20_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.rx.i1_3_lut_LC_15_20_6  (
            .in0(N__55506),
            .in1(N__65136),
            .in2(_gnd_net_),
            .in3(N__55489),
            .lcout(\c0.rx.n29888 ),
            .ltout(\c0.rx.n29888_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_15_20_7 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_15_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_15_20_7 .LUT_INIT=16'b1011000001000000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_15_20_7  (
            .in0(N__55490),
            .in1(N__55476),
            .in2(N__55461),
            .in3(N__55446),
            .lcout(\c0.rx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97617),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_15_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_15_21_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i48_LC_15_21_0  (
            .in0(N__68305),
            .in1(N__78621),
            .in2(N__55398),
            .in3(N__79997),
            .lcout(\c0.data_in_frame_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97630),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_1331_LC_15_21_1 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_1331_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_1331_LC_15_21_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.rx.i2_3_lut_adj_1331_LC_15_21_1  (
            .in0(N__58497),
            .in1(N__58524),
            .in2(_gnd_net_),
            .in3(N__58554),
            .lcout(\c0.rx.n18092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30344_2_lut_LC_15_21_2 .C_ON=1'b0;
    defparam \c0.rx.i30344_2_lut_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30344_2_lut_LC_15_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i30344_2_lut_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__77081),
            .in2(_gnd_net_),
            .in3(N__58498),
            .lcout(),
            .ltout(\c0.rx.n35769_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_LC_15_21_3 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \c0.rx.i3_4_lut_LC_15_21_3  (
            .in0(N__55926),
            .in1(N__77026),
            .in2(N__55806),
            .in3(N__55800),
            .lcout(\c0.rx.n35738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_15_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_15_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_15_21_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i29_LC_15_21_5  (
            .in0(N__78332),
            .in1(N__83732),
            .in2(N__55774),
            .in3(N__84230),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97630),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_1332_LC_15_21_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_1332_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_1332_LC_15_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_1332_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__77025),
            .in2(_gnd_net_),
            .in3(N__77082),
            .lcout(),
            .ltout(\c0.rx.n33223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30607_4_lut_LC_15_21_7 .C_ON=1'b0;
    defparam \c0.rx.i30607_4_lut_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30607_4_lut_LC_15_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i30607_4_lut_LC_15_21_7  (
            .in0(N__58499),
            .in1(N__58525),
            .in2(N__55743),
            .in3(N__58555),
            .lcout(\c0.rx.n35950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i106_LC_15_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i106_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i106_LC_15_22_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i106_LC_15_22_1  (
            .in0(N__68588),
            .in1(N__78574),
            .in2(N__55728),
            .in3(N__75229),
            .lcout(\c0.data_in_frame_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1352_LC_15_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1352_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1352_LC_15_22_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1352_LC_15_22_2  (
            .in0(N__78431),
            .in1(N__57797),
            .in2(N__58020),
            .in3(N__92750),
            .lcout(\c0.n33233 ),
            .ltout(\c0.n33233_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i188_LC_15_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i188_LC_15_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i188_LC_15_22_3 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \c0.data_in_frame_0__i188_LC_15_22_3  (
            .in0(N__78987),
            .in1(N__62261),
            .in2(N__55698),
            .in3(N__58921),
            .lcout(\c0.data_in_frame_23_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1937_LC_15_22_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1937_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1937_LC_15_22_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i11_4_lut_adj_1937_LC_15_22_4  (
            .in0(N__55695),
            .in1(N__55665),
            .in2(N__55656),
            .in3(N__61767),
            .lcout(\c0.n29_adj_4761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_2050_LC_15_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_2050_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_2050_LC_15_22_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.i1_2_lut_adj_2050_LC_15_22_5  (
            .in0(N__78685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74390),
            .lcout(\c0.n33257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1501_LC_15_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1501_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1501_LC_15_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1501_LC_15_23_0  (
            .in0(N__56059),
            .in1(N__62325),
            .in2(N__56040),
            .in3(N__59228),
            .lcout(\c0.n18487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i192_LC_15_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i192_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i192_LC_15_23_1 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \c0.data_in_frame_0__i192_LC_15_23_1  (
            .in0(N__80120),
            .in1(N__72799),
            .in2(N__62259),
            .in3(N__56021),
            .lcout(\c0.data_in_frame_23_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1806_LC_15_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1806_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1806_LC_15_23_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1806_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__56290),
            .in2(_gnd_net_),
            .in3(N__58726),
            .lcout(\c0.n33813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i112_LC_15_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i112_LC_15_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i112_LC_15_23_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i112_LC_15_23_4  (
            .in0(N__78640),
            .in1(N__68580),
            .in2(N__55991),
            .in3(N__80121),
            .lcout(\c0.data_in_frame_13_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i146_LC_15_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i146_LC_15_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i146_LC_15_23_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i146_LC_15_23_6  (
            .in0(N__80299),
            .in1(N__56291),
            .in2(N__72879),
            .in3(N__75230),
            .lcout(\c0.data_in_frame_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97661),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i19_LC_15_23_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i19_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i19_LC_15_23_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i19_LC_15_23_7  (
            .in0(N__72046),
            .in1(N__61503),
            .in2(_gnd_net_),
            .in3(N__86041),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97661),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1934_LC_15_24_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1934_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1934_LC_15_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1934_LC_15_24_0  (
            .in0(N__79545),
            .in1(N__56135),
            .in2(N__58743),
            .in3(N__55956),
            .lcout(),
            .ltout(\c0.n34727_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1940_LC_15_24_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1940_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1940_LC_15_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_1940_LC_15_24_1  (
            .in0(N__68766),
            .in1(N__56145),
            .in2(N__55947),
            .in3(N__55944),
            .lcout(\c0.n33_adj_4764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1935_LC_15_24_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1935_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1935_LC_15_24_2 .LUT_INIT=16'b1101111011101101;
    LogicCell40 \c0.i6_4_lut_adj_1935_LC_15_24_2  (
            .in0(N__56166),
            .in1(N__56151),
            .in2(N__66026),
            .in3(N__58803),
            .lcout(\c0.n24_adj_4760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i226_LC_15_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i226_LC_15_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i226_LC_15_24_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i226_LC_15_24_3  (
            .in0(N__75351),
            .in1(N__73908),
            .in2(N__56139),
            .in3(N__79847),
            .lcout(\c0.data_in_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i164_LC_15_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i164_LC_15_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i164_LC_15_24_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i164_LC_15_24_4  (
            .in0(N__73907),
            .in1(N__78965),
            .in2(N__56277),
            .in3(N__72869),
            .lcout(\c0.data_in_frame_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i163_LC_15_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i163_LC_15_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i163_LC_15_24_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i163_LC_15_24_6  (
            .in0(N__73906),
            .in1(N__72868),
            .in2(N__56091),
            .in3(N__80711),
            .lcout(\c0.data_in_frame_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i186_LC_15_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i186_LC_15_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i186_LC_15_25_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i186_LC_15_25_0  (
            .in0(N__75365),
            .in1(N__62229),
            .in2(N__65771),
            .in3(N__72870),
            .lcout(\c0.data_in_frame_23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97692),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1682_LC_15_25_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1682_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1682_LC_15_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1682_LC_15_25_1  (
            .in0(N__56382),
            .in1(N__56352),
            .in2(_gnd_net_),
            .in3(N__56331),
            .lcout(),
            .ltout(\c0.n17531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1666_LC_15_25_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1666_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1666_LC_15_25_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1666_LC_15_25_2  (
            .in0(N__72521),
            .in1(N__56259),
            .in2(N__56127),
            .in3(N__68785),
            .lcout(\c0.n33539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1696_LC_15_25_3 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1696_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1696_LC_15_25_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i18_4_lut_adj_1696_LC_15_25_3  (
            .in0(N__56455),
            .in1(N__58789),
            .in2(N__56124),
            .in3(N__72522),
            .lcout(\c0.n42_adj_4703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1685_LC_15_25_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1685_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1685_LC_15_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1685_LC_15_25_4  (
            .in0(N__56100),
            .in1(N__56087),
            .in2(_gnd_net_),
            .in3(N__56310),
            .lcout(\c0.n18568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1563_LC_15_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1563_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1563_LC_15_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1563_LC_15_25_5  (
            .in0(N__56381),
            .in1(N__56351),
            .in2(N__56301),
            .in3(N__56330),
            .lcout(\c0.n18974 ),
            .ltout(\c0.n18974_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1664_LC_15_25_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1664_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1664_LC_15_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1664_LC_15_25_6  (
            .in0(N__56273),
            .in1(N__58857),
            .in2(N__56304),
            .in3(N__56454),
            .lcout(\c0.n35211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1629_LC_15_25_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1629_LC_15_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1629_LC_15_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1629_LC_15_25_7  (
            .in0(N__56300),
            .in1(N__56272),
            .in2(_gnd_net_),
            .in3(N__58733),
            .lcout(\c0.n6_adj_4661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i99_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i99_LC_15_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i99_LC_15_26_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i99_LC_15_26_0  (
            .in0(N__80688),
            .in1(N__58380),
            .in2(N__73921),
            .in3(N__56249),
            .lcout(\c0.data_in_frame_12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i122_LC_15_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i122_LC_15_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i122_LC_15_26_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.data_in_frame_0__i122_LC_15_26_1  (
            .in0(N__58378),
            .in1(N__62258),
            .in2(N__56229),
            .in3(N__75335),
            .lcout(\c0.data_in_frame_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_2026_LC_15_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_2026_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_2026_LC_15_26_2 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_2026_LC_15_26_2  (
            .in0(N__67939),
            .in1(N__74543),
            .in2(N__56199),
            .in3(_gnd_net_),
            .lcout(\c0.n32310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1561_LC_15_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1561_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1561_LC_15_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1561_LC_15_26_3  (
            .in0(N__58922),
            .in1(N__65761),
            .in2(_gnd_net_),
            .in3(N__67938),
            .lcout(\c0.n33864 ),
            .ltout(\c0.n33864_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1692_LC_15_26_4 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1692_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1692_LC_15_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_1692_LC_15_26_4  (
            .in0(N__59056),
            .in1(N__59160),
            .in2(N__56181),
            .in3(N__56177),
            .lcout(\c0.n40_adj_4700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i178_LC_15_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i178_LC_15_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i178_LC_15_26_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i178_LC_15_26_5  (
            .in0(N__75289),
            .in1(N__89759),
            .in2(N__73045),
            .in3(N__59057),
            .lcout(\c0.data_in_frame_22_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i117_LC_15_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i117_LC_15_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i117_LC_15_26_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i117_LC_15_26_6  (
            .in0(N__89758),
            .in1(N__58379),
            .in2(N__56520),
            .in3(N__84254),
            .lcout(\c0.data_in_frame_14_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i131_LC_15_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i131_LC_15_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i131_LC_15_26_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i131_LC_15_26_7  (
            .in0(N__81271),
            .in1(N__72986),
            .in2(N__56728),
            .in3(N__80689),
            .lcout(\c0.data_in_frame_16_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97708),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1653_LC_15_27_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1653_LC_15_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1653_LC_15_27_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i12_4_lut_adj_1653_LC_15_27_0  (
            .in0(N__56505),
            .in1(N__56397),
            .in2(N__56496),
            .in3(N__56460),
            .lcout(\c0.n32026 ),
            .ltout(\c0.n32026_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1637_LC_15_27_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1637_LC_15_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1637_LC_15_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1637_LC_15_27_1  (
            .in0(N__74347),
            .in1(N__74273),
            .in2(N__56427),
            .in3(N__65589),
            .lcout(\c0.n33991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_15_27_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_15_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_15_27_2  (
            .in0(N__56424),
            .in1(N__79463),
            .in2(N__56646),
            .in3(N__56418),
            .lcout(\c0.n24_adj_4671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_15_27_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_15_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_15_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_LC_15_27_3  (
            .in0(N__74346),
            .in1(N__65677),
            .in2(N__74279),
            .in3(N__56390),
            .lcout(\c0.n10_adj_4669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1777_LC_15_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1777_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1777_LC_15_27_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1777_LC_15_27_4  (
            .in0(_gnd_net_),
            .in1(N__74263),
            .in2(_gnd_net_),
            .in3(N__74345),
            .lcout(\c0.n18415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1639_LC_15_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1639_LC_15_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1639_LC_15_27_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1639_LC_15_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__65938),
            .in3(N__62039),
            .lcout(\c0.n6_adj_4666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1705_LC_15_27_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1705_LC_15_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1705_LC_15_27_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1705_LC_15_27_7  (
            .in0(N__79544),
            .in1(N__65678),
            .in2(N__74225),
            .in3(N__56391),
            .lcout(\c0.n7_adj_4662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1649_LC_15_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1649_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1649_LC_15_28_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1649_LC_15_28_0  (
            .in0(_gnd_net_),
            .in1(N__67937),
            .in2(_gnd_net_),
            .in3(N__74549),
            .lcout(\c0.n6462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1800_LC_15_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1800_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1800_LC_15_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1800_LC_15_28_1  (
            .in0(_gnd_net_),
            .in1(N__56721),
            .in2(_gnd_net_),
            .in3(N__56688),
            .lcout(\c0.n33618 ),
            .ltout(\c0.n33618_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1698_LC_15_28_2 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1698_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1698_LC_15_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1698_LC_15_28_2  (
            .in0(N__56586),
            .in1(N__74550),
            .in2(N__56658),
            .in3(N__62316),
            .lcout(\c0.n41_adj_4704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1651_LC_15_28_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1651_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1651_LC_15_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1651_LC_15_28_3  (
            .in0(N__56624),
            .in1(N__62407),
            .in2(N__56655),
            .in3(N__65478),
            .lcout(\c0.n22_adj_4670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_1694_LC_15_28_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_1694_LC_15_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_1694_LC_15_28_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i15_4_lut_adj_1694_LC_15_28_4  (
            .in0(N__56637),
            .in1(N__56625),
            .in2(N__74714),
            .in3(N__66386),
            .lcout(\c0.n39_adj_4702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1774_LC_15_28_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1774_LC_15_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1774_LC_15_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1774_LC_15_28_5  (
            .in0(N__62411),
            .in1(N__58959),
            .in2(_gnd_net_),
            .in3(N__56532),
            .lcout(\c0.n31417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1785_LC_15_28_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1785_LC_15_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1785_LC_15_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1785_LC_15_28_6  (
            .in0(N__56585),
            .in1(N__56560),
            .in2(_gnd_net_),
            .in3(N__56541),
            .lcout(\c0.n17702 ),
            .ltout(\c0.n17702_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1513_LC_15_28_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1513_LC_15_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1513_LC_15_28_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1513_LC_15_28_7  (
            .in0(N__59366),
            .in1(_gnd_net_),
            .in2(N__56526),
            .in3(N__58958),
            .lcout(\c0.n33598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_2_lut_LC_16_6_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_2_lut_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_2_lut_LC_16_6_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1482_2_lut_LC_16_6_0  (
            .in0(N__60147),
            .in1(N__60146),
            .in2(N__56998),
            .in3(N__56523),
            .lcout(\quad_counter0.n2219 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\quad_counter0.n30230 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_3_lut_LC_16_6_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_3_lut_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_3_lut_LC_16_6_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1482_3_lut_LC_16_6_1  (
            .in0(N__56913),
            .in1(N__56912),
            .in2(N__57037),
            .in3(N__56895),
            .lcout(\quad_counter0.n2218 ),
            .ltout(),
            .carryin(\quad_counter0.n30230 ),
            .carryout(\quad_counter0.n30231 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_4_lut_LC_16_6_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_4_lut_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_4_lut_LC_16_6_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1482_4_lut_LC_16_6_2  (
            .in0(N__56892),
            .in1(N__56891),
            .in2(N__56999),
            .in3(N__56868),
            .lcout(\quad_counter0.n2217 ),
            .ltout(),
            .carryin(\quad_counter0.n30231 ),
            .carryout(\quad_counter0.n30232 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_5_lut_LC_16_6_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_5_lut_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_5_lut_LC_16_6_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1482_5_lut_LC_16_6_3  (
            .in0(N__56864),
            .in1(N__56863),
            .in2(N__57002),
            .in3(N__56844),
            .lcout(\quad_counter0.n2216 ),
            .ltout(),
            .carryin(\quad_counter0.n30232 ),
            .carryout(\quad_counter0.n30233 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_6_lut_LC_16_6_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_6_lut_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_6_lut_LC_16_6_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1482_6_lut_LC_16_6_4  (
            .in0(N__56841),
            .in1(N__56840),
            .in2(N__57000),
            .in3(N__56823),
            .lcout(\quad_counter0.n2215 ),
            .ltout(),
            .carryin(\quad_counter0.n30233 ),
            .carryout(\quad_counter0.n30234 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_7_lut_LC_16_6_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_7_lut_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_7_lut_LC_16_6_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1482_7_lut_LC_16_6_5  (
            .in0(N__56820),
            .in1(N__56819),
            .in2(N__57003),
            .in3(N__56802),
            .lcout(\quad_counter0.n2214 ),
            .ltout(),
            .carryin(\quad_counter0.n30234 ),
            .carryout(\quad_counter0.n30235 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_8_lut_LC_16_6_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_8_lut_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_8_lut_LC_16_6_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1482_8_lut_LC_16_6_6  (
            .in0(N__56799),
            .in1(N__56798),
            .in2(N__57001),
            .in3(N__56781),
            .lcout(\quad_counter0.n2213 ),
            .ltout(),
            .carryin(\quad_counter0.n30235 ),
            .carryout(\quad_counter0.n30236 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_9_lut_LC_16_6_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_9_lut_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_9_lut_LC_16_6_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1482_9_lut_LC_16_6_7  (
            .in0(N__56778),
            .in1(N__56777),
            .in2(N__57038),
            .in3(N__56757),
            .lcout(\quad_counter0.n2212 ),
            .ltout(),
            .carryin(\quad_counter0.n30236 ),
            .carryout(\quad_counter0.n30237 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_10_lut_LC_16_7_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1482_10_lut_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_10_lut_LC_16_7_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1482_10_lut_LC_16_7_0  (
            .in0(N__56754),
            .in1(N__56753),
            .in2(N__57039),
            .in3(N__56733),
            .lcout(\quad_counter0.n2211 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\quad_counter0.n30238 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1482_11_lut_LC_16_7_1 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1482_11_lut_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1482_11_lut_LC_16_7_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1482_11_lut_LC_16_7_1  (
            .in0(N__57065),
            .in1(N__57066),
            .in2(N__57036),
            .in3(N__57042),
            .lcout(\quad_counter0.n2210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30730_1_lut_LC_16_7_2 .C_ON=1'b0;
    defparam \quad_counter0.i30730_1_lut_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30730_1_lut_LC_16_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter0.i30730_1_lut_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57023),
            .lcout(\quad_counter0.n36157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_delayed_76_LC_16_7_6 .C_ON=1'b0;
    defparam \quad_counter1.A_delayed_76_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.A_delayed_76_LC_16_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter1.A_delayed_76_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59446),
            .lcout(\quad_counter1.A_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97538),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_3_lut_LC_16_8_0 .C_ON=1'b0;
    defparam \quad_counter0.i5_3_lut_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_3_lut_LC_16_8_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \quad_counter0.i5_3_lut_LC_16_8_0  (
            .in0(N__59588),
            .in1(N__59555),
            .in2(_gnd_net_),
            .in3(N__59627),
            .lcout(\quad_counter0.n14_adj_4418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1204_LC_16_10_0 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1204_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1204_LC_16_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1204_LC_16_10_0  (
            .in0(N__63525),
            .in1(N__63072),
            .in2(N__63492),
            .in3(N__63393),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_4_lut_adj_1206_LC_16_10_1 .C_ON=1'b0;
    defparam \quad_counter0.i1_4_lut_adj_1206_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_4_lut_adj_1206_LC_16_10_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i1_4_lut_adj_1206_LC_16_10_1  (
            .in0(N__63456),
            .in1(N__63426),
            .in2(N__56961),
            .in3(N__63321),
            .lcout(\quad_counter0.n7_adj_4393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i6_4_lut_adj_1242_LC_16_10_4 .C_ON=1'b0;
    defparam \quad_counter0.i6_4_lut_adj_1242_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i6_4_lut_adj_1242_LC_16_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i6_4_lut_adj_1242_LC_16_10_4  (
            .in0(N__59574),
            .in1(N__59541),
            .in2(N__59613),
            .in3(N__57237),
            .lcout(),
            .ltout(\quad_counter0.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i8_4_lut_adj_1243_LC_16_10_5 .C_ON=1'b0;
    defparam \quad_counter0.i8_4_lut_adj_1243_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i8_4_lut_adj_1243_LC_16_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i8_4_lut_adj_1243_LC_16_10_5  (
            .in0(N__56958),
            .in1(N__59520),
            .in2(N__56949),
            .in3(N__59499),
            .lcout(n34523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i10_4_lut_adj_1241_LC_16_11_0 .C_ON=1'b0;
    defparam \quad_counter0.i10_4_lut_adj_1241_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i10_4_lut_adj_1241_LC_16_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i10_4_lut_adj_1241_LC_16_11_0  (
            .in0(N__56946),
            .in1(N__56937),
            .in2(N__56928),
            .in3(N__56919),
            .lcout(\quad_counter0.n28_adj_4342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30648_3_lut_LC_16_11_1 .C_ON=1'b0;
    defparam \quad_counter0.i30648_3_lut_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30648_3_lut_LC_16_11_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter0.i30648_3_lut_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__57075),
            .in2(N__57177),
            .in3(N__57297),
            .lcout(),
            .ltout(\quad_counter0.n35977_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i47_4_lut_LC_16_11_2 .C_ON=1'b0;
    defparam \quad_counter0.i47_4_lut_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i47_4_lut_LC_16_11_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \quad_counter0.i47_4_lut_LC_16_11_2  (
            .in0(N__57183),
            .in1(N__57264),
            .in2(N__57252),
            .in3(N__57249),
            .lcout(\quad_counter0.n34205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i13_4_lut_adj_1208_LC_16_11_4 .C_ON=1'b0;
    defparam \quad_counter0.i13_4_lut_adj_1208_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i13_4_lut_adj_1208_LC_16_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i13_4_lut_adj_1208_LC_16_11_4  (
            .in0(N__57231),
            .in1(N__57225),
            .in2(N__57219),
            .in3(N__57210),
            .lcout(),
            .ltout(\quad_counter0.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i16_4_lut_LC_16_11_5 .C_ON=1'b0;
    defparam \quad_counter0.i16_4_lut_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i16_4_lut_LC_16_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i16_4_lut_LC_16_11_5  (
            .in0(N__57204),
            .in1(N__57198),
            .in2(N__57192),
            .in3(N__57189),
            .lcout(\quad_counter0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_2_lut_LC_16_12_0 .C_ON=1'b1;
    defparam \quad_counter0.add_8361_2_lut_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_2_lut_LC_16_12_0 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter0.add_8361_2_lut_LC_16_12_0  (
            .in0(N__57339),
            .in1(N__59985),
            .in2(_gnd_net_),
            .in3(N__57168),
            .lcout(\quad_counter0.n35978 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\quad_counter0.n30453 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_3_lut_LC_16_12_1 .C_ON=1'b1;
    defparam \quad_counter0.add_8361_3_lut_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_3_lut_LC_16_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_8361_3_lut_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__98966),
            .in2(N__57165),
            .in3(N__57138),
            .lcout(\quad_counter0.n12904 ),
            .ltout(),
            .carryin(\quad_counter0.n30453 ),
            .carryout(\quad_counter0.n30454 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_4_lut_LC_16_12_2 .C_ON=1'b1;
    defparam \quad_counter0.add_8361_4_lut_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_4_lut_LC_16_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_8361_4_lut_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57135),
            .in3(N__57108),
            .lcout(\quad_counter0.n12903 ),
            .ltout(),
            .carryin(\quad_counter0.n30454 ),
            .carryout(\quad_counter0.n30455 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_5_lut_LC_16_12_3 .C_ON=1'b1;
    defparam \quad_counter0.add_8361_5_lut_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_5_lut_LC_16_12_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter0.add_8361_5_lut_LC_16_12_3  (
            .in0(N__57105),
            .in1(_gnd_net_),
            .in2(N__57099),
            .in3(N__57069),
            .lcout(\quad_counter0.n9 ),
            .ltout(),
            .carryin(\quad_counter0.n30455 ),
            .carryout(\quad_counter0.n30456 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_6_lut_LC_16_12_4 .C_ON=1'b1;
    defparam \quad_counter0.add_8361_6_lut_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_6_lut_LC_16_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_8361_6_lut_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57393),
            .in3(N__57366),
            .lcout(\quad_counter0.n12901 ),
            .ltout(),
            .carryin(\quad_counter0.n30456 ),
            .carryout(\quad_counter0.n30457 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_7_lut_LC_16_12_5 .C_ON=1'b1;
    defparam \quad_counter0.add_8361_7_lut_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_7_lut_LC_16_12_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter0.add_8361_7_lut_LC_16_12_5  (
            .in0(N__57363),
            .in1(N__57357),
            .in2(_gnd_net_),
            .in3(N__57333),
            .lcout(\quad_counter0.n8_adj_4375 ),
            .ltout(),
            .carryin(\quad_counter0.n30457 ),
            .carryout(\quad_counter0.n30458 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_8361_8_lut_LC_16_12_6 .C_ON=1'b0;
    defparam \quad_counter0.add_8361_8_lut_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_8361_8_lut_LC_16_12_6 .LUT_INIT=16'b1110110111011110;
    LogicCell40 \quad_counter0.add_8361_8_lut_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__57330),
            .in2(N__57324),
            .in3(N__57300),
            .lcout(\quad_counter0.n10_adj_4347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_4_lut_adj_1219_LC_16_13_0 .C_ON=1'b0;
    defparam \quad_counter0.i2_4_lut_adj_1219_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_4_lut_adj_1219_LC_16_13_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i2_4_lut_adj_1219_LC_16_13_0  (
            .in0(N__60683),
            .in1(N__57282),
            .in2(N__60661),
            .in3(N__60785),
            .lcout(\quad_counter0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23623_2_lut_LC_16_13_3 .C_ON=1'b0;
    defparam \quad_counter0.i23623_2_lut_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23623_2_lut_LC_16_13_3 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \quad_counter0.i23623_2_lut_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__60202),
            .in2(N__60226),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\quad_counter0.n28339_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1217_LC_16_13_4 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1217_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1217_LC_16_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1217_LC_16_13_4  (
            .in0(N__60626),
            .in1(N__60712),
            .in2(N__57285),
            .in3(N__60740),
            .lcout(\quad_counter0.n10_adj_4400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_2_lut_adj_1216_LC_16_13_5 .C_ON=1'b0;
    defparam \quad_counter0.i1_2_lut_adj_1216_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_2_lut_adj_1216_LC_16_13_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i1_2_lut_adj_1216_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60571),
            .in3(N__60536),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i7_4_lut_adj_1218_LC_16_13_6 .C_ON=1'b0;
    defparam \quad_counter0.i7_4_lut_adj_1218_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i7_4_lut_adj_1218_LC_16_13_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i7_4_lut_adj_1218_LC_16_13_6  (
            .in0(N__60869),
            .in1(N__60904),
            .in2(N__57276),
            .in3(N__60842),
            .lcout(\quad_counter0.n16_adj_4401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1602_LC_16_14_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1602_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1602_LC_16_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i2_2_lut_adj_1602_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__90695),
            .in2(_gnd_net_),
            .in3(N__95741),
            .lcout(),
            .ltout(\c0.n6_adj_4647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1603_LC_16_14_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1603_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1603_LC_16_14_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \c0.i3_4_lut_adj_1603_LC_16_14_1  (
            .in0(N__89974),
            .in1(N__90231),
            .in2(N__57495),
            .in3(N__95966),
            .lcout(\c0.n28313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__2__5435_LC_16_15_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__2__5435_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__2__5435_LC_16_15_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_11__2__5435_LC_16_15_0  (
            .in0(N__85071),
            .in1(N__84639),
            .in2(N__86367),
            .in3(N__57420),
            .lcout(data_out_frame_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__2__5459_LC_16_15_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__2__5459_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__2__5459_LC_16_15_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.data_out_frame_8__2__5459_LC_16_15_1  (
            .in0(N__84638),
            .in1(N__85072),
            .in2(N__57462),
            .in3(N__72381),
            .lcout(data_out_frame_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36203_bdd_4_lut_LC_16_15_4 .C_ON=1'b0;
    defparam \c0.n36203_bdd_4_lut_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.n36203_bdd_4_lut_LC_16_15_4 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n36203_bdd_4_lut_LC_16_15_4  (
            .in0(N__57476),
            .in1(N__57399),
            .in2(N__90380),
            .in3(N__57458),
            .lcout(\c0.n36206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2064_LC_16_15_6.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2064_LC_16_15_6.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2064_LC_16_15_6.LUT_INIT=16'b1100110010101100;
    LogicCell40 i24_3_lut_4_lut_adj_2064_LC_16_15_6 (
            .in0(N__60759),
            .in1(N__60954),
            .in2(N__95789),
            .in3(N__90774),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__2__5443_LC_16_16_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__2__5443_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__2__5443_LC_16_16_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_10__2__5443_LC_16_16_0  (
            .in0(N__57408),
            .in1(N__84615),
            .in2(N__85163),
            .in3(N__72273),
            .lcout(data_out_frame_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97568),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2065_LC_16_16_1.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2065_LC_16_16_1.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2065_LC_16_16_1.LUT_INIT=16'b1010111010100010;
    LogicCell40 i24_3_lut_4_lut_adj_2065_LC_16_16_1 (
            .in0(N__71739),
            .in1(N__95772),
            .in2(N__90785),
            .in3(N__57543),
            .lcout(n10_adj_4806),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_16_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_16_16_2 .LUT_INIT=16'b1100000011111010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_16_16_2  (
            .in0(N__57429),
            .in1(N__68118),
            .in2(N__96109),
            .in3(N__90044),
            .lcout(\c0.n6_adj_4514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30774_LC_16_16_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30774_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30774_LC_16_16_5 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_30774_LC_16_16_5  (
            .in0(N__57419),
            .in1(N__57407),
            .in2(N__90371),
            .in3(N__96016),
            .lcout(\c0.n36203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__0__5461_LC_16_16_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__0__5461_LC_16_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__0__5461_LC_16_16_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_8__0__5461_LC_16_16_7  (
            .in0(N__84614),
            .in1(N__85033),
            .in2(N__73236),
            .in3(N__57588),
            .lcout(data_out_frame_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_16_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_16_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_16_17_0  (
            .in0(N__96021),
            .in1(N__61034),
            .in2(_gnd_net_),
            .in3(N__60923),
            .lcout(\c0.n11_adj_4655 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36191_bdd_4_lut_LC_16_17_1 .C_ON=1'b0;
    defparam \c0.n36191_bdd_4_lut_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.n36191_bdd_4_lut_LC_16_17_1 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n36191_bdd_4_lut_LC_16_17_1  (
            .in0(N__57576),
            .in1(N__61023),
            .in2(N__90378),
            .in3(N__64761),
            .lcout(),
            .ltout(\c0.n36194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30665_4_lut_LC_16_17_2 .C_ON=1'b0;
    defparam \c0.i30665_4_lut_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i30665_4_lut_LC_16_17_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.i30665_4_lut_LC_16_17_2  (
            .in0(N__90339),
            .in1(N__90040),
            .in2(N__57552),
            .in3(N__57549),
            .lcout(n36094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i7_4_lut_LC_16_17_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i7_4_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i7_4_lut_LC_16_17_3 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i7_4_lut_LC_16_17_3  (
            .in0(N__57537),
            .in1(N__90047),
            .in2(N__90377),
            .in3(N__61077),
            .lcout(\c0.n7_adj_4499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_17_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_16_17_5  (
            .in0(N__57527),
            .in1(N__57515),
            .in2(_gnd_net_),
            .in3(N__96020),
            .lcout(\c0.n5_adj_4515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__3__5474_LC_16_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__3__5474_LC_16_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__3__5474_LC_16_17_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_6__3__5474_LC_16_17_6  (
            .in0(N__57516),
            .in1(N__84625),
            .in2(N__85250),
            .in3(N__79147),
            .lcout(data_out_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97577),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_per_millisecond_i0_i0_LC_16_18_0 .C_ON=1'b0;
    defparam \quad_counter0.count_per_millisecond_i0_i0_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_per_millisecond_i0_i0_LC_16_18_0 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \quad_counter0.count_per_millisecond_i0_i0_LC_16_18_0  (
            .in0(N__100726),
            .in1(N__60252),
            .in2(N__85631),
            .in3(N__60273),
            .lcout(data_out_frame_29__7__N_1240),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__6__5423_LC_16_18_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__6__5423_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__6__5423_LC_16_18_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_12__6__5423_LC_16_18_3  (
            .in0(N__84624),
            .in1(N__85142),
            .in2(N__77295),
            .in3(N__57507),
            .lcout(data_out_frame_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30391_3_lut_LC_16_18_5 .C_ON=1'b0;
    defparam \c0.i30391_3_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30391_3_lut_LC_16_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i30391_3_lut_LC_16_18_5  (
            .in0(N__95676),
            .in1(N__57681),
            .in2(_gnd_net_),
            .in3(N__90793),
            .lcout(n35818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__6__5439_LC_16_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__6__5439_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__6__5439_LC_16_18_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_10__6__5439_LC_16_18_7  (
            .in0(N__84623),
            .in1(N__85141),
            .in2(N__86280),
            .in3(N__61017),
            .lcout(data_out_frame_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i34_LC_16_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i34_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i34_LC_16_19_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i34_LC_16_19_0  (
            .in0(N__83977),
            .in1(N__73914),
            .in2(N__75344),
            .in3(N__57667),
            .lcout(\c0.data_in_frame_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_16_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_16_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_16_19_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i18_LC_16_19_1  (
            .in0(N__80298),
            .in1(N__83979),
            .in2(N__57639),
            .in3(N__75296),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_16_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_16_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_16_19_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i15_LC_16_19_2  (
            .in0(N__83976),
            .in1(N__87294),
            .in2(N__64825),
            .in3(N__73623),
            .lcout(data_in_frame_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i2_LC_16_19_3 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i2_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i2_LC_16_19_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i2_LC_16_19_3  (
            .in0(N__72188),
            .in1(N__58678),
            .in2(_gnd_net_),
            .in3(N__77630),
            .lcout(control_mode_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__6__5415_LC_16_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__6__5415_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__6__5415_LC_16_19_4 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \c0.data_out_frame_13__6__5415_LC_16_19_4  (
            .in0(N__85052),
            .in1(N__94324),
            .in2(N__84700),
            .in3(N__57600),
            .lcout(data_out_frame_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_16_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_16_19_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i14_LC_16_19_5  (
            .in0(N__75050),
            .in1(N__83978),
            .in2(N__87306),
            .in3(N__72415),
            .lcout(data_in_frame_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30585_3_lut_LC_16_19_6 .C_ON=1'b0;
    defparam \c0.i30585_3_lut_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30585_3_lut_LC_16_19_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \c0.i30585_3_lut_LC_16_19_6  (
            .in0(N__61377),
            .in1(N__96108),
            .in2(_gnd_net_),
            .in3(N__90051),
            .lcout(\c0.n36012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_adj_1330_LC_16_20_0 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_adj_1330_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_adj_1330_LC_16_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i3_4_lut_adj_1330_LC_16_20_0  (
            .in0(N__57695),
            .in1(N__58583),
            .in2(N__58602),
            .in3(N__57718),
            .lcout(\c0.rx.n33168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_16_20_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_16_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_16_20_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_16_20_1  (
            .in0(N__57705),
            .in1(N__58478),
            .in2(N__57723),
            .in3(N__58457),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_16_20_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_16_20_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_16_20_2  (
            .in0(N__57772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_rx_data_ready_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_16_20_3 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_16_20_3 .LUT_INIT=16'b0100000000110011;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_16_20_3  (
            .in0(N__76980),
            .in1(N__65078),
            .in2(N__58062),
            .in3(N__65122),
            .lcout(),
            .ltout(\c0.rx.n19345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_16_20_4 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_16_20_4  (
            .in0(N__65123),
            .in1(N__76981),
            .in2(N__58065),
            .in3(N__57787),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_adj_1327_LC_16_20_5 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_adj_1327_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_adj_1327_LC_16_20_5 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.rx.i3_4_lut_adj_1327_LC_16_20_5  (
            .in0(N__76979),
            .in1(N__65077),
            .in2(N__58061),
            .in3(N__65121),
            .lcout(\c0.rx.n17939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i26_LC_16_20_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i26_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i26_LC_16_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i26_LC_16_20_6  (
            .in0(N__76561),
            .in1(N__64656),
            .in2(_gnd_net_),
            .in3(N__72260),
            .lcout(encoder1_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23184_2_lut_3_lut_LC_16_20_7 .C_ON=1'b0;
    defparam \c0.i23184_2_lut_3_lut_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i23184_2_lut_3_lut_LC_16_20_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.i23184_2_lut_3_lut_LC_16_20_7  (
            .in0(N__58005),
            .in1(N__57771),
            .in2(_gnd_net_),
            .in3(N__92838),
            .lcout(\c0.n27890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_16_21_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_16_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_2_lut_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__57722),
            .in2(_gnd_net_),
            .in3(N__57699),
            .lcout(n226),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\c0.rx.n30061 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_16_21_1 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i1_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_16_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__57696),
            .in2(_gnd_net_),
            .in3(N__57684),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.rx.n30061 ),
            .carryout(\c0.rx.n30062 ),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \c0.rx.r_Clock_Count__i2_LC_16_21_2 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i2_LC_16_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_16_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__58601),
            .in2(_gnd_net_),
            .in3(N__58587),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.rx.n30062 ),
            .carryout(\c0.rx.n30063 ),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \c0.rx.r_Clock_Count__i3_LC_16_21_3 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i3_LC_16_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_16_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__58584),
            .in2(_gnd_net_),
            .in3(N__58572),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.rx.n30063 ),
            .carryout(\c0.rx.n30064 ),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \c0.rx.r_Clock_Count__i4_LC_16_21_4 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i4_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_16_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__77083),
            .in2(_gnd_net_),
            .in3(N__58569),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.rx.n30064 ),
            .carryout(\c0.rx.n30065 ),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \c0.rx.r_Clock_Count__i5_LC_16_21_5 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i5_LC_16_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_16_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__58559),
            .in2(_gnd_net_),
            .in3(N__58536),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.rx.n30065 ),
            .carryout(\c0.rx.n30066 ),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \c0.rx.r_Clock_Count__i6_LC_16_21_6 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i6_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_16_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__58529),
            .in2(_gnd_net_),
            .in3(N__58506),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.rx.n30066 ),
            .carryout(\c0.rx.n30067 ),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \c0.rx.r_Clock_Count__i7_LC_16_21_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_16_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_16_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__58500),
            .in2(_gnd_net_),
            .in3(N__58503),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97613),
            .ce(N__58482),
            .sr(N__58461));
    defparam \quad_counter0.count_i0_i29_LC_16_22_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i29_LC_16_22_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i29_LC_16_22_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i29_LC_16_22_0  (
            .in0(N__61539),
            .in1(N__86043),
            .in2(_gnd_net_),
            .in3(N__79030),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97627),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i76_LC_16_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i76_LC_16_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i76_LC_16_22_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i76_LC_16_22_1  (
            .in0(N__87295),
            .in1(N__58322),
            .in2(N__58087),
            .in3(N__78986),
            .lcout(\c0.data_in_frame_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97627),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_16_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_16_22_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i49_LC_16_22_2  (
            .in0(N__89797),
            .in1(N__83943),
            .in2(N__58709),
            .in3(N__80930),
            .lcout(\c0.data_in_frame_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97627),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i22_LC_16_22_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i22_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i22_LC_16_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i22_LC_16_22_3  (
            .in0(N__86042),
            .in1(N__61578),
            .in2(_gnd_net_),
            .in3(N__76713),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97627),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i175_LC_16_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i175_LC_16_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i175_LC_16_22_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i175_LC_16_22_4  (
            .in0(N__78641),
            .in1(N__73625),
            .in2(N__61701),
            .in3(N__78430),
            .lcout(\c0.data_in_frame_21_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97627),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_16_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_16_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_16_22_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i11_LC_16_22_6  (
            .in0(N__87297),
            .in1(N__83942),
            .in2(N__58679),
            .in3(N__80708),
            .lcout(data_in_frame_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97627),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i191_LC_16_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i191_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i191_LC_16_23_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.data_in_frame_0__i191_LC_16_23_1  (
            .in0(N__73624),
            .in1(N__62260),
            .in2(N__58793),
            .in3(N__72803),
            .lcout(\c0.data_in_frame_23_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1781_LC_16_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1781_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1781_LC_16_23_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1781_LC_16_23_2  (
            .in0(N__67940),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58920),
            .lcout(\c0.n33329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23156_2_lut_LC_16_23_3 .C_ON=1'b0;
    defparam \c0.i23156_2_lut_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i23156_2_lut_LC_16_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i23156_2_lut_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(N__91209),
            .in2(_gnd_net_),
            .in3(N__91110),
            .lcout(\c0.n27862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2066_LC_16_23_5.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2066_LC_16_23_5.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2066_LC_16_23_5.LUT_INIT=16'b1111010010110000;
    LogicCell40 i24_3_lut_4_lut_adj_2066_LC_16_23_5 (
            .in0(N__90795),
            .in1(N__95795),
            .in2(N__71568),
            .in3(N__58629),
            .lcout(n10_adj_4820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i182_LC_16_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i182_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i182_LC_16_23_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i182_LC_16_23_6  (
            .in0(N__75008),
            .in1(N__89798),
            .in2(N__72880),
            .in3(N__58871),
            .lcout(\c0.data_in_frame_22_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97641),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i21_LC_16_23_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i21_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i21_LC_16_23_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i21_LC_16_23_7  (
            .in0(N__61587),
            .in1(N__86080),
            .in2(_gnd_net_),
            .in3(N__61608),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97641),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1502_LC_16_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1502_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1502_LC_16_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1502_LC_16_24_0  (
            .in0(N__74341),
            .in1(N__61700),
            .in2(N__74292),
            .in3(N__59276),
            .lcout(\c0.n32346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1512_LC_16_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1512_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1512_LC_16_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1512_LC_16_24_1  (
            .in0(N__61699),
            .in1(N__74286),
            .in2(_gnd_net_),
            .in3(N__74340),
            .lcout(),
            .ltout(\c0.n33506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1779_LC_16_24_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1779_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1779_LC_16_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1779_LC_16_24_2  (
            .in0(N__58758),
            .in1(N__65639),
            .in2(N__58839),
            .in3(N__58836),
            .lcout(),
            .ltout(\c0.n12_adj_4710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1780_LC_16_24_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1780_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1780_LC_16_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1780_LC_16_24_3  (
            .in0(N__69075),
            .in1(N__68911),
            .in2(N__58824),
            .in3(N__59109),
            .lcout(\c0.n18784 ),
            .ltout(\c0.n18784_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1912_LC_16_24_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1912_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1912_LC_16_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1912_LC_16_24_4  (
            .in0(N__61671),
            .in1(N__58820),
            .in2(N__58806),
            .in3(N__79509),
            .lcout(\c0.n10_adj_4749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1782_LC_16_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1782_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1782_LC_16_24_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1782_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__65328),
            .in2(_gnd_net_),
            .in3(N__58782),
            .lcout(\c0.n33726 ),
            .ltout(\c0.n33726_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1910_LC_16_24_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1910_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1910_LC_16_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1910_LC_16_24_6  (
            .in0(N__58752),
            .in1(N__69249),
            .in2(N__58746),
            .in3(N__68742),
            .lcout(\c0.n15_adj_4747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i165_LC_16_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i165_LC_16_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i165_LC_16_25_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i165_LC_16_25_0  (
            .in0(N__72866),
            .in1(N__84146),
            .in2(N__58887),
            .in3(N__73909),
            .lcout(\c0.data_in_frame_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1654_LC_16_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1654_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1654_LC_16_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1654_LC_16_25_1  (
            .in0(_gnd_net_),
            .in1(N__58883),
            .in2(_gnd_net_),
            .in3(N__58734),
            .lcout(\c0.n32320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1638_LC_16_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1638_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1638_LC_16_25_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1638_LC_16_25_2  (
            .in0(N__58928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78725),
            .lcout(\c0.n33632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i158_LC_16_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i158_LC_16_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i158_LC_16_25_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i158_LC_16_25_3  (
            .in0(N__75009),
            .in1(N__72867),
            .in2(N__78221),
            .in3(N__58955),
            .lcout(\c0.data_in_frame_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1643_LC_16_25_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1643_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1643_LC_16_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1643_LC_16_25_4  (
            .in0(N__58929),
            .in1(N__73298),
            .in2(N__68718),
            .in3(N__65435),
            .lcout(\c0.n35307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1931_LC_16_25_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1931_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1931_LC_16_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1931_LC_16_25_5  (
            .in0(N__73299),
            .in1(N__65411),
            .in2(N__78729),
            .in3(N__58893),
            .lcout(\c0.n12_adj_4759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i27_LC_16_25_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i27_LC_16_25_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i27_LC_16_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i27_LC_16_25_6  (
            .in0(N__86081),
            .in1(N__61551),
            .in2(_gnd_net_),
            .in3(N__79117),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1663_LC_16_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1663_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1663_LC_16_25_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1663_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__58882),
            .in2(_gnd_net_),
            .in3(N__58872),
            .lcout(\c0.n6_adj_4675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1930_LC_16_26_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1930_LC_16_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1930_LC_16_26_0 .LUT_INIT=16'b1001011011111111;
    LogicCell40 \c0.i7_4_lut_adj_1930_LC_16_26_0  (
            .in0(N__68838),
            .in1(N__58847),
            .in2(N__66138),
            .in3(N__59067),
            .lcout(\c0.n25_adj_4758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i239_LC_16_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i239_LC_16_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i239_LC_16_26_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i239_LC_16_26_1  (
            .in0(N__58848),
            .in1(N__74449),
            .in2(N__73674),
            .in3(N__78656),
            .lcout(\c0.data_in_frame_29_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i176_LC_16_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i176_LC_16_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i176_LC_16_26_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i176_LC_16_26_2  (
            .in0(N__61721),
            .in1(N__80144),
            .in2(N__78657),
            .in3(N__78429),
            .lcout(\c0.data_in_frame_21_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i169_LC_16_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i169_LC_16_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i169_LC_16_26_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i169_LC_16_26_3  (
            .in0(N__80977),
            .in1(N__78655),
            .in2(N__78432),
            .in3(N__59090),
            .lcout(\c0.data_in_frame_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i233_LC_16_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i233_LC_16_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i233_LC_16_26_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i233_LC_16_26_4  (
            .in0(N__78654),
            .in1(N__59076),
            .in2(N__74456),
            .in3(N__80978),
            .lcout(\c0.data_in_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1926_LC_16_26_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1926_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1926_LC_16_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1926_LC_16_26_5  (
            .in0(N__59075),
            .in1(N__68619),
            .in2(_gnd_net_),
            .in3(N__66105),
            .lcout(\c0.n35181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1768_LC_16_26_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1768_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1768_LC_16_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1768_LC_16_26_6  (
            .in0(N__61720),
            .in1(N__59315),
            .in2(N__59061),
            .in3(N__59043),
            .lcout(\c0.n33374 ),
            .ltout(\c0.n33374_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1529_LC_16_26_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1529_LC_16_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1529_LC_16_26_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1529_LC_16_26_7  (
            .in0(N__66057),
            .in1(N__79576),
            .in2(N__59025),
            .in3(N__68910),
            .lcout(\c0.n33957 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i231_LC_16_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i231_LC_16_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i231_LC_16_27_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i231_LC_16_27_0  (
            .in0(N__79807),
            .in1(N__73920),
            .in2(N__59021),
            .in3(N__73577),
            .lcout(\c0.data_in_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97704),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_adj_1697_LC_16_27_1 .C_ON=1'b0;
    defparam \c0.i22_4_lut_adj_1697_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_adj_1697_LC_16_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_adj_1697_LC_16_27_1  (
            .in0(N__59001),
            .in1(N__65793),
            .in2(N__58992),
            .in3(N__58983),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1642_LC_16_27_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1642_LC_16_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1642_LC_16_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1642_LC_16_27_2  (
            .in0(N__74564),
            .in1(N__65601),
            .in2(N__73143),
            .in3(N__58977),
            .lcout(\c0.n16120 ),
            .ltout(\c0.n16120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1644_LC_16_27_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1644_LC_16_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1644_LC_16_27_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i2_3_lut_adj_1644_LC_16_27_3  (
            .in0(_gnd_net_),
            .in1(N__58971),
            .in2(N__58962),
            .in3(N__66173),
            .lcout(\c0.n33463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1534_LC_16_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1534_LC_16_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1534_LC_16_27_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1534_LC_16_27_4  (
            .in0(N__59367),
            .in1(N__61722),
            .in2(_gnd_net_),
            .in3(N__59316),
            .lcout(\c0.n31444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i194_LC_16_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i194_LC_16_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i194_LC_16_27_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i194_LC_16_27_5  (
            .in0(N__75339),
            .in1(N__81275),
            .in2(N__61670),
            .in3(N__79808),
            .lcout(\c0.data_in_frame_24_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97704),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1533_LC_16_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1533_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1533_LC_16_28_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1533_LC_16_28_0  (
            .in0(N__74760),
            .in1(N__79578),
            .in2(_gnd_net_),
            .in3(N__74790),
            .lcout(\c0.n33490 ),
            .ltout(\c0.n33490_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1699_LC_16_28_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1699_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1699_LC_16_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1699_LC_16_28_1  (
            .in0(N__59259),
            .in1(N__59253),
            .in2(N__59244),
            .in3(N__59241),
            .lcout(),
            .ltout(\c0.n25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1704_LC_16_28_2 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1704_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1704_LC_16_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_1704_LC_16_28_2  (
            .in0(N__61659),
            .in1(N__66075),
            .in2(N__59235),
            .in3(N__75392),
            .lcout(),
            .ltout(\c0.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1746_LC_16_28_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1746_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1746_LC_16_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_1746_LC_16_28_3  (
            .in0(N__62388),
            .in1(N__65910),
            .in2(N__59232),
            .in3(N__79377),
            .lcout(\c0.n33976 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1783_LC_16_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1783_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1783_LC_16_28_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1783_LC_16_28_5  (
            .in0(_gnd_net_),
            .in1(N__59229),
            .in2(_gnd_net_),
            .in3(N__59184),
            .lcout(\c0.n33969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1891_LC_16_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1891_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1891_LC_16_28_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1891_LC_16_28_6  (
            .in0(_gnd_net_),
            .in1(N__59150),
            .in2(_gnd_net_),
            .in3(N__61992),
            .lcout(\c0.n18228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1622_LC_16_29_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1622_LC_16_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1622_LC_16_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1622_LC_16_29_3  (
            .in0(N__68667),
            .in1(N__59108),
            .in2(N__68940),
            .in3(N__69158),
            .lcout(\c0.n20_adj_4656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23548_2_lut_LC_17_3_0 .C_ON=1'b0;
    defparam \quad_counter1.i23548_2_lut_LC_17_3_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23548_2_lut_LC_17_3_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23548_2_lut_LC_17_3_0  (
            .in0(_gnd_net_),
            .in1(N__81877),
            .in2(_gnd_net_),
            .in3(N__66345),
            .lcout(\quad_counter1.n28263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23543_2_lut_LC_17_4_0 .C_ON=1'b0;
    defparam \quad_counter1.i23543_2_lut_LC_17_4_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23543_2_lut_LC_17_4_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23543_2_lut_LC_17_4_0  (
            .in0(_gnd_net_),
            .in1(N__81928),
            .in2(_gnd_net_),
            .in3(N__66737),
            .lcout(),
            .ltout(\quad_counter1.n28257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1306_LC_17_4_1 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1306_LC_17_4_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1306_LC_17_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1306_LC_17_4_1  (
            .in0(N__66688),
            .in1(N__67063),
            .in2(N__59478),
            .in3(N__66710),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_adj_1307_LC_17_4_2 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_adj_1307_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_adj_1307_LC_17_4_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i3_4_lut_adj_1307_LC_17_4_2  (
            .in0(N__66640),
            .in1(N__66967),
            .in2(N__59475),
            .in3(N__66664),
            .lcout(\quad_counter1.n16_adj_4473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_17_4_6 .C_ON=1'b0;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.A_filtered_I_0_2_lut_LC_17_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter1.A_filtered_I_0_2_lut_LC_17_4_6  (
            .in0(_gnd_net_),
            .in1(N__59439),
            .in2(_gnd_net_),
            .in3(N__59468),
            .lcout(\quad_counter1.count_direction ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1085_1_lut_2_lut_LC_17_4_7 .C_ON=1'b0;
    defparam \quad_counter1.i1085_1_lut_2_lut_LC_17_4_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1085_1_lut_2_lut_LC_17_4_7 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \quad_counter1.i1085_1_lut_2_lut_LC_17_4_7  (
            .in0(N__59467),
            .in1(_gnd_net_),
            .in2(N__59447),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n2230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.B_delayed_77_LC_17_5_5 .C_ON=1'b0;
    defparam \quad_counter1.B_delayed_77_LC_17_5_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.B_delayed_77_LC_17_5_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \quad_counter1.B_delayed_77_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(N__59393),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.B_delayed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97537),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23648_2_lut_LC_17_7_4 .C_ON=1'b0;
    defparam \quad_counter0.i23648_2_lut_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23648_2_lut_LC_17_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23648_2_lut_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(N__63000),
            .in2(_gnd_net_),
            .in3(N__62957),
            .lcout(\quad_counter0.n28365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_adj_1324_LC_17_7_6 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_adj_1324_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_adj_1324_LC_17_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \quad_counter1.i3_4_lut_adj_1324_LC_17_7_6  (
            .in0(N__59472),
            .in1(N__59454),
            .in2(N__59448),
            .in3(N__59397),
            .lcout(count_enable_adj_4814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i0_LC_17_8_0 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i0_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i0_LC_17_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i0_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__59628),
            .in2(_gnd_net_),
            .in3(N__59616),
            .lcout(\quad_counter0.millisecond_counter_0 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\quad_counter0.n30140 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i1_LC_17_8_1 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i1_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i1_LC_17_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i1_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__59603),
            .in2(_gnd_net_),
            .in3(N__59592),
            .lcout(\quad_counter0.millisecond_counter_1 ),
            .ltout(),
            .carryin(\quad_counter0.n30140 ),
            .carryout(\quad_counter0.n30141 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i2_LC_17_8_2 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i2_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i2_LC_17_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i2_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__59589),
            .in2(_gnd_net_),
            .in3(N__59577),
            .lcout(\quad_counter0.millisecond_counter_2 ),
            .ltout(),
            .carryin(\quad_counter0.n30141 ),
            .carryout(\quad_counter0.n30142 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i3_LC_17_8_3 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i3_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i3_LC_17_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i3_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__59573),
            .in2(_gnd_net_),
            .in3(N__59559),
            .lcout(\quad_counter0.millisecond_counter_3 ),
            .ltout(),
            .carryin(\quad_counter0.n30142 ),
            .carryout(\quad_counter0.n30143 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i4_LC_17_8_4 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i4_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i4_LC_17_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i4_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__59556),
            .in2(_gnd_net_),
            .in3(N__59544),
            .lcout(\quad_counter0.millisecond_counter_4 ),
            .ltout(),
            .carryin(\quad_counter0.n30143 ),
            .carryout(\quad_counter0.n30144 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i5_LC_17_8_5 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i5_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i5_LC_17_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i5_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__59534),
            .in2(_gnd_net_),
            .in3(N__59523),
            .lcout(\quad_counter0.millisecond_counter_5 ),
            .ltout(),
            .carryin(\quad_counter0.n30144 ),
            .carryout(\quad_counter0.n30145 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i6_LC_17_8_6 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i6_LC_17_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i6_LC_17_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i6_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__59513),
            .in2(_gnd_net_),
            .in3(N__59502),
            .lcout(\quad_counter0.millisecond_counter_6 ),
            .ltout(),
            .carryin(\quad_counter0.n30145 ),
            .carryout(\quad_counter0.n30146 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i7_LC_17_8_7 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i7_LC_17_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i7_LC_17_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i7_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__59492),
            .in2(_gnd_net_),
            .in3(N__59481),
            .lcout(\quad_counter0.millisecond_counter_7 ),
            .ltout(),
            .carryin(\quad_counter0.n30146 ),
            .carryout(\quad_counter0.n30147 ),
            .clk(N__97539),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i8_LC_17_9_0 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i8_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i8_LC_17_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i8_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__59979),
            .in2(_gnd_net_),
            .in3(N__59952),
            .lcout(\quad_counter0.millisecond_counter_8 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\quad_counter0.n30148 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i9_LC_17_9_1 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i9_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i9_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i9_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__59946),
            .in2(_gnd_net_),
            .in3(N__59919),
            .lcout(\quad_counter0.millisecond_counter_9 ),
            .ltout(),
            .carryin(\quad_counter0.n30148 ),
            .carryout(\quad_counter0.n30149 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i10_LC_17_9_2 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i10_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i10_LC_17_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i10_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__59913),
            .in2(_gnd_net_),
            .in3(N__59886),
            .lcout(\quad_counter0.millisecond_counter_10 ),
            .ltout(),
            .carryin(\quad_counter0.n30149 ),
            .carryout(\quad_counter0.n30150 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i11_LC_17_9_3 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i11_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i11_LC_17_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i11_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__59880),
            .in2(_gnd_net_),
            .in3(N__59856),
            .lcout(\quad_counter0.millisecond_counter_11 ),
            .ltout(),
            .carryin(\quad_counter0.n30150 ),
            .carryout(\quad_counter0.n30151 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i12_LC_17_9_4 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i12_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i12_LC_17_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i12_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__59836),
            .in2(_gnd_net_),
            .in3(N__59814),
            .lcout(\quad_counter0.millisecond_counter_12 ),
            .ltout(),
            .carryin(\quad_counter0.n30151 ),
            .carryout(\quad_counter0.n30152 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i13_LC_17_9_5 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i13_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i13_LC_17_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i13_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__59794),
            .in2(_gnd_net_),
            .in3(N__59772),
            .lcout(\quad_counter0.millisecond_counter_13 ),
            .ltout(),
            .carryin(\quad_counter0.n30152 ),
            .carryout(\quad_counter0.n30153 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i14_LC_17_9_6 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i14_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i14_LC_17_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i14_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__59746),
            .in2(_gnd_net_),
            .in3(N__59724),
            .lcout(\quad_counter0.millisecond_counter_14 ),
            .ltout(),
            .carryin(\quad_counter0.n30153 ),
            .carryout(\quad_counter0.n30154 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i15_LC_17_9_7 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i15_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i15_LC_17_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i15_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__59695),
            .in2(_gnd_net_),
            .in3(N__59673),
            .lcout(\quad_counter0.millisecond_counter_15 ),
            .ltout(),
            .carryin(\quad_counter0.n30154 ),
            .carryout(\quad_counter0.n30155 ),
            .clk(N__97542),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i16_LC_17_10_0 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i16_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i16_LC_17_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i16_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__59661),
            .in2(_gnd_net_),
            .in3(N__59631),
            .lcout(\quad_counter0.millisecond_counter_16 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\quad_counter0.n30156 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i17_LC_17_10_1 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i17_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i17_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i17_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__60195),
            .in2(_gnd_net_),
            .in3(N__60162),
            .lcout(\quad_counter0.millisecond_counter_17 ),
            .ltout(),
            .carryin(\quad_counter0.n30156 ),
            .carryout(\quad_counter0.n30157 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i18_LC_17_10_2 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i18_LC_17_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i18_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i18_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__63921),
            .in2(_gnd_net_),
            .in3(N__60159),
            .lcout(\quad_counter0.millisecond_counter_18 ),
            .ltout(),
            .carryin(\quad_counter0.n30157 ),
            .carryout(\quad_counter0.n30158 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i19_LC_17_10_3 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i19_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i19_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i19_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__63688),
            .in2(_gnd_net_),
            .in3(N__60156),
            .lcout(\quad_counter0.millisecond_counter_19 ),
            .ltout(),
            .carryin(\quad_counter0.n30158 ),
            .carryout(\quad_counter0.n30159 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i20_LC_17_10_4 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i20_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i20_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i20_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__63053),
            .in2(_gnd_net_),
            .in3(N__60153),
            .lcout(\quad_counter0.millisecond_counter_20 ),
            .ltout(),
            .carryin(\quad_counter0.n30159 ),
            .carryout(\quad_counter0.n30160 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i21_LC_17_10_5 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i21_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i21_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i21_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__62999),
            .in2(_gnd_net_),
            .in3(N__60150),
            .lcout(\quad_counter0.millisecond_counter_21 ),
            .ltout(),
            .carryin(\quad_counter0.n30160 ),
            .carryout(\quad_counter0.n30161 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i22_LC_17_10_6 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i22_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i22_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i22_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__60135),
            .in2(_gnd_net_),
            .in3(N__60111),
            .lcout(\quad_counter0.millisecond_counter_22 ),
            .ltout(),
            .carryin(\quad_counter0.n30161 ),
            .carryout(\quad_counter0.n30162 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i23_LC_17_10_7 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i23_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i23_LC_17_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i23_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__60093),
            .in2(_gnd_net_),
            .in3(N__60066),
            .lcout(\quad_counter0.millisecond_counter_23 ),
            .ltout(),
            .carryin(\quad_counter0.n30162 ),
            .carryout(\quad_counter0.n30163 ),
            .clk(N__97545),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i24_LC_17_11_0 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i24_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i24_LC_17_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i24_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__60044),
            .in2(_gnd_net_),
            .in3(N__60030),
            .lcout(\quad_counter0.millisecond_counter_24 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\quad_counter0.n30164 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i25_LC_17_11_1 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i25_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i25_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i25_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__60007),
            .in2(_gnd_net_),
            .in3(N__60522),
            .lcout(\quad_counter0.millisecond_counter_25 ),
            .ltout(),
            .carryin(\quad_counter0.n30164 ),
            .carryout(\quad_counter0.n30165 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i26_LC_17_11_2 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i26_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i26_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i26_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__60502),
            .in2(_gnd_net_),
            .in3(N__60480),
            .lcout(\quad_counter0.millisecond_counter_26 ),
            .ltout(),
            .carryin(\quad_counter0.n30165 ),
            .carryout(\quad_counter0.n30166 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i27_LC_17_11_3 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i27_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i27_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i27_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__60457),
            .in2(_gnd_net_),
            .in3(N__60438),
            .lcout(\quad_counter0.millisecond_counter_27 ),
            .ltout(),
            .carryin(\quad_counter0.n30166 ),
            .carryout(\quad_counter0.n30167 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i28_LC_17_11_4 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i28_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i28_LC_17_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i28_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__60412),
            .in2(_gnd_net_),
            .in3(N__60396),
            .lcout(\quad_counter0.millisecond_counter_28 ),
            .ltout(),
            .carryin(\quad_counter0.n30167 ),
            .carryout(\quad_counter0.n30168 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i29_LC_17_11_5 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i29_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i29_LC_17_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i29_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__60372),
            .in2(_gnd_net_),
            .in3(N__60354),
            .lcout(\quad_counter0.millisecond_counter_29 ),
            .ltout(),
            .carryin(\quad_counter0.n30168 ),
            .carryout(\quad_counter0.n30169 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i30_LC_17_11_6 .C_ON=1'b1;
    defparam \quad_counter0.millisecond_counter_1425__i30_LC_17_11_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i30_LC_17_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i30_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__60331),
            .in2(_gnd_net_),
            .in3(N__60315),
            .lcout(\quad_counter0.millisecond_counter_30 ),
            .ltout(),
            .carryin(\quad_counter0.n30169 ),
            .carryout(\quad_counter0.n30170 ),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.millisecond_counter_1425__i31_LC_17_11_7 .C_ON=1'b0;
    defparam \quad_counter0.millisecond_counter_1425__i31_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.millisecond_counter_1425__i31_LC_17_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.millisecond_counter_1425__i31_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__60289),
            .in2(_gnd_net_),
            .in3(N__60312),
            .lcout(\quad_counter0.millisecond_counter_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97549),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_prev__i1_LC_17_12_5 .C_ON=1'b0;
    defparam \quad_counter0.count_prev__i1_LC_17_12_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_prev__i1_LC_17_12_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \quad_counter0.count_prev__i1_LC_17_12_5  (
            .in0(N__60248),
            .in1(N__85630),
            .in2(_gnd_net_),
            .in3(N__60272),
            .lcout(count_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97554),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_2_lut_LC_17_13_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_2_lut_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_2_lut_LC_17_13_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1750_2_lut_LC_17_13_0  (
            .in0(N__63926),
            .in1(N__63925),
            .in2(N__64447),
            .in3(N__60207),
            .lcout(\quad_counter0.n2619 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\quad_counter0.n30272 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_3_lut_LC_17_13_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_3_lut_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_3_lut_LC_17_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_3_lut_LC_17_13_1  (
            .in0(N__63894),
            .in1(N__63893),
            .in2(N__64511),
            .in3(N__60729),
            .lcout(\quad_counter0.n2618 ),
            .ltout(),
            .carryin(\quad_counter0.n30272 ),
            .carryout(\quad_counter0.n30273 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_4_lut_LC_17_13_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_4_lut_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_4_lut_LC_17_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1750_4_lut_LC_17_13_2  (
            .in0(N__64382),
            .in1(N__64381),
            .in2(N__64448),
            .in3(N__60699),
            .lcout(\quad_counter0.n2617 ),
            .ltout(),
            .carryin(\quad_counter0.n30273 ),
            .carryout(\quad_counter0.n30274 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_5_lut_LC_17_13_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_5_lut_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_5_lut_LC_17_13_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1750_5_lut_LC_17_13_3  (
            .in0(N__64405),
            .in1(N__64407),
            .in2(N__64451),
            .in3(N__60672),
            .lcout(\quad_counter0.n2616 ),
            .ltout(),
            .carryin(\quad_counter0.n30274 ),
            .carryout(\quad_counter0.n30275 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_6_lut_LC_17_13_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_6_lut_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_6_lut_LC_17_13_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1750_6_lut_LC_17_13_4  (
            .in0(N__64331),
            .in1(N__64330),
            .in2(N__64449),
            .in3(N__60642),
            .lcout(\quad_counter0.n2615 ),
            .ltout(),
            .carryin(\quad_counter0.n30275 ),
            .carryout(\quad_counter0.n30276 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_7_lut_LC_17_13_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_7_lut_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_7_lut_LC_17_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1750_7_lut_LC_17_13_5  (
            .in0(N__64310),
            .in1(N__64309),
            .in2(N__64452),
            .in3(N__60615),
            .lcout(\quad_counter0.n2614 ),
            .ltout(),
            .carryin(\quad_counter0.n30276 ),
            .carryout(\quad_counter0.n30277 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_8_lut_LC_17_13_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_8_lut_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_8_lut_LC_17_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1750_8_lut_LC_17_13_6  (
            .in0(N__64352),
            .in1(N__64351),
            .in2(N__64450),
            .in3(N__60582),
            .lcout(\quad_counter0.n2613 ),
            .ltout(),
            .carryin(\quad_counter0.n30277 ),
            .carryout(\quad_counter0.n30278 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_9_lut_LC_17_13_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_9_lut_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_9_lut_LC_17_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_9_lut_LC_17_13_7  (
            .in0(N__63876),
            .in1(N__63875),
            .in2(N__64512),
            .in3(N__60552),
            .lcout(\quad_counter0.n2612 ),
            .ltout(),
            .carryin(\quad_counter0.n30278 ),
            .carryout(\quad_counter0.n30279 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_10_lut_LC_17_14_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_10_lut_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_10_lut_LC_17_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_10_lut_LC_17_14_0  (
            .in0(N__63858),
            .in1(N__63857),
            .in2(N__64513),
            .in3(N__60525),
            .lcout(\quad_counter0.n2611 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\quad_counter0.n30280 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_11_lut_LC_17_14_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_11_lut_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_11_lut_LC_17_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_11_lut_LC_17_14_1  (
            .in0(N__63839),
            .in1(N__63838),
            .in2(N__64508),
            .in3(N__60885),
            .lcout(\quad_counter0.n2610 ),
            .ltout(),
            .carryin(\quad_counter0.n30280 ),
            .carryout(\quad_counter0.n30281 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_12_lut_LC_17_14_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_12_lut_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_12_lut_LC_17_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_12_lut_LC_17_14_2  (
            .in0(N__64287),
            .in1(N__64286),
            .in2(N__64514),
            .in3(N__60858),
            .lcout(\quad_counter0.n2609 ),
            .ltout(),
            .carryin(\quad_counter0.n30281 ),
            .carryout(\quad_counter0.n30282 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_13_lut_LC_17_14_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_13_lut_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_13_lut_LC_17_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_13_lut_LC_17_14_3  (
            .in0(N__63819),
            .in1(N__63818),
            .in2(N__64509),
            .in3(N__60831),
            .lcout(\quad_counter0.n2608 ),
            .ltout(),
            .carryin(\quad_counter0.n30282 ),
            .carryout(\quad_counter0.n30283 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_14_lut_LC_17_14_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1750_14_lut_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_14_lut_LC_17_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_14_lut_LC_17_14_4  (
            .in0(N__64560),
            .in1(N__64559),
            .in2(N__64515),
            .in3(N__60804),
            .lcout(\quad_counter0.n2607 ),
            .ltout(),
            .carryin(\quad_counter0.n30283 ),
            .carryout(\quad_counter0.n30284 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1750_15_lut_LC_17_14_5 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1750_15_lut_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1750_15_lut_LC_17_14_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1750_15_lut_LC_17_14_5  (
            .in0(N__64542),
            .in1(N__64541),
            .in2(N__64510),
            .in3(N__60801),
            .lcout(\quad_counter0.n2606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__3__5450_LC_17_15_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__3__5450_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__3__5450_LC_17_15_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_9__3__5450_LC_17_15_1  (
            .in0(N__60774),
            .in1(N__84637),
            .in2(N__85464),
            .in3(N__85227),
            .lcout(data_out_frame_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97572),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30749_LC_17_15_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30749_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30749_LC_17_15_3 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_30749_LC_17_15_3  (
            .in0(N__90320),
            .in1(N__81303),
            .in2(N__96176),
            .in3(N__60947),
            .lcout(),
            .ltout(\c0.n36161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36161_bdd_4_lut_LC_17_15_4 .C_ON=1'b0;
    defparam \c0.n36161_bdd_4_lut_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.n36161_bdd_4_lut_LC_17_15_4 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n36161_bdd_4_lut_LC_17_15_4  (
            .in0(N__60935),
            .in1(N__60773),
            .in2(N__60765),
            .in3(N__90321),
            .lcout(),
            .ltout(\c0.n36164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30654_4_lut_LC_17_15_5 .C_ON=1'b0;
    defparam \c0.i30654_4_lut_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30654_4_lut_LC_17_15_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.i30654_4_lut_LC_17_15_5  (
            .in0(N__90322),
            .in1(N__67524),
            .in2(N__60762),
            .in3(N__90027),
            .lcout(n36082),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__0__5437_LC_17_16_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__0__5437_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__0__5437_LC_17_16_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \c0.data_out_frame_11__0__5437_LC_17_16_0  (
            .in0(N__84617),
            .in1(N__61071),
            .in2(N__85233),
            .in3(N__79190),
            .lcout(data_out_frame_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__0__5445_LC_17_16_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__0__5445_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__0__5445_LC_17_16_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_10__0__5445_LC_17_16_3  (
            .in0(N__61059),
            .in1(N__84618),
            .in2(N__68037),
            .in3(N__85158),
            .lcout(data_out_frame_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30409_4_lut_LC_17_16_4 .C_ON=1'b0;
    defparam \c0.i30409_4_lut_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i30409_4_lut_LC_17_16_4 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \c0.i30409_4_lut_LC_17_16_4  (
            .in0(N__90039),
            .in1(N__60969),
            .in2(N__90375),
            .in3(N__60963),
            .lcout(),
            .ltout(\c0.n35836_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30411_4_lut_LC_17_16_5 .C_ON=1'b0;
    defparam \c0.i30411_4_lut_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30411_4_lut_LC_17_16_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.i30411_4_lut_LC_17_16_5  (
            .in0(N__90728),
            .in1(N__90884),
            .in2(N__60957),
            .in3(N__75957),
            .lcout(n35838),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__3__5442_LC_17_16_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__3__5442_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__3__5442_LC_17_16_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \c0.data_out_frame_10__3__5442_LC_17_16_6  (
            .in0(N__84616),
            .in1(N__60948),
            .in2(N__85232),
            .in3(N__77504),
            .lcout(data_out_frame_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97581),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__3__5458_LC_17_16_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__3__5458_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__3__5458_LC_17_16_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_8__3__5458_LC_17_16_7  (
            .in0(N__60936),
            .in1(N__84619),
            .in2(N__77145),
            .in3(N__85159),
            .lcout(data_out_frame_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97581),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i0_LC_17_17_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i0_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i0_LC_17_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i0_LC_17_17_0  (
            .in0(N__76520),
            .in1(N__64242),
            .in2(_gnd_net_),
            .in3(N__101270),
            .lcout(encoder1_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97587),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i19_LC_17_17_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i19_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i19_LC_17_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i19_LC_17_17_1  (
            .in0(N__76521),
            .in1(N__64614),
            .in2(_gnd_net_),
            .in3(N__83220),
            .lcout(encoder1_position_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__7__5422_LC_17_17_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__7__5422_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__7__5422_LC_17_17_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_12__7__5422_LC_17_17_2  (
            .in0(N__85197),
            .in1(N__84604),
            .in2(N__68184),
            .in3(N__60924),
            .lcout(data_out_frame_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30593_4_lut_LC_17_17_3 .C_ON=1'b0;
    defparam \c0.i30593_4_lut_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i30593_4_lut_LC_17_17_3 .LUT_INIT=16'b1100000001010000;
    LogicCell40 \c0.i30593_4_lut_LC_17_17_3  (
            .in0(N__90319),
            .in1(N__71718),
            .in2(N__96175),
            .in3(N__90046),
            .lcout(\c0.n36021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30769_LC_17_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30769_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30769_LC_17_17_4 .LUT_INIT=16'b1011110010110000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_30769_LC_17_17_4  (
            .in0(N__61070),
            .in1(N__90318),
            .in2(N__96174),
            .in3(N__61058),
            .lcout(\c0.n36197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__7__5414_LC_17_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__7__5414_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__7__5414_LC_17_17_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_13__7__5414_LC_17_17_6  (
            .in0(N__85198),
            .in1(N__61035),
            .in2(N__97962),
            .in3(N__84605),
            .lcout(data_out_frame_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97587),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i7_LC_17_17_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i7_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i7_LC_17_17_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i7_LC_17_17_7  (
            .in0(N__76522),
            .in1(N__64590),
            .in2(_gnd_net_),
            .in3(N__97951),
            .lcout(encoder1_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__6__5431_LC_17_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__6__5431_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__6__5431_LC_17_18_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_11__6__5431_LC_17_18_0  (
            .in0(N__61005),
            .in1(N__84690),
            .in2(N__85177),
            .in3(N__71890),
            .lcout(data_out_frame_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__6__5447_LC_17_18_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__6__5447_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__6__5447_LC_17_18_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.data_out_frame_9__6__5447_LC_17_18_1  (
            .in0(N__84689),
            .in1(N__85068),
            .in2(N__60996),
            .in3(N__75836),
            .lcout(data_out_frame_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30764_LC_17_18_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30764_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30764_LC_17_18_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_30764_LC_17_18_2  (
            .in0(N__61118),
            .in1(N__90317),
            .in2(N__67767),
            .in3(N__96055),
            .lcout(\c0.n36191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30759_LC_17_18_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30759_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30759_LC_17_18_3 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_30759_LC_17_18_3  (
            .in0(N__90315),
            .in1(N__61016),
            .in2(N__96123),
            .in3(N__61004),
            .lcout(),
            .ltout(\c0.n36185_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36185_bdd_4_lut_LC_17_18_4 .C_ON=1'b0;
    defparam \c0.n36185_bdd_4_lut_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.n36185_bdd_4_lut_LC_17_18_4 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n36185_bdd_4_lut_LC_17_18_4  (
            .in0(N__61395),
            .in1(N__60992),
            .in2(N__60984),
            .in3(N__90316),
            .lcout(\c0.n36188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__1__5452_LC_17_18_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__1__5452_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__1__5452_LC_17_18_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_9__1__5452_LC_17_18_5  (
            .in0(N__84688),
            .in1(N__85067),
            .in2(N__71808),
            .in3(N__61247),
            .lcout(data_out_frame_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1980_LC_17_18_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1980_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1980_LC_17_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1980_LC_17_18_6  (
            .in0(N__67893),
            .in1(N__61233),
            .in2(_gnd_net_),
            .in3(N__61215),
            .lcout(\c0.n18479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__5__5480_LC_17_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__5__5480_LC_17_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__5__5480_LC_17_18_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__5__5480_LC_17_18_7  (
            .in0(N__84687),
            .in1(N__85066),
            .in2(N__76815),
            .in3(N__61107),
            .lcout(data_out_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97596),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i10_LC_17_19_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i10_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i10_LC_17_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i10_LC_17_19_1  (
            .in0(N__76562),
            .in1(N__64575),
            .in2(_gnd_net_),
            .in3(N__83117),
            .lcout(encoder1_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__5__5432_LC_17_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__5__5432_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__5__5432_LC_17_19_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_11__5__5432_LC_17_19_2  (
            .in0(N__85203),
            .in1(N__84684),
            .in2(N__85515),
            .in3(N__67463),
            .lcout(data_out_frame_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__7__5430_LC_17_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__7__5430_LC_17_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__7__5430_LC_17_19_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_11__7__5430_LC_17_19_4  (
            .in0(N__85204),
            .in1(N__61122),
            .in2(N__67871),
            .in3(N__84686),
            .lcout(data_out_frame_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97606),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i23_LC_17_19_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i23_LC_17_19_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i23_LC_17_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i23_LC_17_19_5  (
            .in0(N__76563),
            .in1(N__64671),
            .in2(_gnd_net_),
            .in3(N__67866),
            .lcout(encoder1_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__7__5462_LC_17_19_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__7__5462_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__7__5462_LC_17_19_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_7__7__5462_LC_17_19_6  (
            .in0(N__85205),
            .in1(N__84685),
            .in2(N__72600),
            .in3(N__71918),
            .lcout(data_out_frame_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30657_4_lut_LC_17_19_7 .C_ON=1'b0;
    defparam \c0.i30657_4_lut_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30657_4_lut_LC_17_19_7 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \c0.i30657_4_lut_LC_17_19_7  (
            .in0(N__90064),
            .in1(N__96135),
            .in2(N__90391),
            .in3(N__61106),
            .lcout(\c0.n36086 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__2__5467_LC_17_20_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__2__5467_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__2__5467_LC_17_20_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_7__2__5467_LC_17_20_0  (
            .in0(N__85210),
            .in1(N__84682),
            .in2(N__77700),
            .in3(N__61091),
            .lcout(data_out_frame_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_17_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_17_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_17_20_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i53_LC_17_20_1  (
            .in0(N__89795),
            .in1(N__83699),
            .in2(N__61340),
            .in3(N__84231),
            .lcout(\c0.data_in_frame_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__5__5472_LC_17_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__5__5472_LC_17_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__5__5472_LC_17_20_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_6__5__5472_LC_17_20_2  (
            .in0(N__61320),
            .in1(N__84680),
            .in2(N__85252),
            .in3(N__79060),
            .lcout(data_out_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__5__5464_LC_17_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__5__5464_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__5__5464_LC_17_20_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.data_out_frame_7__5__5464_LC_17_20_3  (
            .in0(N__84679),
            .in1(N__85211),
            .in2(N__61308),
            .in3(N__61617),
            .lcout(data_out_frame_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_17_20_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_17_20_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_17_20_4  (
            .in0(N__61319),
            .in1(N__96122),
            .in2(_gnd_net_),
            .in3(N__61304),
            .lcout(),
            .ltout(\c0.n5_adj_4619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30394_4_lut_LC_17_20_5 .C_ON=1'b0;
    defparam \c0.i30394_4_lut_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30394_4_lut_LC_17_20_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.i30394_4_lut_LC_17_20_5  (
            .in0(N__61296),
            .in1(N__90396),
            .in2(N__61290),
            .in3(N__90084),
            .lcout(\c0.n35821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__6__5471_LC_17_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__6__5471_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__6__5471_LC_17_20_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_6__6__5471_LC_17_20_6  (
            .in0(N__85209),
            .in1(N__84681),
            .in2(N__76860),
            .in3(N__61286),
            .lcout(data_out_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1444_LC_17_20_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1444_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1444_LC_17_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1444_LC_17_20_7  (
            .in0(N__61616),
            .in1(N__72062),
            .in2(_gnd_net_),
            .in3(N__76807),
            .lcout(\c0.n18124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__4__5441_LC_17_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__4__5441_LC_17_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__4__5441_LC_17_21_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_10__4__5441_LC_17_21_0  (
            .in0(N__85212),
            .in1(N__84669),
            .in2(N__77352),
            .in3(N__65205),
            .lcout(data_out_frame_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30397_4_lut_LC_17_21_1 .C_ON=1'b0;
    defparam \c0.i30397_4_lut_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i30397_4_lut_LC_17_21_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \c0.i30397_4_lut_LC_17_21_1  (
            .in0(N__90086),
            .in1(N__61272),
            .in2(N__90395),
            .in3(N__61263),
            .lcout(\c0.n35824 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__4__5465_LC_17_21_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__4__5465_LC_17_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__4__5465_LC_17_21_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_7__4__5465_LC_17_21_2  (
            .in0(N__85214),
            .in1(N__84670),
            .in2(N__72004),
            .in3(N__65037),
            .lcout(data_out_frame_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_17_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_17_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_17_21_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i8_LC_17_21_3  (
            .in0(N__81270),
            .in1(N__83698),
            .in2(N__61437),
            .in3(N__79998),
            .lcout(\c0.data_in_frame_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__6__5455_LC_17_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__6__5455_LC_17_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__6__5455_LC_17_21_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.data_out_frame_8__6__5455_LC_17_21_5  (
            .in0(N__61391),
            .in1(N__85787),
            .in2(N__84716),
            .in3(N__85216),
            .lcout(data_out_frame_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__6__5479_LC_17_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__6__5479_LC_17_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__6__5479_LC_17_21_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_5__6__5479_LC_17_21_6  (
            .in0(N__85213),
            .in1(N__61376),
            .in2(N__72661),
            .in3(N__84677),
            .lcout(data_out_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97631),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__4__5433_LC_17_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__4__5433_LC_17_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__4__5433_LC_17_21_7 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \c0.data_out_frame_11__4__5433_LC_17_21_7  (
            .in0(N__76662),
            .in1(N__65217),
            .in2(N__84717),
            .in3(N__85215),
            .lcout(data_out_frame_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97631),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_1_LC_17_22_0 .C_ON=1'b1;
    defparam \quad_counter0.add_657_1_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_1_LC_17_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter0.add_657_1_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__61845),
            .in2(N__61917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\quad_counter0.n30108 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_2_lut_LC_17_22_1 .C_ON=1'b1;
    defparam \quad_counter0.add_657_2_lut_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_2_lut_LC_17_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_2_lut_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__61362),
            .in2(N__85603),
            .in3(N__61350),
            .lcout(n2345),
            .ltout(),
            .carryin(\quad_counter0.n30108 ),
            .carryout(\quad_counter0.n30109 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_3_lut_LC_17_22_2 .C_ON=1'b1;
    defparam \quad_counter0.add_657_3_lut_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_3_lut_LC_17_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_3_lut_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__61846),
            .in2(N__71804),
            .in3(N__61347),
            .lcout(n2344),
            .ltout(),
            .carryin(\quad_counter0.n30109 ),
            .carryout(\quad_counter0.n30110 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_4_lut_LC_17_22_3 .C_ON=1'b1;
    defparam \quad_counter0.add_657_4_lut_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_4_lut_LC_17_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_4_lut_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__83320),
            .in2(N__61914),
            .in3(N__61344),
            .lcout(n2343),
            .ltout(),
            .carryin(\quad_counter0.n30110 ),
            .carryout(\quad_counter0.n30111 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_5_lut_LC_17_22_4 .C_ON=1'b1;
    defparam \quad_counter0.add_657_5_lut_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_5_lut_LC_17_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_5_lut_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(N__61850),
            .in2(N__85451),
            .in3(N__61485),
            .lcout(n2342),
            .ltout(),
            .carryin(\quad_counter0.n30111 ),
            .carryout(\quad_counter0.n30112 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_6_lut_LC_17_22_5 .C_ON=1'b1;
    defparam \quad_counter0.add_657_6_lut_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_6_lut_LC_17_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_6_lut_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__85378),
            .in2(N__61915),
            .in3(N__61482),
            .lcout(n2341),
            .ltout(),
            .carryin(\quad_counter0.n30112 ),
            .carryout(\quad_counter0.n30113 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_7_lut_LC_17_22_6 .C_ON=1'b1;
    defparam \quad_counter0.add_657_7_lut_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_7_lut_LC_17_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_7_lut_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__61854),
            .in2(N__96638),
            .in3(N__61479),
            .lcout(n2340),
            .ltout(),
            .carryin(\quad_counter0.n30113 ),
            .carryout(\quad_counter0.n30114 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_8_lut_LC_17_22_7 .C_ON=1'b1;
    defparam \quad_counter0.add_657_8_lut_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_8_lut_LC_17_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_8_lut_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(N__75824),
            .in2(N__61916),
            .in3(N__61476),
            .lcout(n2339),
            .ltout(),
            .carryin(\quad_counter0.n30114 ),
            .carryout(\quad_counter0.n30115 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_9_lut_LC_17_23_0 .C_ON=1'b1;
    defparam \quad_counter0.add_657_9_lut_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_9_lut_LC_17_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_9_lut_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__61861),
            .in2(N__75944),
            .in3(N__61473),
            .lcout(n2338),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\quad_counter0.n30116 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_10_lut_LC_17_23_1 .C_ON=1'b1;
    defparam \quad_counter0.add_657_10_lut_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_10_lut_LC_17_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_10_lut_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__73232),
            .in2(N__61918),
            .in3(N__61470),
            .lcout(n2337),
            .ltout(),
            .carryin(\quad_counter0.n30116 ),
            .carryout(\quad_counter0.n30117 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_11_lut_LC_17_23_2 .C_ON=1'b1;
    defparam \quad_counter0.add_657_11_lut_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_11_lut_LC_17_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_11_lut_LC_17_23_2  (
            .in0(_gnd_net_),
            .in1(N__61865),
            .in2(N__77453),
            .in3(N__61467),
            .lcout(n2336),
            .ltout(),
            .carryin(\quad_counter0.n30117 ),
            .carryout(\quad_counter0.n30118 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_12_lut_LC_17_23_3 .C_ON=1'b1;
    defparam \quad_counter0.add_657_12_lut_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_12_lut_LC_17_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_12_lut_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__72380),
            .in2(N__61919),
            .in3(N__61464),
            .lcout(n2335),
            .ltout(),
            .carryin(\quad_counter0.n30118 ),
            .carryout(\quad_counter0.n30119 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_13_lut_LC_17_23_4 .C_ON=1'b1;
    defparam \quad_counter0.add_657_13_lut_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_13_lut_LC_17_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_13_lut_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(N__61869),
            .in2(N__77141),
            .in3(N__61461),
            .lcout(n2334),
            .ltout(),
            .carryin(\quad_counter0.n30119 ),
            .carryout(\quad_counter0.n30120 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_14_lut_LC_17_23_5 .C_ON=1'b1;
    defparam \quad_counter0.add_657_14_lut_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_14_lut_LC_17_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_14_lut_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__79244),
            .in2(N__61920),
            .in3(N__61524),
            .lcout(n2333),
            .ltout(),
            .carryin(\quad_counter0.n30120 ),
            .carryout(\quad_counter0.n30121 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_15_lut_LC_17_23_6 .C_ON=1'b1;
    defparam \quad_counter0.add_657_15_lut_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_15_lut_LC_17_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_15_lut_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(N__61873),
            .in2(N__77826),
            .in3(N__61521),
            .lcout(n2332),
            .ltout(),
            .carryin(\quad_counter0.n30121 ),
            .carryout(\quad_counter0.n30122 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_16_lut_LC_17_23_7 .C_ON=1'b1;
    defparam \quad_counter0.add_657_16_lut_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_16_lut_LC_17_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_16_lut_LC_17_23_7  (
            .in0(_gnd_net_),
            .in1(N__85777),
            .in2(N__61921),
            .in3(N__61518),
            .lcout(n2331),
            .ltout(),
            .carryin(\quad_counter0.n30122 ),
            .carryout(\quad_counter0.n30123 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_17_lut_LC_17_24_0 .C_ON=1'b1;
    defparam \quad_counter0.add_657_17_lut_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_17_lut_LC_17_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_17_lut_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(N__86495),
            .in2(N__61955),
            .in3(N__61515),
            .lcout(n2330),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\quad_counter0.n30124 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_18_lut_LC_17_24_1 .C_ON=1'b1;
    defparam \quad_counter0.add_657_18_lut_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_18_lut_LC_17_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_18_lut_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__61925),
            .in2(N__86426),
            .in3(N__61512),
            .lcout(n2329),
            .ltout(),
            .carryin(\quad_counter0.n30124 ),
            .carryout(\quad_counter0.n30125 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_19_lut_LC_17_24_2 .C_ON=1'b1;
    defparam \quad_counter0.add_657_19_lut_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_19_lut_LC_17_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_19_lut_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__83279),
            .in2(N__61956),
            .in3(N__61509),
            .lcout(n2328),
            .ltout(),
            .carryin(\quad_counter0.n30125 ),
            .carryout(\quad_counter0.n30126 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_20_lut_LC_17_24_3 .C_ON=1'b1;
    defparam \quad_counter0.add_657_20_lut_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_20_lut_LC_17_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_20_lut_LC_17_24_3  (
            .in0(_gnd_net_),
            .in1(N__61929),
            .in2(N__77699),
            .in3(N__61506),
            .lcout(n2327),
            .ltout(),
            .carryin(\quad_counter0.n30126 ),
            .carryout(\quad_counter0.n30127 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_21_lut_LC_17_24_4 .C_ON=1'b1;
    defparam \quad_counter0.add_657_21_lut_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_21_lut_LC_17_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_21_lut_LC_17_24_4  (
            .in0(_gnd_net_),
            .in1(N__72069),
            .in2(N__61957),
            .in3(N__61491),
            .lcout(n2326),
            .ltout(),
            .carryin(\quad_counter0.n30127 ),
            .carryout(\quad_counter0.n30128 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_22_lut_LC_17_24_5 .C_ON=1'b1;
    defparam \quad_counter0.add_657_22_lut_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_22_lut_LC_17_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_22_lut_LC_17_24_5  (
            .in0(_gnd_net_),
            .in1(N__61933),
            .in2(N__72008),
            .in3(N__61488),
            .lcout(n2325),
            .ltout(),
            .carryin(\quad_counter0.n30128 ),
            .carryout(\quad_counter0.n30129 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_23_lut_LC_17_24_6 .C_ON=1'b1;
    defparam \quad_counter0.add_657_23_lut_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_23_lut_LC_17_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_23_lut_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(N__61615),
            .in2(N__61958),
            .in3(N__61581),
            .lcout(n2324),
            .ltout(),
            .carryin(\quad_counter0.n30129 ),
            .carryout(\quad_counter0.n30130 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_24_lut_LC_17_24_7 .C_ON=1'b1;
    defparam \quad_counter0.add_657_24_lut_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_24_lut_LC_17_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_24_lut_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__61937),
            .in2(N__76752),
            .in3(N__61566),
            .lcout(n2323),
            .ltout(),
            .carryin(\quad_counter0.n30130 ),
            .carryout(\quad_counter0.n30131 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_25_lut_LC_17_25_0 .C_ON=1'b1;
    defparam \quad_counter0.add_657_25_lut_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_25_lut_LC_17_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_25_lut_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__61938),
            .in2(N__72596),
            .in3(N__61563),
            .lcout(n2322),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\quad_counter0.n30132 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_26_lut_LC_17_25_1 .C_ON=1'b1;
    defparam \quad_counter0.add_657_26_lut_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_26_lut_LC_17_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_26_lut_LC_17_25_1  (
            .in0(_gnd_net_),
            .in1(N__78035),
            .in2(N__61959),
            .in3(N__61560),
            .lcout(n2321),
            .ltout(),
            .carryin(\quad_counter0.n30132 ),
            .carryout(\quad_counter0.n30133 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_27_lut_LC_17_25_2 .C_ON=1'b1;
    defparam \quad_counter0.add_657_27_lut_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_27_lut_LC_17_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_27_lut_LC_17_25_2  (
            .in0(_gnd_net_),
            .in1(N__61942),
            .in2(N__73097),
            .in3(N__61557),
            .lcout(n2320),
            .ltout(),
            .carryin(\quad_counter0.n30133 ),
            .carryout(\quad_counter0.n30134 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_28_lut_LC_17_25_3 .C_ON=1'b1;
    defparam \quad_counter0.add_657_28_lut_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_28_lut_LC_17_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_28_lut_LC_17_25_3  (
            .in0(_gnd_net_),
            .in1(N__85920),
            .in2(N__61960),
            .in3(N__61554),
            .lcout(n2319),
            .ltout(),
            .carryin(\quad_counter0.n30134 ),
            .carryout(\quad_counter0.n30135 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_29_lut_LC_17_25_4 .C_ON=1'b1;
    defparam \quad_counter0.add_657_29_lut_LC_17_25_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_29_lut_LC_17_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_29_lut_LC_17_25_4  (
            .in0(_gnd_net_),
            .in1(N__61946),
            .in2(N__79146),
            .in3(N__61545),
            .lcout(n2318),
            .ltout(),
            .carryin(\quad_counter0.n30135 ),
            .carryout(\quad_counter0.n30136 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_30_lut_LC_17_25_5 .C_ON=1'b1;
    defparam \quad_counter0.add_657_30_lut_LC_17_25_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_30_lut_LC_17_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_30_lut_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(N__86198),
            .in2(N__61961),
            .in3(N__61542),
            .lcout(n2317),
            .ltout(),
            .carryin(\quad_counter0.n30136 ),
            .carryout(\quad_counter0.n30137 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_31_lut_LC_17_25_6 .C_ON=1'b1;
    defparam \quad_counter0.add_657_31_lut_LC_17_25_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_31_lut_LC_17_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_31_lut_LC_17_25_6  (
            .in0(_gnd_net_),
            .in1(N__61950),
            .in2(N__79070),
            .in3(N__61527),
            .lcout(n2316),
            .ltout(),
            .carryin(\quad_counter0.n30137 ),
            .carryout(\quad_counter0.n30138 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_32_lut_LC_17_25_7 .C_ON=1'b1;
    defparam \quad_counter0.add_657_32_lut_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_32_lut_LC_17_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.add_657_32_lut_LC_17_25_7  (
            .in0(_gnd_net_),
            .in1(N__76846),
            .in2(N__61962),
            .in3(N__61965),
            .lcout(n2315),
            .ltout(),
            .carryin(\quad_counter0.n30138 ),
            .carryout(\quad_counter0.n30139 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.add_657_33_lut_LC_17_26_0 .C_ON=1'b0;
    defparam \quad_counter0.add_657_33_lut_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.add_657_33_lut_LC_17_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.add_657_33_lut_LC_17_26_0  (
            .in0(N__61954),
            .in1(N__76910),
            .in2(_gnd_net_),
            .in3(N__61776),
            .lcout(n2314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1933_LC_17_26_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1933_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1933_LC_17_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1933_LC_17_26_1  (
            .in0(N__61773),
            .in1(N__74004),
            .in2(N__62040),
            .in3(N__74187),
            .lcout(\c0.n34841 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1640_LC_17_26_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1640_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1640_LC_17_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1640_LC_17_26_3  (
            .in0(N__65891),
            .in1(N__65549),
            .in2(N__61755),
            .in3(N__61739),
            .lcout(\c0.n31451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1680_LC_17_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1680_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1680_LC_17_26_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1680_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__61719),
            .in2(_gnd_net_),
            .in3(N__61698),
            .lcout(\c0.n33948 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1909_LC_17_26_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1909_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1909_LC_17_26_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1909_LC_17_26_5  (
            .in0(_gnd_net_),
            .in1(N__68473),
            .in2(_gnd_net_),
            .in3(N__68663),
            .lcout(\c0.n18193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i237_LC_17_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i237_LC_17_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i237_LC_17_26_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i237_LC_17_26_7  (
            .in0(N__74445),
            .in1(N__84240),
            .in2(N__62345),
            .in3(N__78557),
            .lcout(\c0.data_in_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_13_2_lut_LC_17_27_0 .C_ON=1'b0;
    defparam \c0.i1_rep_13_2_lut_LC_17_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_13_2_lut_LC_17_27_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_rep_13_2_lut_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(N__61663),
            .in2(_gnd_net_),
            .in3(N__66079),
            .lcout(),
            .ltout(\c0.n36530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1923_LC_17_27_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1923_LC_17_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1923_LC_17_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1923_LC_17_27_1  (
            .in0(N__67944),
            .in1(N__61638),
            .in2(N__61620),
            .in3(N__68991),
            .lcout(\c0.n10_adj_4755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1632_LC_17_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1632_LC_17_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1632_LC_17_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1632_LC_17_27_2  (
            .in0(_gnd_net_),
            .in1(N__74522),
            .in2(_gnd_net_),
            .in3(N__66183),
            .lcout(\c0.n32431 ),
            .ltout(\c0.n32431_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1924_LC_17_27_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1924_LC_17_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1924_LC_17_27_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1924_LC_17_27_3  (
            .in0(N__66134),
            .in1(N__74474),
            .in2(N__62355),
            .in3(N__69138),
            .lcout(\c0.n35142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1928_LC_17_27_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1928_LC_17_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1928_LC_17_27_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1928_LC_17_27_5  (
            .in0(N__68825),
            .in1(N__62352),
            .in2(N__62346),
            .in3(N__69350),
            .lcout(\c0.n35314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i196_LC_17_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i196_LC_17_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i196_LC_17_27_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i196_LC_17_27_7  (
            .in0(N__78979),
            .in1(N__81172),
            .in2(N__66084),
            .in3(N__79844),
            .lcout(\c0.data_in_frame_24_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i140_LC_17_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i140_LC_17_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i140_LC_17_28_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i140_LC_17_28_0  (
            .in0(N__87298),
            .in1(N__73011),
            .in2(N__62309),
            .in3(N__78980),
            .lcout(\c0.data_in_frame_17_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1906_LC_17_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1906_LC_17_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1906_LC_17_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1906_LC_17_28_1  (
            .in0(_gnd_net_),
            .in1(N__62025),
            .in2(_gnd_net_),
            .in3(N__65722),
            .lcout(\c0.n18405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i190_LC_17_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i190_LC_17_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i190_LC_17_28_2 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \c0.data_in_frame_0__i190_LC_17_28_2  (
            .in0(N__75066),
            .in1(N__73012),
            .in2(N__62267),
            .in3(N__65735),
            .lcout(\c0.data_in_frame_23_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i189_LC_17_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i189_LC_17_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i189_LC_17_28_3 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_in_frame_0__i189_LC_17_28_3  (
            .in0(N__73009),
            .in1(N__62026),
            .in2(N__62268),
            .in3(N__84243),
            .lcout(\c0.data_in_frame_23_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i133_LC_17_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i133_LC_17_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i133_LC_17_28_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i133_LC_17_28_4  (
            .in0(N__84241),
            .in1(N__73010),
            .in2(N__62003),
            .in3(N__81173),
            .lcout(\c0.data_in_frame_16_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i149_LC_17_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i149_LC_17_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i149_LC_17_28_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i149_LC_17_28_5  (
            .in0(N__73008),
            .in1(N__84242),
            .in2(N__80412),
            .in3(N__62431),
            .lcout(\c0.data_in_frame_18_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97744),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1624_LC_17_28_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1624_LC_17_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1624_LC_17_28_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i9_4_lut_adj_1624_LC_17_28_6  (
            .in0(N__69212),
            .in1(N__68322),
            .in2(N__79632),
            .in3(N__73403),
            .lcout(\c0.n21_adj_4659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_1736_LC_17_28_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_1736_LC_17_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_1736_LC_17_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_1736_LC_17_28_7  (
            .in0(N__68972),
            .in1(N__68688),
            .in2(N__65412),
            .in3(N__62415),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i8_4_lut_adj_1288_LC_18_2_0 .C_ON=1'b0;
    defparam \quad_counter1.i8_4_lut_adj_1288_LC_18_2_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i8_4_lut_adj_1288_LC_18_2_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i8_4_lut_adj_1288_LC_18_2_0  (
            .in0(N__66466),
            .in1(N__66424),
            .in2(N__66624),
            .in3(N__66549),
            .lcout(\quad_counter1.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1291_LC_18_2_1 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1291_LC_18_2_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1291_LC_18_2_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1291_LC_18_2_1  (
            .in0(N__62361),
            .in1(N__66568),
            .in2(N__66520),
            .in3(N__62694),
            .lcout(\quad_counter1.n2936 ),
            .ltout(\quad_counter1.n2936_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30732_1_lut_LC_18_2_2 .C_ON=1'b0;
    defparam \quad_counter1.i30732_1_lut_LC_18_2_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30732_1_lut_LC_18_2_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30732_1_lut_LC_18_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62382),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1287_LC_18_2_3 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1287_LC_18_2_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1287_LC_18_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1287_LC_18_2_3  (
            .in0(N__62379),
            .in1(N__66220),
            .in2(N__66313),
            .in3(N__66283),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4458_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_4_lut_adj_1289_LC_18_2_4 .C_ON=1'b0;
    defparam \quad_counter1.i1_4_lut_adj_1289_LC_18_2_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_4_lut_adj_1289_LC_18_2_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i1_4_lut_adj_1289_LC_18_2_4  (
            .in0(N__66262),
            .in1(N__66445),
            .in2(N__62373),
            .in3(N__66241),
            .lcout(),
            .ltout(\quad_counter1.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1290_LC_18_2_5 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1290_LC_18_2_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1290_LC_18_2_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1290_LC_18_2_5  (
            .in0(N__62370),
            .in1(N__66774),
            .in2(N__62364),
            .in3(N__66586),
            .lcout(\quad_counter1.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_2_lut_LC_18_3_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_2_lut_LC_18_3_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_2_lut_LC_18_3_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2018_2_lut_LC_18_3_0  (
            .in0(N__81879),
            .in1(N__81878),
            .in2(N__62494),
            .in3(N__62523),
            .lcout(\quad_counter1.n3019 ),
            .ltout(),
            .carryin(bfn_18_3_0_),
            .carryout(\quad_counter1.n30580 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_3_lut_LC_18_3_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_3_lut_LC_18_3_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_3_lut_LC_18_3_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_3_lut_LC_18_3_1  (
            .in0(N__66341),
            .in1(N__66340),
            .in2(N__62572),
            .in3(N__62520),
            .lcout(\quad_counter1.n3018 ),
            .ltout(),
            .carryin(\quad_counter1.n30580 ),
            .carryout(\quad_counter1.n30581 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_4_lut_LC_18_3_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_4_lut_LC_18_3_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_4_lut_LC_18_3_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2018_4_lut_LC_18_3_2  (
            .in0(N__66317),
            .in1(N__66318),
            .in2(N__62495),
            .in3(N__62517),
            .lcout(\quad_counter1.n3017 ),
            .ltout(),
            .carryin(\quad_counter1.n30581 ),
            .carryout(\quad_counter1.n30582 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_5_lut_LC_18_3_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_5_lut_LC_18_3_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_5_lut_LC_18_3_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2018_5_lut_LC_18_3_3  (
            .in0(N__66287),
            .in1(N__66288),
            .in2(N__62504),
            .in3(N__62514),
            .lcout(\quad_counter1.n3016 ),
            .ltout(),
            .carryin(\quad_counter1.n30582 ),
            .carryout(\quad_counter1.n30583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_6_lut_LC_18_3_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_6_lut_LC_18_3_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_6_lut_LC_18_3_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2018_6_lut_LC_18_3_4  (
            .in0(N__66264),
            .in1(N__66263),
            .in2(N__62496),
            .in3(N__62511),
            .lcout(\quad_counter1.n3015 ),
            .ltout(),
            .carryin(\quad_counter1.n30583 ),
            .carryout(\quad_counter1.n30584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_7_lut_LC_18_3_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_7_lut_LC_18_3_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_7_lut_LC_18_3_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2018_7_lut_LC_18_3_5  (
            .in0(N__66243),
            .in1(N__66242),
            .in2(N__62505),
            .in3(N__62508),
            .lcout(\quad_counter1.n3014 ),
            .ltout(),
            .carryin(\quad_counter1.n30584 ),
            .carryout(\quad_counter1.n30585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_8_lut_LC_18_3_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_8_lut_LC_18_3_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_8_lut_LC_18_3_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2018_8_lut_LC_18_3_6  (
            .in0(N__66222),
            .in1(N__66221),
            .in2(N__62497),
            .in3(N__62460),
            .lcout(\quad_counter1.n3013 ),
            .ltout(),
            .carryin(\quad_counter1.n30585 ),
            .carryout(\quad_counter1.n30586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_9_lut_LC_18_3_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_9_lut_LC_18_3_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_9_lut_LC_18_3_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_9_lut_LC_18_3_7  (
            .in0(N__66623),
            .in1(N__66622),
            .in2(N__62573),
            .in3(N__62457),
            .lcout(\quad_counter1.n3012 ),
            .ltout(),
            .carryin(\quad_counter1.n30586 ),
            .carryout(\quad_counter1.n30587 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_10_lut_LC_18_4_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_10_lut_LC_18_4_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_10_lut_LC_18_4_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_10_lut_LC_18_4_0  (
            .in0(N__66600),
            .in1(N__66593),
            .in2(N__62604),
            .in3(N__62454),
            .lcout(\quad_counter1.n3011 ),
            .ltout(),
            .carryin(bfn_18_4_0_),
            .carryout(\quad_counter1.n30588 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_11_lut_LC_18_4_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_11_lut_LC_18_4_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_11_lut_LC_18_4_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_11_lut_LC_18_4_1  (
            .in0(N__66570),
            .in1(N__66569),
            .in2(N__62608),
            .in3(N__62643),
            .lcout(\quad_counter1.n3010 ),
            .ltout(),
            .carryin(\quad_counter1.n30588 ),
            .carryout(\quad_counter1.n30589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_12_lut_LC_18_4_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_12_lut_LC_18_4_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_12_lut_LC_18_4_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_12_lut_LC_18_4_2  (
            .in0(N__66548),
            .in1(N__66547),
            .in2(N__62605),
            .in3(N__62640),
            .lcout(\quad_counter1.n3009 ),
            .ltout(),
            .carryin(\quad_counter1.n30589 ),
            .carryout(\quad_counter1.n30590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_13_lut_LC_18_4_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_13_lut_LC_18_4_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_13_lut_LC_18_4_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_13_lut_LC_18_4_3  (
            .in0(N__66524),
            .in1(N__66525),
            .in2(N__62609),
            .in3(N__62637),
            .lcout(\quad_counter1.n3008 ),
            .ltout(),
            .carryin(\quad_counter1.n30590 ),
            .carryout(\quad_counter1.n30591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_14_lut_LC_18_4_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_14_lut_LC_18_4_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_14_lut_LC_18_4_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_14_lut_LC_18_4_4  (
            .in0(N__66491),
            .in1(N__66490),
            .in2(N__62606),
            .in3(N__62634),
            .lcout(\quad_counter1.n3007 ),
            .ltout(),
            .carryin(\quad_counter1.n30591 ),
            .carryout(\quad_counter1.n30592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_15_lut_LC_18_4_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_15_lut_LC_18_4_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_15_lut_LC_18_4_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_15_lut_LC_18_4_5  (
            .in0(N__66468),
            .in1(N__66467),
            .in2(N__62610),
            .in3(N__62631),
            .lcout(\quad_counter1.n3006 ),
            .ltout(),
            .carryin(\quad_counter1.n30592 ),
            .carryout(\quad_counter1.n30593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_16_lut_LC_18_4_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_16_lut_LC_18_4_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_16_lut_LC_18_4_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_16_lut_LC_18_4_6  (
            .in0(N__66447),
            .in1(N__66446),
            .in2(N__62607),
            .in3(N__62628),
            .lcout(\quad_counter1.n3005 ),
            .ltout(),
            .carryin(\quad_counter1.n30593 ),
            .carryout(\quad_counter1.n30594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_17_lut_LC_18_4_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_17_lut_LC_18_4_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_17_lut_LC_18_4_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_17_lut_LC_18_4_7  (
            .in0(N__66426),
            .in1(N__66425),
            .in2(N__62611),
            .in3(N__62625),
            .lcout(\quad_counter1.n3004 ),
            .ltout(),
            .carryin(\quad_counter1.n30594 ),
            .carryout(\quad_counter1.n30595 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_18_lut_LC_18_5_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2018_18_lut_LC_18_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_18_lut_LC_18_5_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_18_lut_LC_18_5_0  (
            .in0(N__66804),
            .in1(N__66800),
            .in2(N__62618),
            .in3(N__62622),
            .lcout(\quad_counter1.n3003 ),
            .ltout(),
            .carryin(bfn_18_5_0_),
            .carryout(\quad_counter1.n30596 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2018_19_lut_LC_18_5_1 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_2018_19_lut_LC_18_5_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2018_19_lut_LC_18_5_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2018_19_lut_LC_18_5_1  (
            .in0(N__66772),
            .in1(N__66773),
            .in2(N__62619),
            .in3(N__62526),
            .lcout(\quad_counter1.n3002 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i6_2_lut_LC_18_5_2 .C_ON=1'b0;
    defparam \quad_counter1.i6_2_lut_LC_18_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i6_2_lut_LC_18_5_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter1.i6_2_lut_LC_18_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__66495),
            .in3(N__66799),
            .lcout(\quad_counter1.n18_adj_4459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1308_LC_18_5_3 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1308_LC_18_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1308_LC_18_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1308_LC_18_5_3  (
            .in0(N__66821),
            .in1(N__67244),
            .in2(N__67309),
            .in3(N__66848),
            .lcout(\quad_counter1.n22_adj_4474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i7_3_lut_LC_18_5_7 .C_ON=1'b0;
    defparam \quad_counter1.i7_3_lut_LC_18_5_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i7_3_lut_LC_18_5_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter1.i7_3_lut_LC_18_5_7  (
            .in0(_gnd_net_),
            .in1(N__67195),
            .in2(N__67282),
            .in3(N__67222),
            .lcout(\quad_counter1.n20_adj_4475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1309_LC_18_6_0 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1309_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1309_LC_18_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1309_LC_18_6_0  (
            .in0(N__62685),
            .in1(N__62676),
            .in2(N__66892),
            .in3(N__66943),
            .lcout(),
            .ltout(\quad_counter1.n24_adj_4476_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1310_LC_18_6_1 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1310_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1310_LC_18_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1310_LC_18_6_1  (
            .in0(N__66916),
            .in1(N__66997),
            .in2(N__62670),
            .in3(N__62667),
            .lcout(\quad_counter1.n3035 ),
            .ltout(\quad_counter1.n3035_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30729_1_lut_LC_18_6_2 .C_ON=1'b0;
    defparam \quad_counter1.i30729_1_lut_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30729_1_lut_LC_18_6_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30729_1_lut_LC_18_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62661),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1201_LC_18_8_1 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1201_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1201_LC_18_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1201_LC_18_8_1  (
            .in0(N__62658),
            .in1(N__62938),
            .in2(N__62904),
            .in3(N__62803),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_4_lut_adj_1202_LC_18_8_2 .C_ON=1'b0;
    defparam \quad_counter0.i2_4_lut_adj_1202_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_4_lut_adj_1202_LC_18_8_2 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i2_4_lut_adj_1202_LC_18_8_2  (
            .in0(N__62836),
            .in1(N__62866),
            .in2(N__62652),
            .in3(N__63199),
            .lcout(),
            .ltout(\quad_counter0.n7_adj_4383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1203_LC_18_8_3 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1203_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1203_LC_18_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1203_LC_18_8_3  (
            .in0(N__62725),
            .in1(N__63232),
            .in2(N__62649),
            .in3(N__63160),
            .lcout(\quad_counter0.n2243 ),
            .ltout(\quad_counter0.n2243_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30728_1_lut_LC_18_8_4 .C_ON=1'b0;
    defparam \quad_counter0.i30728_1_lut_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30728_1_lut_LC_18_8_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30728_1_lut_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62646),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_2_lut_LC_18_9_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_2_lut_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_2_lut_LC_18_9_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1549_2_lut_LC_18_9_0  (
            .in0(N__62998),
            .in1(N__62997),
            .in2(N__62767),
            .in3(N__62973),
            .lcout(\quad_counter0.n2319_adj_4385 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\quad_counter0.n30239 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_3_lut_LC_18_9_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_3_lut_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_3_lut_LC_18_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1549_3_lut_LC_18_9_1  (
            .in0(N__62970),
            .in1(N__62969),
            .in2(N__63116),
            .in3(N__62946),
            .lcout(\quad_counter0.n2318_adj_4386 ),
            .ltout(),
            .carryin(\quad_counter0.n30239 ),
            .carryout(\quad_counter0.n30240 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_4_lut_LC_18_9_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_4_lut_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_4_lut_LC_18_9_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1549_4_lut_LC_18_9_2  (
            .in0(N__62943),
            .in1(N__62939),
            .in2(N__62768),
            .in3(N__62907),
            .lcout(\quad_counter0.n2317_adj_4387 ),
            .ltout(),
            .carryin(\quad_counter0.n30240 ),
            .carryout(\quad_counter0.n30241 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_5_lut_LC_18_9_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_5_lut_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_5_lut_LC_18_9_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1549_5_lut_LC_18_9_3  (
            .in0(N__62902),
            .in1(N__62903),
            .in2(N__62771),
            .in3(N__62871),
            .lcout(\quad_counter0.n2316_adj_4391 ),
            .ltout(),
            .carryin(\quad_counter0.n30241 ),
            .carryout(\quad_counter0.n30242 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_6_lut_LC_18_9_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_6_lut_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_6_lut_LC_18_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1549_6_lut_LC_18_9_4  (
            .in0(N__62867),
            .in1(N__62868),
            .in2(N__62769),
            .in3(N__62841),
            .lcout(\quad_counter0.n2315_adj_4392 ),
            .ltout(),
            .carryin(\quad_counter0.n30242 ),
            .carryout(\quad_counter0.n30243 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_7_lut_LC_18_9_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_7_lut_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_7_lut_LC_18_9_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1549_7_lut_LC_18_9_5  (
            .in0(N__62838),
            .in1(N__62837),
            .in2(N__62772),
            .in3(N__62808),
            .lcout(\quad_counter0.n2314_adj_4388 ),
            .ltout(),
            .carryin(\quad_counter0.n30243 ),
            .carryout(\quad_counter0.n30244 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_8_lut_LC_18_9_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_8_lut_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_8_lut_LC_18_9_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1549_8_lut_LC_18_9_6  (
            .in0(N__62805),
            .in1(N__62804),
            .in2(N__62770),
            .in3(N__62730),
            .lcout(\quad_counter0.n2313 ),
            .ltout(),
            .carryin(\quad_counter0.n30244 ),
            .carryout(\quad_counter0.n30245 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_9_lut_LC_18_9_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_9_lut_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_9_lut_LC_18_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1549_9_lut_LC_18_9_7  (
            .in0(N__62727),
            .in1(N__62726),
            .in2(N__63117),
            .in3(N__62697),
            .lcout(\quad_counter0.n2312 ),
            .ltout(),
            .carryin(\quad_counter0.n30245 ),
            .carryout(\quad_counter0.n30246 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_10_lut_LC_18_10_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_10_lut_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_10_lut_LC_18_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1549_10_lut_LC_18_10_0  (
            .in0(N__63234),
            .in1(N__63233),
            .in2(N__63127),
            .in3(N__63204),
            .lcout(\quad_counter0.n2311 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\quad_counter0.n30247 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_11_lut_LC_18_10_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1549_11_lut_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_11_lut_LC_18_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1549_11_lut_LC_18_10_1  (
            .in0(N__63201),
            .in1(N__63200),
            .in2(N__63129),
            .in3(N__63168),
            .lcout(\quad_counter0.n2310 ),
            .ltout(),
            .carryin(\quad_counter0.n30247 ),
            .carryout(\quad_counter0.n30248 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1549_12_lut_LC_18_10_2 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1549_12_lut_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1549_12_lut_LC_18_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1549_12_lut_LC_18_10_2  (
            .in0(N__63165),
            .in1(N__63164),
            .in2(N__63128),
            .in3(N__63087),
            .lcout(\quad_counter0.n2309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i5_4_lut_adj_1207_LC_18_10_4 .C_ON=1'b0;
    defparam \quad_counter0.i5_4_lut_adj_1207_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i5_4_lut_adj_1207_LC_18_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i5_4_lut_adj_1207_LC_18_10_4  (
            .in0(N__63793),
            .in1(N__63063),
            .in2(N__63259),
            .in3(N__63084),
            .lcout(\quad_counter0.n2342_adj_4384 ),
            .ltout(\quad_counter0.n2342_adj_4384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30727_1_lut_LC_18_10_5 .C_ON=1'b0;
    defparam \quad_counter0.i30727_1_lut_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30727_1_lut_LC_18_10_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30727_1_lut_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__63075),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23645_2_lut_LC_18_10_6 .C_ON=1'b0;
    defparam \quad_counter0.i23645_2_lut_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23645_2_lut_LC_18_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23645_2_lut_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__63048),
            .in2(_gnd_net_),
            .in3(N__63016),
            .lcout(\quad_counter0.n28361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_2_lut_adj_1205_LC_18_10_7 .C_ON=1'b0;
    defparam \quad_counter0.i2_2_lut_adj_1205_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_2_lut_adj_1205_LC_18_10_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter0.i2_2_lut_adj_1205_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__63286),
            .in3(N__63769),
            .lcout(\quad_counter0.n8_adj_4390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_2_lut_LC_18_11_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_2_lut_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_2_lut_LC_18_11_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1616_2_lut_LC_18_11_0  (
            .in0(N__63052),
            .in1(N__63057),
            .in2(N__63361),
            .in3(N__63027),
            .lcout(\quad_counter0.n2419 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\quad_counter0.n30249 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_3_lut_LC_18_11_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_3_lut_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_3_lut_LC_18_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1616_3_lut_LC_18_11_1  (
            .in0(N__63024),
            .in1(N__63023),
            .in2(N__63739),
            .in3(N__63003),
            .lcout(\quad_counter0.n2418 ),
            .ltout(),
            .carryin(\quad_counter0.n30249 ),
            .carryout(\quad_counter0.n30250 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_4_lut_LC_18_11_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_4_lut_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_4_lut_LC_18_11_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1616_4_lut_LC_18_11_2  (
            .in0(N__63524),
            .in1(N__63523),
            .in2(N__63362),
            .in3(N__63495),
            .lcout(\quad_counter0.n2417 ),
            .ltout(),
            .carryin(\quad_counter0.n30250 ),
            .carryout(\quad_counter0.n30251 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_5_lut_LC_18_11_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_5_lut_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_5_lut_LC_18_11_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1616_5_lut_LC_18_11_3  (
            .in0(N__63488),
            .in1(N__63487),
            .in2(N__63365),
            .in3(N__63459),
            .lcout(\quad_counter0.n2416 ),
            .ltout(),
            .carryin(\quad_counter0.n30251 ),
            .carryout(\quad_counter0.n30252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_6_lut_LC_18_11_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_6_lut_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_6_lut_LC_18_11_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1616_6_lut_LC_18_11_4  (
            .in0(N__63455),
            .in1(N__63454),
            .in2(N__63363),
            .in3(N__63429),
            .lcout(\quad_counter0.n2415 ),
            .ltout(),
            .carryin(\quad_counter0.n30252 ),
            .carryout(\quad_counter0.n30253 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_7_lut_LC_18_11_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_7_lut_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_7_lut_LC_18_11_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1616_7_lut_LC_18_11_5  (
            .in0(N__63424),
            .in1(N__63425),
            .in2(N__63366),
            .in3(N__63396),
            .lcout(\quad_counter0.n2414 ),
            .ltout(),
            .carryin(\quad_counter0.n30253 ),
            .carryout(\quad_counter0.n30254 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_8_lut_LC_18_11_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_8_lut_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_8_lut_LC_18_11_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1616_8_lut_LC_18_11_6  (
            .in0(N__63392),
            .in1(N__63391),
            .in2(N__63364),
            .in3(N__63324),
            .lcout(\quad_counter0.n2413 ),
            .ltout(),
            .carryin(\quad_counter0.n30254 ),
            .carryout(\quad_counter0.n30255 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_9_lut_LC_18_11_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_9_lut_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_9_lut_LC_18_11_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1616_9_lut_LC_18_11_7  (
            .in0(N__63320),
            .in1(N__63319),
            .in2(N__63740),
            .in3(N__63291),
            .lcout(\quad_counter0.n2412 ),
            .ltout(),
            .carryin(\quad_counter0.n30255 ),
            .carryout(\quad_counter0.n30256 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_10_lut_LC_18_12_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_10_lut_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_10_lut_LC_18_12_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1616_10_lut_LC_18_12_0  (
            .in0(N__63288),
            .in1(N__63287),
            .in2(N__63753),
            .in3(N__63264),
            .lcout(\quad_counter0.n2411 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\quad_counter0.n30257 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_11_lut_LC_18_12_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_11_lut_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_11_lut_LC_18_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1616_11_lut_LC_18_12_1  (
            .in0(N__63261),
            .in1(N__63260),
            .in2(N__63755),
            .in3(N__63237),
            .lcout(\quad_counter0.n2410 ),
            .ltout(),
            .carryin(\quad_counter0.n30257 ),
            .carryout(\quad_counter0.n30258 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_12_lut_LC_18_12_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1616_12_lut_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_12_lut_LC_18_12_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1616_12_lut_LC_18_12_2  (
            .in0(N__63801),
            .in1(N__63800),
            .in2(N__63754),
            .in3(N__63780),
            .lcout(\quad_counter0.n2409 ),
            .ltout(),
            .carryin(\quad_counter0.n30258 ),
            .carryout(\quad_counter0.n30259 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1616_13_lut_LC_18_12_3 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1616_13_lut_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1616_13_lut_LC_18_12_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1616_13_lut_LC_18_12_3  (
            .in0(N__63776),
            .in1(N__63777),
            .in2(N__63756),
            .in3(N__63708),
            .lcout(\quad_counter0.n2408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_2_lut_LC_18_13_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_2_lut_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_2_lut_LC_18_13_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1683_2_lut_LC_18_13_0  (
            .in0(N__63705),
            .in1(N__63704),
            .in2(N__64222),
            .in3(N__63666),
            .lcout(\quad_counter0.n2519 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\quad_counter0.n30260 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_3_lut_LC_18_13_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_3_lut_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_3_lut_LC_18_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_3_lut_LC_18_13_1  (
            .in0(N__63658),
            .in1(N__63662),
            .in2(N__63969),
            .in3(N__63627),
            .lcout(\quad_counter0.n2518 ),
            .ltout(),
            .carryin(\quad_counter0.n30260 ),
            .carryout(\quad_counter0.n30261 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_4_lut_LC_18_13_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_4_lut_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_4_lut_LC_18_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1683_4_lut_LC_18_13_2  (
            .in0(N__63624),
            .in1(N__63623),
            .in2(N__64223),
            .in3(N__63597),
            .lcout(\quad_counter0.n2517 ),
            .ltout(),
            .carryin(\quad_counter0.n30261 ),
            .carryout(\quad_counter0.n30262 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_5_lut_LC_18_13_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_5_lut_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_5_lut_LC_18_13_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1683_5_lut_LC_18_13_3  (
            .in0(N__70628),
            .in1(N__70627),
            .in2(N__64226),
            .in3(N__63594),
            .lcout(\quad_counter0.n2516 ),
            .ltout(),
            .carryin(\quad_counter0.n30262 ),
            .carryout(\quad_counter0.n30263 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_6_lut_LC_18_13_4 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_6_lut_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_6_lut_LC_18_13_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1683_6_lut_LC_18_13_4  (
            .in0(N__63587),
            .in1(N__63586),
            .in2(N__64224),
            .in3(N__63561),
            .lcout(\quad_counter0.n2515 ),
            .ltout(),
            .carryin(\quad_counter0.n30263 ),
            .carryout(\quad_counter0.n30264 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_7_lut_LC_18_13_5 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_7_lut_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_7_lut_LC_18_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1683_7_lut_LC_18_13_5  (
            .in0(N__63551),
            .in1(N__63550),
            .in2(N__64227),
            .in3(N__63528),
            .lcout(\quad_counter0.n2514 ),
            .ltout(),
            .carryin(\quad_counter0.n30264 ),
            .carryout(\quad_counter0.n30265 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_8_lut_LC_18_13_6 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_8_lut_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_8_lut_LC_18_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter0.mod_61_add_1683_8_lut_LC_18_13_6  (
            .in0(N__70602),
            .in1(N__70601),
            .in2(N__64225),
            .in3(N__64182),
            .lcout(\quad_counter0.n2513 ),
            .ltout(),
            .carryin(\quad_counter0.n30265 ),
            .carryout(\quad_counter0.n30266 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_9_lut_LC_18_13_7 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_9_lut_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_9_lut_LC_18_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_9_lut_LC_18_13_7  (
            .in0(N__64179),
            .in1(N__64174),
            .in2(N__63970),
            .in3(N__64149),
            .lcout(\quad_counter0.n2512 ),
            .ltout(),
            .carryin(\quad_counter0.n30266 ),
            .carryout(\quad_counter0.n30267 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_10_lut_LC_18_14_0 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_10_lut_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_10_lut_LC_18_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_10_lut_LC_18_14_0  (
            .in0(N__64145),
            .in1(N__64144),
            .in2(N__63986),
            .in3(N__64116),
            .lcout(\quad_counter0.n2511 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\quad_counter0.n30268 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_11_lut_LC_18_14_1 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_11_lut_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_11_lut_LC_18_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_11_lut_LC_18_14_1  (
            .in0(N__64109),
            .in1(N__64108),
            .in2(N__63989),
            .in3(N__64083),
            .lcout(\quad_counter0.n2510 ),
            .ltout(),
            .carryin(\quad_counter0.n30268 ),
            .carryout(\quad_counter0.n30269 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_12_lut_LC_18_14_2 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_12_lut_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_12_lut_LC_18_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_12_lut_LC_18_14_2  (
            .in0(N__64078),
            .in1(N__64079),
            .in2(N__63987),
            .in3(N__64053),
            .lcout(\quad_counter0.n2509 ),
            .ltout(),
            .carryin(\quad_counter0.n30269 ),
            .carryout(\quad_counter0.n30270 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_13_lut_LC_18_14_3 .C_ON=1'b1;
    defparam \quad_counter0.mod_61_add_1683_13_lut_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_13_lut_LC_18_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_13_lut_LC_18_14_3  (
            .in0(N__64049),
            .in1(N__64048),
            .in2(N__63990),
            .in3(N__64023),
            .lcout(\quad_counter0.n2508 ),
            .ltout(),
            .carryin(\quad_counter0.n30270 ),
            .carryout(\quad_counter0.n30271 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.mod_61_add_1683_14_lut_LC_18_14_4 .C_ON=1'b0;
    defparam \quad_counter0.mod_61_add_1683_14_lut_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.mod_61_add_1683_14_lut_LC_18_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter0.mod_61_add_1683_14_lut_LC_18_14_4  (
            .in0(N__64018),
            .in1(N__64019),
            .in2(N__63988),
            .in3(N__63930),
            .lcout(\quad_counter0.n2507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i23629_2_lut_LC_18_14_6 .C_ON=1'b0;
    defparam \quad_counter0.i23629_2_lut_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i23629_2_lut_LC_18_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter0.i23629_2_lut_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__63927),
            .in2(_gnd_net_),
            .in3(N__63892),
            .lcout(\quad_counter0.n28345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i6_4_lut_adj_1214_LC_18_14_7 .C_ON=1'b0;
    defparam \quad_counter0.i6_4_lut_adj_1214_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i6_4_lut_adj_1214_LC_18_14_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i6_4_lut_adj_1214_LC_18_14_7  (
            .in0(N__63874),
            .in1(N__63856),
            .in2(N__63840),
            .in3(N__63817),
            .lcout(\quad_counter0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i7_4_lut_LC_18_15_4 .C_ON=1'b0;
    defparam \quad_counter0.i7_4_lut_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i7_4_lut_LC_18_15_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter0.i7_4_lut_LC_18_15_4  (
            .in0(N__64558),
            .in1(N__64537),
            .in2(N__64269),
            .in3(N__64521),
            .lcout(\quad_counter0.n2540 ),
            .ltout(\quad_counter0.n2540_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i30724_1_lut_LC_18_15_5 .C_ON=1'b0;
    defparam \quad_counter0.i30724_1_lut_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i30724_1_lut_LC_18_15_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter0.i30724_1_lut_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__64455),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.n36151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i4_4_lut_adj_1213_LC_18_15_6 .C_ON=1'b0;
    defparam \quad_counter0.i4_4_lut_adj_1213_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i4_4_lut_adj_1213_LC_18_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter0.i4_4_lut_adj_1213_LC_18_15_6  (
            .in0(N__64406),
            .in1(N__64383),
            .in2(N__64362),
            .in3(N__64353),
            .lcout(),
            .ltout(\quad_counter0.n10_adj_4397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i1_4_lut_adj_1215_LC_18_15_7 .C_ON=1'b0;
    defparam \quad_counter0.i1_4_lut_adj_1215_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i1_4_lut_adj_1215_LC_18_15_7 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \quad_counter0.i1_4_lut_adj_1215_LC_18_15_7  (
            .in0(N__64332),
            .in1(N__64311),
            .in2(N__64290),
            .in3(N__64285),
            .lcout(\quad_counter0.n9_adj_4398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_1_LC_18_16_0 .C_ON=1'b1;
    defparam \quad_counter1.add_623_1_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_1_LC_18_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \quad_counter1.add_623_1_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__64869),
            .in2(N__64903),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\quad_counter1.n30076 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_2_lut_LC_18_16_1 .C_ON=1'b1;
    defparam \quad_counter1.add_623_2_lut_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_2_lut_LC_18_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_2_lut_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__64260),
            .in2(N__101277),
            .in3(N__64236),
            .lcout(n2279),
            .ltout(),
            .carryin(\quad_counter1.n30076 ),
            .carryout(\quad_counter1.n30077 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_3_lut_LC_18_16_2 .C_ON=1'b1;
    defparam \quad_counter1.add_623_3_lut_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_3_lut_LC_18_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_3_lut_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__64870),
            .in2(N__84773),
            .in3(N__64233),
            .lcout(n2278),
            .ltout(),
            .carryin(\quad_counter1.n30077 ),
            .carryout(\quad_counter1.n30078 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_4_lut_LC_18_16_3 .C_ON=1'b1;
    defparam \quad_counter1.add_623_4_lut_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_4_lut_LC_18_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_4_lut_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__64876),
            .in2(N__86608),
            .in3(N__64230),
            .lcout(n2277),
            .ltout(),
            .carryin(\quad_counter1.n30078 ),
            .carryout(\quad_counter1.n30079 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_5_lut_LC_18_16_4 .C_ON=1'b1;
    defparam \quad_counter1.add_623_5_lut_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_5_lut_LC_18_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_5_lut_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__64871),
            .in2(N__83529),
            .in3(N__64602),
            .lcout(n2276),
            .ltout(),
            .carryin(\quad_counter1.n30079 ),
            .carryout(\quad_counter1.n30080 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_6_lut_LC_18_16_5 .C_ON=1'b1;
    defparam \quad_counter1.add_623_6_lut_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_6_lut_LC_18_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_6_lut_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__64877),
            .in2(N__85844),
            .in3(N__64599),
            .lcout(n2275),
            .ltout(),
            .carryin(\quad_counter1.n30080 ),
            .carryout(\quad_counter1.n30081 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_7_lut_LC_18_16_6 .C_ON=1'b1;
    defparam \quad_counter1.add_623_7_lut_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_7_lut_LC_18_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_7_lut_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__64872),
            .in2(N__85739),
            .in3(N__64596),
            .lcout(n2274),
            .ltout(),
            .carryin(\quad_counter1.n30081 ),
            .carryout(\quad_counter1.n30082 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_8_lut_LC_18_16_7 .C_ON=1'b1;
    defparam \quad_counter1.add_623_8_lut_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_8_lut_LC_18_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_8_lut_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__64878),
            .in2(N__94323),
            .in3(N__64593),
            .lcout(n2273),
            .ltout(),
            .carryin(\quad_counter1.n30082 ),
            .carryout(\quad_counter1.n30083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_9_lut_LC_18_17_0 .C_ON=1'b1;
    defparam \quad_counter1.add_623_9_lut_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_9_lut_LC_18_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_9_lut_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__64904),
            .in2(N__97961),
            .in3(N__64584),
            .lcout(n2272),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\quad_counter1.n30084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_10_lut_LC_18_17_1 .C_ON=1'b1;
    defparam \quad_counter1.add_623_10_lut_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_10_lut_LC_18_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_10_lut_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__75875),
            .in2(N__64957),
            .in3(N__64581),
            .lcout(n2271),
            .ltout(),
            .carryin(\quad_counter1.n30084 ),
            .carryout(\quad_counter1.n30085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_11_lut_LC_18_17_2 .C_ON=1'b1;
    defparam \quad_counter1.add_623_11_lut_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_11_lut_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_11_lut_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__64908),
            .in2(N__83060),
            .in3(N__64578),
            .lcout(n2270),
            .ltout(),
            .carryin(\quad_counter1.n30085 ),
            .carryout(\quad_counter1.n30086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_12_lut_LC_18_17_3 .C_ON=1'b1;
    defparam \quad_counter1.add_623_12_lut_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_12_lut_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_12_lut_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__83127),
            .in2(N__64958),
            .in3(N__64566),
            .lcout(n2269),
            .ltout(),
            .carryin(\quad_counter1.n30086 ),
            .carryout(\quad_counter1.n30087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_13_lut_LC_18_17_4 .C_ON=1'b1;
    defparam \quad_counter1.add_623_13_lut_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_13_lut_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_13_lut_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__64912),
            .in2(N__83484),
            .in3(N__64563),
            .lcout(n2268),
            .ltout(),
            .carryin(\quad_counter1.n30087 ),
            .carryout(\quad_counter1.n30088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_14_lut_LC_18_17_5 .C_ON=1'b1;
    defparam \quad_counter1.add_623_14_lut_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_14_lut_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_14_lut_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__76054),
            .in2(N__64959),
            .in3(N__64635),
            .lcout(n2267),
            .ltout(),
            .carryin(\quad_counter1.n30088 ),
            .carryout(\quad_counter1.n30089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_15_lut_LC_18_17_6 .C_ON=1'b1;
    defparam \quad_counter1.add_623_15_lut_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_15_lut_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_15_lut_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__64916),
            .in2(N__76096),
            .in3(N__64632),
            .lcout(n2266),
            .ltout(),
            .carryin(\quad_counter1.n30089 ),
            .carryout(\quad_counter1.n30090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_16_lut_LC_18_17_7 .C_ON=1'b1;
    defparam \quad_counter1.add_623_16_lut_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_16_lut_LC_18_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_16_lut_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__77281),
            .in2(N__64960),
            .in3(N__64629),
            .lcout(n2265),
            .ltout(),
            .carryin(\quad_counter1.n30090 ),
            .carryout(\quad_counter1.n30091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_17_lut_LC_18_18_0 .C_ON=1'b1;
    defparam \quad_counter1.add_623_17_lut_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_17_lut_LC_18_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_17_lut_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__64961),
            .in2(N__68183),
            .in3(N__64626),
            .lcout(n2264),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\quad_counter1.n30092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_18_lut_LC_18_18_1 .C_ON=1'b1;
    defparam \quad_counter1.add_623_18_lut_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_18_lut_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_18_lut_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__79179),
            .in2(N__64994),
            .in3(N__64623),
            .lcout(n2263),
            .ltout(),
            .carryin(\quad_counter1.n30092 ),
            .carryout(\quad_counter1.n30093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_19_lut_LC_18_18_2 .C_ON=1'b1;
    defparam \quad_counter1.add_623_19_lut_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_19_lut_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_19_lut_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__64965),
            .in2(N__77873),
            .in3(N__64620),
            .lcout(n2262),
            .ltout(),
            .carryin(\quad_counter1.n30093 ),
            .carryout(\quad_counter1.n30094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_20_lut_LC_18_18_3 .C_ON=1'b1;
    defparam \quad_counter1.add_623_20_lut_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_20_lut_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_20_lut_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__86353),
            .in2(N__64995),
            .in3(N__64617),
            .lcout(n2261),
            .ltout(),
            .carryin(\quad_counter1.n30094 ),
            .carryout(\quad_counter1.n30095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_21_lut_LC_18_18_4 .C_ON=1'b1;
    defparam \quad_counter1.add_623_21_lut_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_21_lut_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_21_lut_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__64969),
            .in2(N__83224),
            .in3(N__64608),
            .lcout(n2260),
            .ltout(),
            .carryin(\quad_counter1.n30095 ),
            .carryout(\quad_counter1.n30096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_22_lut_LC_18_18_5 .C_ON=1'b1;
    defparam \quad_counter1.add_623_22_lut_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_22_lut_LC_18_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_22_lut_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__76651),
            .in2(N__64996),
            .in3(N__64605),
            .lcout(n2259),
            .ltout(),
            .carryin(\quad_counter1.n30096 ),
            .carryout(\quad_counter1.n30097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_23_lut_LC_18_18_6 .C_ON=1'b1;
    defparam \quad_counter1.add_623_23_lut_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_23_lut_LC_18_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_23_lut_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__64973),
            .in2(N__85506),
            .in3(N__64677),
            .lcout(n2258),
            .ltout(),
            .carryin(\quad_counter1.n30097 ),
            .carryout(\quad_counter1.n30098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_24_lut_LC_18_18_7 .C_ON=1'b1;
    defparam \quad_counter1.add_623_24_lut_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_24_lut_LC_18_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_24_lut_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__71892),
            .in2(N__64997),
            .in3(N__64674),
            .lcout(n2257),
            .ltout(),
            .carryin(\quad_counter1.n30098 ),
            .carryout(\quad_counter1.n30099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_25_lut_LC_18_19_0 .C_ON=1'b1;
    defparam \quad_counter1.add_623_25_lut_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_25_lut_LC_18_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_25_lut_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__64977),
            .in2(N__67870),
            .in3(N__64665),
            .lcout(n2256),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\quad_counter1.n30100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_26_lut_LC_18_19_1 .C_ON=1'b1;
    defparam \quad_counter1.add_623_26_lut_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_26_lut_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_26_lut_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__68030),
            .in2(N__64998),
            .in3(N__64662),
            .lcout(n2255),
            .ltout(),
            .carryin(\quad_counter1.n30100 ),
            .carryout(\quad_counter1.n30101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_27_lut_LC_18_19_2 .C_ON=1'b1;
    defparam \quad_counter1.add_623_27_lut_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_27_lut_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_27_lut_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__64981),
            .in2(N__67798),
            .in3(N__64659),
            .lcout(n2254),
            .ltout(),
            .carryin(\quad_counter1.n30101 ),
            .carryout(\quad_counter1.n30102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_28_lut_LC_18_19_3 .C_ON=1'b1;
    defparam \quad_counter1.add_623_28_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_28_lut_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_28_lut_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__72278),
            .in2(N__64999),
            .in3(N__64644),
            .lcout(n2253),
            .ltout(),
            .carryin(\quad_counter1.n30102 ),
            .carryout(\quad_counter1.n30103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_29_lut_LC_18_19_4 .C_ON=1'b1;
    defparam \quad_counter1.add_623_29_lut_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_29_lut_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_29_lut_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__64985),
            .in2(N__77499),
            .in3(N__64641),
            .lcout(n2252),
            .ltout(),
            .carryin(\quad_counter1.n30103 ),
            .carryout(\quad_counter1.n30104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_30_lut_LC_18_19_5 .C_ON=1'b1;
    defparam \quad_counter1.add_623_30_lut_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_30_lut_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_30_lut_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__77343),
            .in2(N__65000),
            .in3(N__64638),
            .lcout(n2251),
            .ltout(),
            .carryin(\quad_counter1.n30104 ),
            .carryout(\quad_counter1.n30105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_31_lut_LC_18_19_6 .C_ON=1'b1;
    defparam \quad_counter1.add_623_31_lut_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_31_lut_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_31_lut_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__64989),
            .in2(N__77943),
            .in3(N__65007),
            .lcout(n2250),
            .ltout(),
            .carryin(\quad_counter1.n30105 ),
            .carryout(\quad_counter1.n30106 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_32_lut_LC_18_19_7 .C_ON=1'b1;
    defparam \quad_counter1.add_623_32_lut_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_32_lut_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_623_32_lut_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__86273),
            .in2(N__65001),
            .in3(N__65004),
            .lcout(n2249),
            .ltout(),
            .carryin(\quad_counter1.n30106 ),
            .carryout(\quad_counter1.n30107 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_623_33_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \quad_counter1.add_623_33_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_623_33_lut_LC_18_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter1.add_623_33_lut_LC_18_20_0  (
            .in0(N__85689),
            .in1(N__64993),
            .in2(_gnd_net_),
            .in3(N__64833),
            .lcout(n2248),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i6_LC_18_20_1 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i6_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i6_LC_18_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.control_mode_i0_i6_LC_18_20_1  (
            .in0(N__77618),
            .in1(N__72651),
            .in2(_gnd_net_),
            .in3(N__64830),
            .lcout(control_mode_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97632),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1745_LC_18_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1745_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1745_LC_18_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1745_LC_18_20_2  (
            .in0(N__72650),
            .in1(N__77558),
            .in2(N__79069),
            .in3(N__78038),
            .lcout(\c0.n33902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i27_LC_18_20_3 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i27_LC_18_20_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i27_LC_18_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i27_LC_18_20_3  (
            .in0(N__76540),
            .in1(N__64776),
            .in2(_gnd_net_),
            .in3(N__77489),
            .lcout(encoder1_position_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97632),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i22_LC_18_20_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i22_LC_18_20_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i22_LC_18_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i22_LC_18_20_4  (
            .in0(N__64770),
            .in1(N__76542),
            .in2(_gnd_net_),
            .in3(N__71889),
            .lcout(encoder1_position_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97632),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__7__5454_LC_18_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__7__5454_LC_18_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__7__5454_LC_18_20_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_8__7__5454_LC_18_20_5  (
            .in0(N__85100),
            .in1(N__84683),
            .in2(N__86499),
            .in3(N__64754),
            .lcout(data_out_frame_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97632),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i3_LC_18_20_6 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i3_LC_18_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i3_LC_18_20_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.control_mode_i0_i3_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__72148),
            .in2(N__64740),
            .in3(N__77619),
            .lcout(control_mode_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97632),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i28_LC_18_20_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i28_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i28_LC_18_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i28_LC_18_20_7  (
            .in0(N__76541),
            .in1(N__64683),
            .in2(_gnd_net_),
            .in3(N__77344),
            .lcout(encoder1_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97632),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_21_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_18_21_0  (
            .in0(N__90385),
            .in1(N__65025),
            .in2(N__90104),
            .in3(N__65187),
            .lcout(),
            .ltout(\c0.n36173_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36173_bdd_4_lut_4_lut_LC_18_21_1 .C_ON=1'b0;
    defparam \c0.n36173_bdd_4_lut_4_lut_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.n36173_bdd_4_lut_4_lut_LC_18_21_1 .LUT_INIT=16'b1111000011000010;
    LogicCell40 \c0.n36173_bdd_4_lut_4_lut_LC_18_21_1  (
            .in0(N__65175),
            .in1(N__90093),
            .in2(N__65154),
            .in3(N__96119),
            .lcout(n36176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30387_4_lut_LC_18_21_2 .C_ON=1'b0;
    defparam \c0.i30387_4_lut_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i30387_4_lut_LC_18_21_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.i30387_4_lut_LC_18_21_2  (
            .in0(N__90386),
            .in1(N__68133),
            .in2(N__90103),
            .in3(N__65193),
            .lcout(),
            .ltout(\c0.n35814_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30670_4_lut_LC_18_21_3 .C_ON=1'b0;
    defparam \c0.i30670_4_lut_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i30670_4_lut_LC_18_21_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.i30670_4_lut_LC_18_21_3  (
            .in0(N__68412),
            .in1(N__90094),
            .in2(N__65151),
            .in3(N__90387),
            .lcout(n36099),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1956_LC_18_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1956_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1956_LC_18_21_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i1_2_lut_adj_1956_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(N__68272),
            .in2(_gnd_net_),
            .in3(N__78689),
            .lcout(\c0.n33249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i30699_3_lut_LC_18_21_6 .C_ON=1'b0;
    defparam \c0.rx.i30699_3_lut_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i30699_3_lut_LC_18_21_6 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.rx.i30699_3_lut_LC_18_21_6  (
            .in0(N__65147),
            .in1(N__65088),
            .in2(_gnd_net_),
            .in3(N__76992),
            .lcout(\c0.rx.n34953 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_18_21_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_18_21_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_18_21_7  (
            .in0(N__68387),
            .in1(N__65036),
            .in2(_gnd_net_),
            .in3(N__96118),
            .lcout(\c0.n5_adj_4707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i0_LC_18_22_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i0_LC_18_22_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i0_LC_18_22_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i0_LC_18_22_0  (
            .in0(N__86118),
            .in1(N__65019),
            .in2(_gnd_net_),
            .in3(N__85593),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97662),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i3_LC_18_22_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i3_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i3_LC_18_22_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i3_LC_18_22_1  (
            .in0(N__85441),
            .in1(N__65013),
            .in2(_gnd_net_),
            .in3(N__86119),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97662),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i6_LC_18_22_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i6_LC_18_22_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i6_LC_18_22_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i6_LC_18_22_2  (
            .in0(N__86120),
            .in1(N__65283),
            .in2(_gnd_net_),
            .in3(N__75825),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_18_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_18_22_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i44_LC_18_22_3  (
            .in0(N__68303),
            .in1(N__78556),
            .in2(N__65262),
            .in3(N__78995),
            .lcout(\c0.data_in_frame_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97662),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i17_LC_18_22_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i17_LC_18_22_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i17_LC_18_22_4 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \quad_counter1.count_i0_i17_LC_18_22_4  (
            .in0(N__77856),
            .in1(N__65235),
            .in2(N__76583),
            .in3(_gnd_net_),
            .lcout(encoder1_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97662),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i24_LC_18_22_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i24_LC_18_22_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i24_LC_18_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i24_LC_18_22_5  (
            .in0(N__68028),
            .in1(N__65226),
            .in2(_gnd_net_),
            .in3(N__76565),
            .lcout(encoder1_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30386_3_lut_LC_18_22_6 .C_ON=1'b0;
    defparam \c0.i30386_3_lut_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30386_3_lut_LC_18_22_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i30386_3_lut_LC_18_22_6  (
            .in0(N__96120),
            .in1(N__65216),
            .in2(_gnd_net_),
            .in3(N__65204),
            .lcout(\c0.n35813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30618_2_lut_LC_18_22_7 .C_ON=1'b0;
    defparam \c0.i30618_2_lut_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30618_2_lut_LC_18_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i30618_2_lut_LC_18_22_7  (
            .in0(N__68048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__96121),
            .lcout(\c0.n35964 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i207_LC_18_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i207_LC_18_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i207_LC_18_23_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i207_LC_18_23_0  (
            .in0(N__79816),
            .in1(N__87240),
            .in2(N__65846),
            .in3(N__73655),
            .lcout(\c0.data_in_frame_25_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1344_LC_18_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1344_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1344_LC_18_23_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1344_LC_18_23_1  (
            .in0(N__91468),
            .in1(N__91555),
            .in2(N__91365),
            .in3(N__91648),
            .lcout(\c0.n12_adj_4519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i20_LC_18_23_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i20_LC_18_23_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i20_LC_18_23_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i20_LC_18_23_2  (
            .in0(N__71983),
            .in1(N__65181),
            .in2(_gnd_net_),
            .in3(N__86117),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_2053_LC_18_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_2053_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_2053_LC_18_23_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_2053_LC_18_23_3  (
            .in0(N__91469),
            .in1(N__91556),
            .in2(N__91366),
            .in3(N__91649),
            .lcout(\c0.n12_adj_4526 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1661_LC_18_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1661_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1661_LC_18_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1661_LC_18_23_4  (
            .in0(N__69244),
            .in1(N__65317),
            .in2(_gnd_net_),
            .in3(N__65836),
            .lcout(\c0.n33407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i14_LC_18_23_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i14_LC_18_23_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i14_LC_18_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i14_LC_18_23_5  (
            .in0(N__86116),
            .in1(N__65379),
            .in2(_gnd_net_),
            .in3(N__85781),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1600_LC_18_23_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1600_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1600_LC_18_23_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.i1_4_lut_adj_1600_LC_18_23_6  (
            .in0(N__65373),
            .in1(N__91467),
            .in2(N__90497),
            .in3(N__91352),
            .lcout(\c0.n18084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i208_LC_18_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i208_LC_18_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i208_LC_18_23_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i208_LC_18_23_7  (
            .in0(N__87239),
            .in1(N__80016),
            .in2(N__65324),
            .in3(N__79817),
            .lcout(\c0.data_in_frame_25_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97676),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1938_LC_18_24_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1938_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1938_LC_18_24_0 .LUT_INIT=16'b1111111011101111;
    LogicCell40 \c0.i10_4_lut_adj_1938_LC_18_24_0  (
            .in0(N__69324),
            .in1(N__69261),
            .in2(N__73257),
            .in3(N__66104),
            .lcout(),
            .ltout(\c0.n28_adj_4762_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1941_LC_18_24_1 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1941_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1941_LC_18_24_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i17_4_lut_adj_1941_LC_18_24_1  (
            .in0(N__65304),
            .in1(N__65973),
            .in2(N__65295),
            .in3(N__65685),
            .lcout(n35693),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i30_LC_18_24_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i30_LC_18_24_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i30_LC_18_24_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i30_LC_18_24_2  (
            .in0(N__76564),
            .in1(N__65292),
            .in2(_gnd_net_),
            .in3(N__86258),
            .lcout(encoder1_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i177_LC_18_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i177_LC_18_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i177_LC_18_24_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i177_LC_18_24_3  (
            .in0(N__89760),
            .in1(N__80974),
            .in2(N__66025),
            .in3(N__72925),
            .lcout(\c0.data_in_frame_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1939_LC_18_24_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1939_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1939_LC_18_24_4 .LUT_INIT=16'b1111111110110111;
    LogicCell40 \c0.i13_4_lut_adj_1939_LC_18_24_4  (
            .in0(N__65418),
            .in1(N__65706),
            .in2(N__65820),
            .in3(N__65697),
            .lcout(\c0.n31_adj_4763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i184_LC_18_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i184_LC_18_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i184_LC_18_24_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i184_LC_18_24_5  (
            .in0(N__89761),
            .in1(N__72924),
            .in2(N__65673),
            .in3(N__80017),
            .lcout(\c0.data_in_frame_22_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97693),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1739_LC_18_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1739_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1739_LC_18_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1739_LC_18_25_0  (
            .in0(N__79477),
            .in1(N__78357),
            .in2(N__65526),
            .in3(N__65474),
            .lcout(\c0.n31374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1772_LC_18_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1772_LC_18_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1772_LC_18_25_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1772_LC_18_25_1  (
            .in0(N__65525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65473),
            .lcout(\c0.n18961 ),
            .ltout(\c0.n18961_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1641_LC_18_25_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1641_LC_18_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1641_LC_18_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1641_LC_18_25_2  (
            .in0(N__68710),
            .in1(N__65616),
            .in2(N__65604),
            .in3(N__65532),
            .lcout(\c0.n14_adj_4668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1527_LC_18_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1527_LC_18_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1527_LC_18_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1527_LC_18_25_3  (
            .in0(N__65523),
            .in1(N__65471),
            .in2(_gnd_net_),
            .in3(N__65588),
            .lcout(\c0.n32263 ),
            .ltout(\c0.n32263_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1523_LC_18_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1523_LC_18_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1523_LC_18_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1523_LC_18_25_4  (
            .in0(_gnd_net_),
            .in1(N__78724),
            .in2(N__65535),
            .in3(N__78356),
            .lcout(\c0.n33576 ),
            .ltout(\c0.n33576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1738_LC_18_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1738_LC_18_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1738_LC_18_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1738_LC_18_25_5  (
            .in0(N__65524),
            .in1(N__65472),
            .in2(N__65445),
            .in3(N__79476),
            .lcout(\c0.n33577 ),
            .ltout(\c0.n33577_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1927_LC_18_25_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1927_LC_18_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1927_LC_18_25_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1927_LC_18_25_6  (
            .in0(N__73689),
            .in1(N__68687),
            .in2(N__65442),
            .in3(N__65439),
            .lcout(\c0.n14_adj_4757 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_1701_LC_18_25_7 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_1701_LC_18_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_1701_LC_18_25_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_1701_LC_18_25_7  (
            .in0(N__65946),
            .in1(N__68856),
            .in2(N__73169),
            .in3(N__74715),
            .lcout(\c0.n30_adj_4706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1929_LC_18_26_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1929_LC_18_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1929_LC_18_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1929_LC_18_26_0  (
            .in0(N__65898),
            .in1(N__65875),
            .in2(N__65847),
            .in3(N__74218),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1667_LC_18_26_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1667_LC_18_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1667_LC_18_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1667_LC_18_26_2  (
            .in0(N__68793),
            .in1(N__72708),
            .in2(_gnd_net_),
            .in3(N__73399),
            .lcout(\c0.n33819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1766_LC_18_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1766_LC_18_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1766_LC_18_26_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1766_LC_18_26_3  (
            .in0(_gnd_net_),
            .in1(N__65731),
            .in2(_gnd_net_),
            .in3(N__65744),
            .lcout(),
            .ltout(\c0.n32294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_1695_LC_18_26_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_1695_LC_18_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_1695_LC_18_26_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i13_4_lut_adj_1695_LC_18_26_4  (
            .in0(N__66017),
            .in1(N__65808),
            .in2(N__65796),
            .in3(N__68953),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_1528_LC_18_26_5 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1528_LC_18_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1528_LC_18_26_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1528_LC_18_26_5  (
            .in0(N__65781),
            .in1(N__79475),
            .in2(N__65775),
            .in3(N__66367),
            .lcout(\c0.n8_adj_4622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1522_LC_18_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1522_LC_18_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1522_LC_18_26_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1522_LC_18_26_6  (
            .in0(N__65745),
            .in1(_gnd_net_),
            .in2(N__65736),
            .in3(N__65960),
            .lcout(\c0.n34006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1688_LC_18_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1688_LC_18_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1688_LC_18_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1688_LC_18_27_1  (
            .in0(_gnd_net_),
            .in1(N__69111),
            .in2(_gnd_net_),
            .in3(N__68631),
            .lcout(\c0.n33816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1631_LC_18_27_2 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1631_LC_18_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1631_LC_18_27_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_adj_1631_LC_18_27_2  (
            .in0(N__66201),
            .in1(N__74018),
            .in2(N__74806),
            .in3(N__66195),
            .lcout(\c0.n32316 ),
            .ltout(\c0.n32316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1623_LC_18_27_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1623_LC_18_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1623_LC_18_27_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1623_LC_18_27_3  (
            .in0(N__74492),
            .in1(N__68630),
            .in2(N__66177),
            .in3(N__66174),
            .lcout(),
            .ltout(\c0.n19_adj_4658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1625_LC_18_27_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1625_LC_18_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1625_LC_18_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1625_LC_18_27_4  (
            .in0(N__66162),
            .in1(N__69275),
            .in2(N__66156),
            .in3(N__66153),
            .lcout(),
            .ltout(\c0.n5_adj_4660_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1626_LC_18_27_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1626_LC_18_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1626_LC_18_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1626_LC_18_27_5  (
            .in0(N__69349),
            .in1(N__74156),
            .in2(N__66141),
            .in3(N__66133),
            .lcout(\c0.n33792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1917_LC_18_27_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1917_LC_18_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1917_LC_18_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1917_LC_18_27_7  (
            .in0(N__68984),
            .in1(N__66083),
            .in2(N__74022),
            .in3(N__66056),
            .lcout(\c0.n17_adj_4753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i230_LC_18_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i230_LC_18_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i230_LC_18_28_0 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i230_LC_18_28_0  (
            .in0(N__75062),
            .in1(N__66042),
            .in2(N__73950),
            .in3(N__79867),
            .lcout(\c0.data_in_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30362_4_lut_LC_18_28_3 .C_ON=1'b0;
    defparam \c0.i30362_4_lut_LC_18_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i30362_4_lut_LC_18_28_3 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.i30362_4_lut_LC_18_28_3  (
            .in0(N__66041),
            .in1(N__66033),
            .in2(N__66027),
            .in3(N__65979),
            .lcout(\c0.n35787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i210_LC_18_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i210_LC_18_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i210_LC_18_28_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i210_LC_18_28_4  (
            .in0(N__75361),
            .in1(N__80320),
            .in2(N__65964),
            .in3(N__79866),
            .lcout(\c0.data_in_frame_26_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i232_LC_18_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i232_LC_18_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i232_LC_18_28_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i232_LC_18_28_5  (
            .in0(N__79865),
            .in1(N__80057),
            .in2(N__69180),
            .in3(N__73946),
            .lcout(\c0.data_in_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97762),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1657_LC_18_28_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1657_LC_18_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1657_LC_18_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1657_LC_18_28_6  (
            .in0(N__74094),
            .in1(N__73371),
            .in2(N__74499),
            .in3(N__66408),
            .lcout(),
            .ltout(\c0.n10_adj_4673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1658_LC_18_28_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1658_LC_18_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1658_LC_18_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1658_LC_18_28_7  (
            .in0(_gnd_net_),
            .in1(N__66390),
            .in2(N__66375),
            .in3(N__66372),
            .lcout(\c0.n31784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_2_lut_LC_19_2_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_2_lut_LC_19_2_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_2_lut_LC_19_2_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1951_2_lut_LC_19_2_0  (
            .in0(N__81843),
            .in1(N__81842),
            .in2(N__69565),
            .in3(N__66321),
            .lcout(\quad_counter1.n2919 ),
            .ltout(),
            .carryin(bfn_19_2_0_),
            .carryout(\quad_counter1.n30564 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_3_lut_LC_19_2_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_3_lut_LC_19_2_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_3_lut_LC_19_2_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_3_lut_LC_19_2_1  (
            .in0(N__69426),
            .in1(N__69425),
            .in2(N__69524),
            .in3(N__66291),
            .lcout(\quad_counter1.n2918 ),
            .ltout(),
            .carryin(\quad_counter1.n30564 ),
            .carryout(\quad_counter1.n30565 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_4_lut_LC_19_2_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_4_lut_LC_19_2_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_4_lut_LC_19_2_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1951_4_lut_LC_19_2_2  (
            .in0(N__69399),
            .in1(N__69398),
            .in2(N__69566),
            .in3(N__66267),
            .lcout(\quad_counter1.n2917 ),
            .ltout(),
            .carryin(\quad_counter1.n30565 ),
            .carryout(\quad_counter1.n30566 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_5_lut_LC_19_2_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_5_lut_LC_19_2_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_5_lut_LC_19_2_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1951_5_lut_LC_19_2_3  (
            .in0(N__69375),
            .in1(N__69374),
            .in2(N__69569),
            .in3(N__66246),
            .lcout(\quad_counter1.n2916 ),
            .ltout(),
            .carryin(\quad_counter1.n30566 ),
            .carryout(\quad_counter1.n30567 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_6_lut_LC_19_2_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_6_lut_LC_19_2_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_6_lut_LC_19_2_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1951_6_lut_LC_19_2_4  (
            .in0(N__69732),
            .in1(N__69731),
            .in2(N__69567),
            .in3(N__66225),
            .lcout(\quad_counter1.n2915 ),
            .ltout(),
            .carryin(\quad_counter1.n30567 ),
            .carryout(\quad_counter1.n30568 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_7_lut_LC_19_2_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_7_lut_LC_19_2_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_7_lut_LC_19_2_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1951_7_lut_LC_19_2_5  (
            .in0(N__69705),
            .in1(N__69704),
            .in2(N__69570),
            .in3(N__66204),
            .lcout(\quad_counter1.n2914 ),
            .ltout(),
            .carryin(\quad_counter1.n30568 ),
            .carryout(\quad_counter1.n30569 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_8_lut_LC_19_2_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_8_lut_LC_19_2_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_8_lut_LC_19_2_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1951_8_lut_LC_19_2_6  (
            .in0(N__69681),
            .in1(N__69677),
            .in2(N__69568),
            .in3(N__66603),
            .lcout(\quad_counter1.n2913 ),
            .ltout(),
            .carryin(\quad_counter1.n30569 ),
            .carryout(\quad_counter1.n30570 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_9_lut_LC_19_2_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_9_lut_LC_19_2_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_9_lut_LC_19_2_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_9_lut_LC_19_2_7  (
            .in0(N__74601),
            .in1(N__74597),
            .in2(N__69525),
            .in3(N__66573),
            .lcout(\quad_counter1.n2912 ),
            .ltout(),
            .carryin(\quad_counter1.n30570 ),
            .carryout(\quad_counter1.n30571 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_10_lut_LC_19_3_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_10_lut_LC_19_3_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_10_lut_LC_19_3_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_10_lut_LC_19_3_0  (
            .in0(N__69648),
            .in1(N__69647),
            .in2(N__69515),
            .in3(N__66552),
            .lcout(\quad_counter1.n2911 ),
            .ltout(),
            .carryin(bfn_19_3_0_),
            .carryout(\quad_counter1.n30572 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_11_lut_LC_19_3_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_11_lut_LC_19_3_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_11_lut_LC_19_3_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_11_lut_LC_19_3_1  (
            .in0(N__74667),
            .in1(N__74666),
            .in2(N__69519),
            .in3(N__66528),
            .lcout(\quad_counter1.n2910 ),
            .ltout(),
            .carryin(\quad_counter1.n30572 ),
            .carryout(\quad_counter1.n30573 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_12_lut_LC_19_3_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_12_lut_LC_19_3_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_12_lut_LC_19_3_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_12_lut_LC_19_3_2  (
            .in0(N__74625),
            .in1(N__74624),
            .in2(N__69516),
            .in3(N__66498),
            .lcout(\quad_counter1.n2909 ),
            .ltout(),
            .carryin(\quad_counter1.n30573 ),
            .carryout(\quad_counter1.n30574 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_13_lut_LC_19_3_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_13_lut_LC_19_3_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_13_lut_LC_19_3_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_13_lut_LC_19_3_3  (
            .in0(N__69620),
            .in1(N__69621),
            .in2(N__69520),
            .in3(N__66471),
            .lcout(\quad_counter1.n2908 ),
            .ltout(),
            .carryin(\quad_counter1.n30574 ),
            .carryout(\quad_counter1.n30575 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_14_lut_LC_19_3_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_14_lut_LC_19_3_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_14_lut_LC_19_3_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_14_lut_LC_19_3_4  (
            .in0(N__69594),
            .in1(N__69593),
            .in2(N__69517),
            .in3(N__66450),
            .lcout(\quad_counter1.n2907 ),
            .ltout(),
            .carryin(\quad_counter1.n30575 ),
            .carryout(\quad_counter1.n30576 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_15_lut_LC_19_3_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_15_lut_LC_19_3_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_15_lut_LC_19_3_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_15_lut_LC_19_3_5  (
            .in0(N__74646),
            .in1(N__74645),
            .in2(N__69521),
            .in3(N__66429),
            .lcout(\quad_counter1.n2906 ),
            .ltout(),
            .carryin(\quad_counter1.n30576 ),
            .carryout(\quad_counter1.n30577 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_16_lut_LC_19_3_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_16_lut_LC_19_3_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_16_lut_LC_19_3_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_16_lut_LC_19_3_6  (
            .in0(N__69840),
            .in1(N__69836),
            .in2(N__69518),
            .in3(N__66807),
            .lcout(\quad_counter1.n2905 ),
            .ltout(),
            .carryin(\quad_counter1.n30577 ),
            .carryout(\quad_counter1.n30578 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_17_lut_LC_19_3_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1951_17_lut_LC_19_3_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_17_lut_LC_19_3_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_17_lut_LC_19_3_7  (
            .in0(N__69810),
            .in1(N__69805),
            .in2(N__69522),
            .in3(N__66780),
            .lcout(\quad_counter1.n2904 ),
            .ltout(),
            .carryin(\quad_counter1.n30578 ),
            .carryout(\quad_counter1.n30579 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1951_18_lut_LC_19_4_0 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1951_18_lut_LC_19_4_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1951_18_lut_LC_19_4_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1951_18_lut_LC_19_4_0  (
            .in0(N__69772),
            .in1(N__69773),
            .in2(N__69523),
            .in3(N__66777),
            .lcout(\quad_counter1.n2903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_2_lut_LC_19_5_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_2_lut_LC_19_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_2_lut_LC_19_5_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2085_2_lut_LC_19_5_0  (
            .in0(N__81930),
            .in1(N__81929),
            .in2(N__67045),
            .in3(N__66753),
            .lcout(\quad_counter1.n3119 ),
            .ltout(),
            .carryin(bfn_19_5_0_),
            .carryout(\quad_counter1.n30597 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_3_lut_LC_19_5_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_3_lut_LC_19_5_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_3_lut_LC_19_5_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_3_lut_LC_19_5_1  (
            .in0(N__66750),
            .in1(N__66749),
            .in2(N__67178),
            .in3(N__66726),
            .lcout(\quad_counter1.n3118 ),
            .ltout(),
            .carryin(\quad_counter1.n30597 ),
            .carryout(\quad_counter1.n30598 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_4_lut_LC_19_5_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_4_lut_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_4_lut_LC_19_5_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2085_4_lut_LC_19_5_2  (
            .in0(N__66723),
            .in1(N__66722),
            .in2(N__67046),
            .in3(N__66699),
            .lcout(\quad_counter1.n3117 ),
            .ltout(),
            .carryin(\quad_counter1.n30598 ),
            .carryout(\quad_counter1.n30599 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_5_lut_LC_19_5_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_5_lut_LC_19_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_5_lut_LC_19_5_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2085_5_lut_LC_19_5_3  (
            .in0(N__66696),
            .in1(N__66695),
            .in2(N__67049),
            .in3(N__66675),
            .lcout(\quad_counter1.n3116 ),
            .ltout(),
            .carryin(\quad_counter1.n30599 ),
            .carryout(\quad_counter1.n30600 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_6_lut_LC_19_5_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_6_lut_LC_19_5_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_6_lut_LC_19_5_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2085_6_lut_LC_19_5_4  (
            .in0(N__66672),
            .in1(N__66671),
            .in2(N__67047),
            .in3(N__66651),
            .lcout(\quad_counter1.n3115 ),
            .ltout(),
            .carryin(\quad_counter1.n30600 ),
            .carryout(\quad_counter1.n30601 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_7_lut_LC_19_5_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_7_lut_LC_19_5_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_7_lut_LC_19_5_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2085_7_lut_LC_19_5_5  (
            .in0(N__66648),
            .in1(N__66647),
            .in2(N__67050),
            .in3(N__66627),
            .lcout(\quad_counter1.n3114 ),
            .ltout(),
            .carryin(\quad_counter1.n30601 ),
            .carryout(\quad_counter1.n30602 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_8_lut_LC_19_5_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_8_lut_LC_19_5_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_8_lut_LC_19_5_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2085_8_lut_LC_19_5_6  (
            .in0(N__67071),
            .in1(N__67070),
            .in2(N__67048),
            .in3(N__67008),
            .lcout(\quad_counter1.n3113 ),
            .ltout(),
            .carryin(\quad_counter1.n30602 ),
            .carryout(\quad_counter1.n30603 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_9_lut_LC_19_5_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_9_lut_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_9_lut_LC_19_5_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_9_lut_LC_19_5_7  (
            .in0(N__67005),
            .in1(N__67004),
            .in2(N__67179),
            .in3(N__66978),
            .lcout(\quad_counter1.n3112 ),
            .ltout(),
            .carryin(\quad_counter1.n30603 ),
            .carryout(\quad_counter1.n30604 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_10_lut_LC_19_6_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_10_lut_LC_19_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_10_lut_LC_19_6_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_10_lut_LC_19_6_0  (
            .in0(N__66975),
            .in1(N__66974),
            .in2(N__67167),
            .in3(N__66954),
            .lcout(\quad_counter1.n3111 ),
            .ltout(),
            .carryin(bfn_19_6_0_),
            .carryout(\quad_counter1.n30605 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_11_lut_LC_19_6_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_11_lut_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_11_lut_LC_19_6_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_11_lut_LC_19_6_1  (
            .in0(N__66951),
            .in1(N__66950),
            .in2(N__67171),
            .in3(N__66927),
            .lcout(\quad_counter1.n3110 ),
            .ltout(),
            .carryin(\quad_counter1.n30605 ),
            .carryout(\quad_counter1.n30606 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_12_lut_LC_19_6_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_12_lut_LC_19_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_12_lut_LC_19_6_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_12_lut_LC_19_6_2  (
            .in0(N__66924),
            .in1(N__66923),
            .in2(N__67168),
            .in3(N__66897),
            .lcout(\quad_counter1.n3109 ),
            .ltout(),
            .carryin(\quad_counter1.n30606 ),
            .carryout(\quad_counter1.n30607 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_13_lut_LC_19_6_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_13_lut_LC_19_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_13_lut_LC_19_6_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_13_lut_LC_19_6_3  (
            .in0(N__66894),
            .in1(N__66893),
            .in2(N__67172),
            .in3(N__66864),
            .lcout(\quad_counter1.n3108 ),
            .ltout(),
            .carryin(\quad_counter1.n30607 ),
            .carryout(\quad_counter1.n30608 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_14_lut_LC_19_6_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_14_lut_LC_19_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_14_lut_LC_19_6_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_14_lut_LC_19_6_4  (
            .in0(N__66861),
            .in1(N__66860),
            .in2(N__67169),
            .in3(N__66837),
            .lcout(\quad_counter1.n3107 ),
            .ltout(),
            .carryin(\quad_counter1.n30608 ),
            .carryout(\quad_counter1.n30609 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_15_lut_LC_19_6_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_15_lut_LC_19_6_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_15_lut_LC_19_6_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_15_lut_LC_19_6_5  (
            .in0(N__66834),
            .in1(N__66833),
            .in2(N__67173),
            .in3(N__66810),
            .lcout(\quad_counter1.n3106 ),
            .ltout(),
            .carryin(\quad_counter1.n30609 ),
            .carryout(\quad_counter1.n30610 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_16_lut_LC_19_6_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_16_lut_LC_19_6_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_16_lut_LC_19_6_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_16_lut_LC_19_6_6  (
            .in0(N__67311),
            .in1(N__67310),
            .in2(N__67170),
            .in3(N__67287),
            .lcout(\quad_counter1.n3105 ),
            .ltout(),
            .carryin(\quad_counter1.n30610 ),
            .carryout(\quad_counter1.n30611 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_17_lut_LC_19_6_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_17_lut_LC_19_6_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_17_lut_LC_19_6_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_17_lut_LC_19_6_7  (
            .in0(N__67284),
            .in1(N__67283),
            .in2(N__67174),
            .in3(N__67260),
            .lcout(\quad_counter1.n3104 ),
            .ltout(),
            .carryin(\quad_counter1.n30611 ),
            .carryout(\quad_counter1.n30612 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_18_lut_LC_19_7_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_18_lut_LC_19_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_18_lut_LC_19_7_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_18_lut_LC_19_7_0  (
            .in0(N__67256),
            .in1(N__67257),
            .in2(N__67175),
            .in3(N__67233),
            .lcout(\quad_counter1.n3103 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\quad_counter1.n30613 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_19_lut_LC_19_7_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2085_19_lut_LC_19_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_19_lut_LC_19_7_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_19_lut_LC_19_7_1  (
            .in0(N__67230),
            .in1(N__67229),
            .in2(N__67177),
            .in3(N__67209),
            .lcout(\quad_counter1.n3102 ),
            .ltout(),
            .carryin(\quad_counter1.n30613 ),
            .carryout(\quad_counter1.n30614 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2085_20_lut_LC_19_7_2 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_2085_20_lut_LC_19_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2085_20_lut_LC_19_7_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2085_20_lut_LC_19_7_2  (
            .in0(N__67206),
            .in1(N__67205),
            .in2(N__67176),
            .in3(N__67083),
            .lcout(\quad_counter1.n3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_adj_1311_LC_19_7_3 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_adj_1311_LC_19_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_adj_1311_LC_19_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \quad_counter1.i2_2_lut_adj_1311_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__69991),
            .in2(_gnd_net_),
            .in3(N__70114),
            .lcout(\quad_counter1.n8_adj_4477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_2_lut_LC_19_7_4 .C_ON=1'b0;
    defparam \quad_counter1.i4_2_lut_LC_19_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_2_lut_LC_19_7_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter1.i4_2_lut_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__70393),
            .in3(N__70903),
            .lcout(),
            .ltout(\quad_counter1.n18_adj_4479_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1316_LC_19_7_5 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1316_LC_19_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1316_LC_19_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1316_LC_19_7_5  (
            .in0(N__71003),
            .in1(N__70496),
            .in2(N__67080),
            .in3(N__67077),
            .lcout(\quad_counter1.n26_adj_4482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1314_LC_19_7_6 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1314_LC_19_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1314_LC_19_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1314_LC_19_7_6  (
            .in0(N__70339),
            .in1(N__70948),
            .in2(N__70246),
            .in3(N__70291),
            .lcout(\quad_counter1.n24_adj_4480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1320_LC_19_8_5 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1320_LC_19_8_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1320_LC_19_8_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1320_LC_19_8_5  (
            .in0(N__70039),
            .in1(N__81429),
            .in2(N__70273),
            .in3(N__70087),
            .lcout(\quad_counter1.n19_adj_4485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_2_lut_adj_1321_LC_19_9_0 .C_ON=1'b0;
    defparam \quad_counter1.i1_2_lut_adj_1321_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_2_lut_adj_1321_LC_19_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i1_2_lut_adj_1321_LC_19_9_0  (
            .in0(_gnd_net_),
            .in1(N__70871),
            .in2(_gnd_net_),
            .in3(N__69862),
            .lcout(\quad_counter1.n16_adj_4486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1322_LC_19_9_1 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1322_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1322_LC_19_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1322_LC_19_9_1  (
            .in0(N__70715),
            .in1(N__70417),
            .in2(N__70477),
            .in3(N__69919),
            .lcout(\quad_counter1.n24_adj_4487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1319_LC_19_9_3 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1319_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1319_LC_19_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1319_LC_19_9_3  (
            .in0(N__70315),
            .in1(N__70979),
            .in2(N__71041),
            .in3(N__70363),
            .lcout(),
            .ltout(\quad_counter1.n26_adj_4484_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i13_4_lut_adj_1323_LC_19_9_4 .C_ON=1'b0;
    defparam \quad_counter1.i13_4_lut_adj_1323_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i13_4_lut_adj_1323_LC_19_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i13_4_lut_adj_1323_LC_19_9_4  (
            .in0(N__70213),
            .in1(N__67332),
            .in2(N__67326),
            .in3(N__70523),
            .lcout(\quad_counter1.n28_adj_4488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_2_lut_LC_19_11_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_2_lut_LC_19_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_2_lut_LC_19_11_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2219_2_lut_LC_19_11_0  (
            .in0(N__82008),
            .in1(N__82007),
            .in2(N__67423),
            .in3(N__67323),
            .lcout(\quad_counter1.n3319 ),
            .ltout(),
            .carryin(bfn_19_11_0_),
            .carryout(\quad_counter1.n30634 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_3_lut_LC_19_11_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_3_lut_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_3_lut_LC_19_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_3_lut_LC_19_11_1  (
            .in0(N__81549),
            .in1(N__81548),
            .in2(N__67652),
            .in3(N__67320),
            .lcout(\quad_counter1.n3318 ),
            .ltout(),
            .carryin(\quad_counter1.n30634 ),
            .carryout(\quad_counter1.n30635 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_4_lut_LC_19_11_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_4_lut_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_4_lut_LC_19_11_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2219_4_lut_LC_19_11_2  (
            .in0(N__81522),
            .in1(N__81521),
            .in2(N__67424),
            .in3(N__67317),
            .lcout(\quad_counter1.n3317 ),
            .ltout(),
            .carryin(\quad_counter1.n30635 ),
            .carryout(\quad_counter1.n30636 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_5_lut_LC_19_11_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_5_lut_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_5_lut_LC_19_11_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2219_5_lut_LC_19_11_3  (
            .in0(N__81459),
            .in1(N__81454),
            .in2(N__67427),
            .in3(N__67314),
            .lcout(\quad_counter1.n3316 ),
            .ltout(),
            .carryin(\quad_counter1.n30636 ),
            .carryout(\quad_counter1.n30637 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_6_lut_LC_19_11_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_6_lut_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_6_lut_LC_19_11_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2219_6_lut_LC_19_11_4  (
            .in0(N__70097),
            .in1(N__70098),
            .in2(N__67425),
            .in3(N__67362),
            .lcout(\quad_counter1.n3315 ),
            .ltout(),
            .carryin(\quad_counter1.n30637 ),
            .carryout(\quad_counter1.n30638 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_7_lut_LC_19_11_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_7_lut_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_7_lut_LC_19_11_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2219_7_lut_LC_19_11_5  (
            .in0(N__70050),
            .in1(N__70049),
            .in2(N__67428),
            .in3(N__67359),
            .lcout(\quad_counter1.n3314 ),
            .ltout(),
            .carryin(\quad_counter1.n30638 ),
            .carryout(\quad_counter1.n30639 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_8_lut_LC_19_11_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_8_lut_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_8_lut_LC_19_11_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2219_8_lut_LC_19_11_6  (
            .in0(N__81490),
            .in1(N__81492),
            .in2(N__67426),
            .in3(N__67356),
            .lcout(\quad_counter1.n3313 ),
            .ltout(),
            .carryin(\quad_counter1.n30639 ),
            .carryout(\quad_counter1.n30640 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_9_lut_LC_19_11_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_9_lut_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_9_lut_LC_19_11_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_9_lut_LC_19_11_7  (
            .in0(N__69929),
            .in1(N__69930),
            .in2(N__67653),
            .in3(N__67353),
            .lcout(\quad_counter1.n3312 ),
            .ltout(),
            .carryin(\quad_counter1.n30640 ),
            .carryout(\quad_counter1.n30641 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_10_lut_LC_19_12_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_10_lut_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_10_lut_LC_19_12_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_10_lut_LC_19_12_0  (
            .in0(N__69876),
            .in1(N__69875),
            .in2(N__67642),
            .in3(N__67350),
            .lcout(\quad_counter1.n3311 ),
            .ltout(),
            .carryin(bfn_19_12_0_),
            .carryout(\quad_counter1.n30642 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_11_lut_LC_19_12_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_11_lut_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_11_lut_LC_19_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_11_lut_LC_19_12_1  (
            .in0(N__70536),
            .in1(N__70535),
            .in2(N__67646),
            .in3(N__67347),
            .lcout(\quad_counter1.n3310 ),
            .ltout(),
            .carryin(\quad_counter1.n30642 ),
            .carryout(\quad_counter1.n30643 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_12_lut_LC_19_12_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_12_lut_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_12_lut_LC_19_12_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_12_lut_LC_19_12_2  (
            .in0(N__70485),
            .in1(N__70484),
            .in2(N__67643),
            .in3(N__67344),
            .lcout(\quad_counter1.n3309 ),
            .ltout(),
            .carryin(\quad_counter1.n30643 ),
            .carryout(\quad_counter1.n30644 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_13_lut_LC_19_12_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_13_lut_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_13_lut_LC_19_12_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_13_lut_LC_19_12_3  (
            .in0(N__70428),
            .in1(N__70424),
            .in2(N__67647),
            .in3(N__67341),
            .lcout(\quad_counter1.n3308 ),
            .ltout(),
            .carryin(\quad_counter1.n30644 ),
            .carryout(\quad_counter1.n30645 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_14_lut_LC_19_12_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_14_lut_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_14_lut_LC_19_12_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_14_lut_LC_19_12_4  (
            .in0(N__70373),
            .in1(N__70374),
            .in2(N__67644),
            .in3(N__67338),
            .lcout(\quad_counter1.n3307 ),
            .ltout(),
            .carryin(\quad_counter1.n30645 ),
            .carryout(\quad_counter1.n30646 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_15_lut_LC_19_12_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_15_lut_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_15_lut_LC_19_12_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_15_lut_LC_19_12_5  (
            .in0(N__70326),
            .in1(N__70322),
            .in2(N__67648),
            .in3(N__67335),
            .lcout(\quad_counter1.n3306 ),
            .ltout(),
            .carryin(\quad_counter1.n30646 ),
            .carryout(\quad_counter1.n30647 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_16_lut_LC_19_12_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_16_lut_LC_19_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_16_lut_LC_19_12_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_16_lut_LC_19_12_6  (
            .in0(N__70277),
            .in1(N__70278),
            .in2(N__67645),
            .in3(N__67449),
            .lcout(\quad_counter1.n3305 ),
            .ltout(),
            .carryin(\quad_counter1.n30647 ),
            .carryout(\quad_counter1.n30648 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_17_lut_LC_19_12_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_17_lut_LC_19_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_17_lut_LC_19_12_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_17_lut_LC_19_12_7  (
            .in0(N__70223),
            .in1(N__70224),
            .in2(N__67649),
            .in3(N__67446),
            .lcout(\quad_counter1.n3304 ),
            .ltout(),
            .carryin(\quad_counter1.n30648 ),
            .carryout(\quad_counter1.n30649 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_18_lut_LC_19_13_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_18_lut_LC_19_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_18_lut_LC_19_13_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_18_lut_LC_19_13_0  (
            .in0(N__71049),
            .in1(N__71048),
            .in2(N__67633),
            .in3(N__67443),
            .lcout(\quad_counter1.n3303 ),
            .ltout(),
            .carryin(bfn_19_13_0_),
            .carryout(\quad_counter1.n30650 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_19_lut_LC_19_13_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_19_lut_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_19_lut_LC_19_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_19_lut_LC_19_13_1  (
            .in0(N__70992),
            .in1(N__70991),
            .in2(N__67650),
            .in3(N__67440),
            .lcout(\quad_counter1.n3302 ),
            .ltout(),
            .carryin(\quad_counter1.n30650 ),
            .carryout(\quad_counter1.n30651 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_20_lut_LC_19_13_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_20_lut_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_20_lut_LC_19_13_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_20_lut_LC_19_13_2  (
            .in0(N__70935),
            .in1(N__70934),
            .in2(N__67634),
            .in3(N__67437),
            .lcout(\quad_counter1.n3301 ),
            .ltout(),
            .carryin(\quad_counter1.n30651 ),
            .carryout(\quad_counter1.n30652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_21_lut_LC_19_13_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2219_21_lut_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_21_lut_LC_19_13_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_21_lut_LC_19_13_3  (
            .in0(N__70884),
            .in1(N__70883),
            .in2(N__67651),
            .in3(N__67434),
            .lcout(\quad_counter1.n3300 ),
            .ltout(),
            .carryin(\quad_counter1.n30652 ),
            .carryout(\quad_counter1.n30653 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2219_22_lut_LC_19_13_4 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_2219_22_lut_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2219_22_lut_LC_19_13_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2219_22_lut_LC_19_13_4  (
            .in0(N__70728),
            .in1(N__70727),
            .in2(N__67635),
            .in3(N__67431),
            .lcout(\quad_counter1.n3299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30721_1_lut_LC_19_13_5 .C_ON=1'b0;
    defparam \quad_counter1.i30721_1_lut_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30721_1_lut_LC_19_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter1.i30721_1_lut_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__67588),
            .lcout(\quad_counter1.n36148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i14_4_lut_LC_19_13_6 .C_ON=1'b0;
    defparam \quad_counter1.i14_4_lut_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i14_4_lut_LC_19_13_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i14_4_lut_LC_19_13_6  (
            .in0(N__67383),
            .in1(N__70933),
            .in2(N__67374),
            .in3(N__67662),
            .lcout(\quad_counter1.n3233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__3__5426_LC_19_15_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__3__5426_LC_19_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__3__5426_LC_19_15_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \c0.data_out_frame_12__3__5426_LC_19_15_0  (
            .in0(N__85176),
            .in1(N__83477),
            .in2(N__84561),
            .in3(N__67536),
            .lcout(data_out_frame_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1374_LC_19_15_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1374_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1374_LC_19_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1374_LC_19_15_1  (
            .in0(N__91439),
            .in1(N__91554),
            .in2(N__91367),
            .in3(N__91628),
            .lcout(\c0.n12_adj_4536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i1_LC_19_15_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i1_LC_19_15_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i1_LC_19_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i1_LC_19_15_5  (
            .in0(N__84746),
            .in1(N__67542),
            .in2(_gnd_net_),
            .in3(N__76482),
            .lcout(encoder1_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_19_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_19_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_19_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_19_16_0  (
            .in0(N__76194),
            .in1(N__67535),
            .in2(_gnd_net_),
            .in3(N__96111),
            .lcout(\c0.n11_adj_4517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i15_LC_19_16_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i15_LC_19_16_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i15_LC_19_16_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i15_LC_19_16_1  (
            .in0(N__67509),
            .in1(N__76479),
            .in2(_gnd_net_),
            .in3(N__68168),
            .lcout(encoder1_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97597),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i3_LC_19_16_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i3_LC_19_16_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i3_LC_19_16_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i3_LC_19_16_4  (
            .in0(N__67500),
            .in1(N__76480),
            .in2(_gnd_net_),
            .in3(N__83522),
            .lcout(encoder1_position_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_19_16_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_19_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_19_16_5  (
            .in0(N__96110),
            .in1(N__84273),
            .in2(_gnd_net_),
            .in3(N__67478),
            .lcout(\c0.n11_adj_4507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__1__5428_LC_19_16_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__1__5428_LC_19_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__1__5428_LC_19_16_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_12__1__5428_LC_19_16_6  (
            .in0(N__67479),
            .in1(N__84699),
            .in2(N__85231),
            .in3(N__83054),
            .lcout(data_out_frame_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30754_LC_19_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30754_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_0__bdd_4_lut_30754_LC_19_17_0 .LUT_INIT=16'b1100101011110000;
    LogicCell40 \c0.byte_transmit_counter_0__bdd_4_lut_30754_LC_19_17_0  (
            .in0(N__71756),
            .in1(N__67470),
            .in2(N__96167),
            .in3(N__90372),
            .lcout(),
            .ltout(\c0.n36179_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n36179_bdd_4_lut_LC_19_17_1 .C_ON=1'b0;
    defparam \c0.n36179_bdd_4_lut_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.n36179_bdd_4_lut_LC_19_17_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n36179_bdd_4_lut_LC_19_17_1  (
            .in0(N__90373),
            .in1(N__67673),
            .in2(N__67725),
            .in3(N__67722),
            .lcout(),
            .ltout(\c0.n36182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30669_4_lut_LC_19_17_2 .C_ON=1'b0;
    defparam \c0.i30669_4_lut_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i30669_4_lut_LC_19_17_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.i30669_4_lut_LC_19_17_2  (
            .in0(N__67980),
            .in1(N__90085),
            .in2(N__67701),
            .in3(N__90374),
            .lcout(),
            .ltout(n36098_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_3_lut_4_lut_adj_2067_LC_19_17_3.C_ON=1'b0;
    defparam i24_3_lut_4_lut_adj_2067_LC_19_17_3.SEQ_MODE=4'b0000;
    defparam i24_3_lut_4_lut_adj_2067_LC_19_17_3.LUT_INIT=16'b1011100010101010;
    LogicCell40 i24_3_lut_4_lut_adj_2067_LC_19_17_3 (
            .in0(N__83352),
            .in1(N__90778),
            .in2(N__67698),
            .in3(N__95776),
            .lcout(n10_adj_4821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i9_LC_19_17_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i9_LC_19_17_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i9_LC_19_17_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i9_LC_19_17_4  (
            .in0(N__76474),
            .in1(N__67695),
            .in2(_gnd_net_),
            .in3(N__83058),
            .lcout(encoder1_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97607),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i11_LC_19_17_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i11_LC_19_17_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i11_LC_19_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i11_LC_19_17_6  (
            .in0(N__76473),
            .in1(N__67689),
            .in2(_gnd_net_),
            .in3(N__83466),
            .lcout(encoder1_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97607),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i13_LC_19_17_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i13_LC_19_17_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i13_LC_19_17_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i13_LC_19_17_7  (
            .in0(N__76475),
            .in1(N__67683),
            .in2(_gnd_net_),
            .in3(N__76090),
            .lcout(encoder1_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97607),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__5__5424_LC_19_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__5__5424_LC_19_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__5__5424_LC_19_18_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \c0.data_out_frame_12__5__5424_LC_19_18_0  (
            .in0(N__67994),
            .in1(N__84711),
            .in2(N__85175),
            .in3(N__76083),
            .lcout(data_out_frame_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97619),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__5__5456_LC_19_18_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__5__5456_LC_19_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__5__5456_LC_19_18_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.data_out_frame_8__5__5456_LC_19_18_1  (
            .in0(N__84710),
            .in1(N__85056),
            .in2(N__67677),
            .in3(N__77825),
            .lcout(data_out_frame_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97619),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1482_LC_19_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1482_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1482_LC_19_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1482_LC_19_18_2  (
            .in0(_gnd_net_),
            .in1(N__76082),
            .in2(_gnd_net_),
            .in3(N__77272),
            .lcout(),
            .ltout(\c0.n18357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_19_18_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_19_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_LC_19_18_3  (
            .in0(N__68169),
            .in1(N__83041),
            .in2(N__67770),
            .in3(N__83128),
            .lcout(\c0.n39_adj_4567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__7__5438_LC_19_18_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__7__5438_LC_19_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__7__5438_LC_19_18_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \c0.data_out_frame_10__7__5438_LC_19_18_4  (
            .in0(N__85684),
            .in1(N__67763),
            .in2(N__85174),
            .in3(N__84712),
            .lcout(data_out_frame_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97619),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i16_LC_19_18_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i16_LC_19_18_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i16_LC_19_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i16_LC_19_18_5  (
            .in0(N__76476),
            .in1(N__67749),
            .in2(_gnd_net_),
            .in3(N__79180),
            .lcout(encoder1_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97619),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i14_LC_19_18_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i14_LC_19_18_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i14_LC_19_18_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i14_LC_19_18_6  (
            .in0(N__77285),
            .in1(N__67743),
            .in2(_gnd_net_),
            .in3(N__76478),
            .lcout(encoder1_position_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97619),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i21_LC_19_18_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i21_LC_19_18_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i21_LC_19_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i21_LC_19_18_7  (
            .in0(N__76477),
            .in1(N__67737),
            .in2(_gnd_net_),
            .in3(N__85500),
            .lcout(encoder1_position_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97619),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1449_LC_19_19_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1449_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1449_LC_19_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1449_LC_19_19_0  (
            .in0(N__68029),
            .in1(N__76739),
            .in2(_gnd_net_),
            .in3(N__72003),
            .lcout(\c0.n18689 ),
            .ltout(\c0.n18689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1442_LC_19_19_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1442_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1442_LC_19_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1442_LC_19_19_1  (
            .in0(N__67838),
            .in1(_gnd_net_),
            .in2(N__67731),
            .in3(N__96626),
            .lcout(\c0.n33755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_3_lut_LC_19_19_2 .C_ON=1'b0;
    defparam \c0.i13_3_lut_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_3_lut_LC_19_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i13_3_lut_LC_19_19_2  (
            .in0(N__83467),
            .in1(N__72274),
            .in2(_gnd_net_),
            .in3(N__85683),
            .lcout(),
            .ltout(\c0.n38_adj_4568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_19_19_3 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_19_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_LC_19_19_3  (
            .in0(N__77336),
            .in1(N__67956),
            .in2(N__67728),
            .in3(N__72589),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i29_LC_19_19_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i29_LC_19_19_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i29_LC_19_19_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.count_i0_i29_LC_19_19_4  (
            .in0(N__77936),
            .in1(N__76481),
            .in2(_gnd_net_),
            .in3(N__67962),
            .lcout(encoder1_position_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97633),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_19_19_5 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_19_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_LC_19_19_5  (
            .in0(N__76214),
            .in1(N__72197),
            .in2(N__67839),
            .in3(N__76301),
            .lcout(\c0.n43_adj_4569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i25_LC_19_19_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i25_LC_19_19_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i25_LC_19_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i25_LC_19_19_6  (
            .in0(N__76523),
            .in1(N__67950),
            .in2(_gnd_net_),
            .in3(N__67814),
            .lcout(encoder1_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97633),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i174_LC_19_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i174_LC_19_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i174_LC_19_20_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i174_LC_19_20_0  (
            .in0(N__78421),
            .in1(N__75083),
            .in2(N__67936),
            .in3(N__78573),
            .lcout(\c0.data_in_frame_21_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_19_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_19_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_19_20_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i42_LC_19_20_1  (
            .in0(N__78572),
            .in1(N__75326),
            .in2(N__68296),
            .in3(N__67889),
            .lcout(\c0.data_in_frame_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1441_LC_19_20_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1441_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1441_LC_19_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1441_LC_19_20_3  (
            .in0(N__75922),
            .in1(N__72304),
            .in2(N__67875),
            .in3(N__72099),
            .lcout(\c0.n33400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1443_LC_19_20_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1443_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1443_LC_19_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1443_LC_19_20_4  (
            .in0(N__71928),
            .in1(N__75923),
            .in2(N__76261),
            .in3(N__67789),
            .lcout(\c0.n31673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i18_LC_19_20_5 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i18_LC_19_20_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i18_LC_19_20_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i18_LC_19_20_5  (
            .in0(N__67824),
            .in1(N__76584),
            .in2(_gnd_net_),
            .in3(N__86348),
            .lcout(encoder1_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1448_LC_19_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1448_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1448_LC_19_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1448_LC_19_20_6  (
            .in0(_gnd_net_),
            .in1(N__75826),
            .in2(_gnd_net_),
            .in3(N__67788),
            .lcout(\c0.n33305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1399_LC_19_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1399_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1399_LC_19_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1399_LC_19_20_7  (
            .in0(_gnd_net_),
            .in1(N__68170),
            .in2(_gnd_net_),
            .in3(N__77821),
            .lcout(\c0.n18892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_19_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_19_21_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_19_21_0  (
            .in0(N__68126),
            .in1(N__68366),
            .in2(N__96178),
            .in3(_gnd_net_),
            .lcout(\c0.n11_adj_4576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__4__5425_LC_19_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__4__5425_LC_19_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__4__5425_LC_19_21_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \c0.data_out_frame_12__4__5425_LC_19_21_1  (
            .in0(N__76059),
            .in1(N__84713),
            .in2(N__85275),
            .in3(N__68127),
            .lcout(data_out_frame_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97663),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__3__5482_LC_19_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__3__5482_LC_19_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__3__5482_LC_19_21_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__3__5482_LC_19_21_3  (
            .in0(N__85245),
            .in1(N__84714),
            .in2(N__72158),
            .in3(N__68111),
            .lcout(data_out_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97663),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i1_LC_19_21_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i1_LC_19_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i1_LC_19_21_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i1_LC_19_21_4  (
            .in0(N__72308),
            .in1(N__68097),
            .in2(_gnd_net_),
            .in3(N__77627),
            .lcout(control_mode_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97663),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__4__5481_LC_19_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__4__5481_LC_19_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__4__5481_LC_19_21_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__4__5481_LC_19_21_5  (
            .in0(N__85246),
            .in1(N__84715),
            .in2(N__77559),
            .in3(N__68049),
            .lcout(data_out_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97663),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1440_LC_19_21_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1440_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1440_LC_19_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1440_LC_19_21_7  (
            .in0(N__71871),
            .in1(N__85374),
            .in2(N__96630),
            .in3(N__68018),
            .lcout(\c0.n33615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_19_22_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_19_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_19_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_19_22_0  (
            .in0(N__67995),
            .in1(N__67970),
            .in2(_gnd_net_),
            .in3(N__96155),
            .lcout(\c0.n11_adj_4621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__5__5416_LC_19_22_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__5__5416_LC_19_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__5__5416_LC_19_22_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_13__5__5416_LC_19_22_2  (
            .in0(N__84704),
            .in1(N__85173),
            .in2(N__85743),
            .in3(N__67971),
            .lcout(data_out_frame_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__4__5473_LC_19_22_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__4__5473_LC_19_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__4__5473_LC_19_22_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_6__4__5473_LC_19_22_3  (
            .in0(N__85172),
            .in1(N__84705),
            .in2(N__86205),
            .in3(N__68388),
            .lcout(data_out_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97677),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i1_LC_19_22_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i1_LC_19_22_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i1_LC_19_22_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i1_LC_19_22_4  (
            .in0(N__71790),
            .in1(N__68376),
            .in2(_gnd_net_),
            .in3(N__86111),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__4__5417_LC_19_22_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__4__5417_LC_19_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__4__5417_LC_19_22_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_13__4__5417_LC_19_22_5  (
            .in0(N__85171),
            .in1(N__68367),
            .in2(N__85845),
            .in3(N__84706),
            .lcout(data_out_frame_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97677),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i18_LC_19_22_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i18_LC_19_22_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i18_LC_19_22_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i18_LC_19_22_6  (
            .in0(N__77676),
            .in1(N__68355),
            .in2(_gnd_net_),
            .in3(N__86110),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97677),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i31_LC_19_22_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i31_LC_19_22_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i31_LC_19_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i31_LC_19_22_7  (
            .in0(N__86112),
            .in1(N__68343),
            .in2(_gnd_net_),
            .in3(N__76889),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97677),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i197_LC_19_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i197_LC_19_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i197_LC_19_23_0 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i197_LC_19_23_0  (
            .in0(N__84234),
            .in1(N__68655),
            .in2(N__81174),
            .in3(N__79833),
            .lcout(\c0.data_in_frame_24_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97694),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i7_LC_19_23_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i7_LC_19_23_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i7_LC_19_23_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i7_LC_19_23_1  (
            .in0(N__75930),
            .in1(N__68331),
            .in2(_gnd_net_),
            .in3(N__86108),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97694),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1645_LC_19_23_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1645_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1645_LC_19_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1645_LC_19_23_2  (
            .in0(N__69012),
            .in1(N__69079),
            .in2(_gnd_net_),
            .in3(N__74725),
            .lcout(\c0.n35140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_19_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_19_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_19_23_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i45_LC_19_23_3  (
            .in0(N__68265),
            .in1(N__78559),
            .in2(N__68213),
            .in3(N__84235),
            .lcout(\c0.data_in_frame_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97694),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i13_LC_19_23_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i13_LC_19_23_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i13_LC_19_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i13_LC_19_23_4  (
            .in0(N__86107),
            .in1(N__68193),
            .in2(_gnd_net_),
            .in3(N__77819),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97694),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i179_LC_19_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i179_LC_19_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i179_LC_19_23_5 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i179_LC_19_23_5  (
            .in0(N__80676),
            .in1(N__69013),
            .in2(N__89794),
            .in3(N__72982),
            .lcout(\c0.data_in_frame_22_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97694),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i109_LC_19_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i109_LC_19_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i109_LC_19_23_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i109_LC_19_23_7  (
            .in0(N__68563),
            .in1(N__78558),
            .in2(N__68519),
            .in3(N__84233),
            .lcout(\c0.data_in_frame_13_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97694),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i15_LC_19_24_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i15_LC_19_24_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i15_LC_19_24_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i15_LC_19_24_1  (
            .in0(N__86045),
            .in1(N__68484),
            .in2(_gnd_net_),
            .in3(N__86473),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i195_LC_19_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i195_LC_19_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i195_LC_19_24_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i195_LC_19_24_2  (
            .in0(N__80710),
            .in1(N__81116),
            .in2(N__68475),
            .in3(N__79834),
            .lcout(\c0.data_in_frame_24_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97710),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i10_LC_19_24_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i10_LC_19_24_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i10_LC_19_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i10_LC_19_24_3  (
            .in0(N__86044),
            .in1(N__68445),
            .in2(_gnd_net_),
            .in3(N__72366),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97710),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i8_LC_19_24_4 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i8_LC_19_24_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i8_LC_19_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i8_LC_19_24_4  (
            .in0(N__86046),
            .in1(N__68433),
            .in2(_gnd_net_),
            .in3(N__73221),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_8__4__5457_LC_19_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_8__4__5457_LC_19_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_8__4__5457_LC_19_24_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_8__4__5457_LC_19_24_5  (
            .in0(N__68421),
            .in1(N__85234),
            .in2(N__79248),
            .in3(N__84708),
            .lcout(data_out_frame_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30385_3_lut_LC_19_24_6 .C_ON=1'b0;
    defparam \c0.i30385_3_lut_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30385_3_lut_LC_19_24_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i30385_3_lut_LC_19_24_6  (
            .in0(N__68399),
            .in1(N__68420),
            .in2(_gnd_net_),
            .in3(N__96177),
            .lcout(\c0.n35812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_9__4__5449_LC_19_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_9__4__5449_LC_19_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_9__4__5449_LC_19_24_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_9__4__5449_LC_19_24_7  (
            .in0(N__68400),
            .in1(N__84707),
            .in2(N__85379),
            .in3(N__85235),
            .lcout(data_out_frame_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1686_LC_19_25_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1686_LC_19_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1686_LC_19_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1686_LC_19_25_0  (
            .in0(N__72700),
            .in1(N__69017),
            .in2(_gnd_net_),
            .in3(N__68789),
            .lcout(\c0.n33775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1936_LC_19_25_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1936_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1936_LC_19_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1936_LC_19_25_1  (
            .in0(N__73268),
            .in1(N__68618),
            .in2(N__73353),
            .in3(N__74157),
            .lcout(\c0.n35416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i223_LC_19_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i223_LC_19_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i223_LC_19_25_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i223_LC_19_25_2  (
            .in0(N__78287),
            .in1(N__73671),
            .in2(N__69299),
            .in3(N__79820),
            .lcout(\c0.data_in_frame_27_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i224_LC_19_25_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i224_LC_19_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i224_LC_19_25_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i224_LC_19_25_3  (
            .in0(N__79818),
            .in1(N__80145),
            .in2(N__68738),
            .in3(N__78288),
            .lcout(\c0.data_in_frame_27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97727),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i30_LC_19_25_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i30_LC_19_25_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i30_LC_19_25_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i30_LC_19_25_5  (
            .in0(N__68751),
            .in1(N__86114),
            .in2(_gnd_net_),
            .in3(N__76839),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i205_LC_19_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i205_LC_19_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i205_LC_19_25_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i205_LC_19_25_6  (
            .in0(N__87241),
            .in1(N__84203),
            .in2(N__68714),
            .in3(N__79819),
            .lcout(\c0.data_in_frame_25_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1662_LC_19_25_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1662_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1662_LC_19_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1662_LC_19_25_7  (
            .in0(N__68731),
            .in1(N__68706),
            .in2(_gnd_net_),
            .in3(N__69292),
            .lcout(\c0.n33594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1424_LC_19_26_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1424_LC_19_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1424_LC_19_26_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1424_LC_19_26_1  (
            .in0(N__68662),
            .in1(N__68954),
            .in2(N__69096),
            .in3(N__68912),
            .lcout(\c0.n34009 ),
            .ltout(\c0.n34009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1671_LC_19_26_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1671_LC_19_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1671_LC_19_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1671_LC_19_26_2  (
            .in0(N__79627),
            .in1(N__69109),
            .in2(N__68622),
            .in3(N__73367),
            .lcout(\c0.n31355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i217_LC_19_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i217_LC_19_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i217_LC_19_26_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i217_LC_19_26_4  (
            .in0(N__79821),
            .in1(N__69110),
            .in2(N__78296),
            .in3(N__80926),
            .lcout(\c0.data_in_frame_27_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i215_LC_19_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i215_LC_19_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i215_LC_19_26_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i215_LC_19_26_5  (
            .in0(N__69095),
            .in1(N__73673),
            .in2(N__80361),
            .in3(N__79822),
            .lcout(\c0.data_in_frame_26_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1652_LC_19_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1652_LC_19_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1652_LC_19_26_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1652_LC_19_26_6  (
            .in0(N__69084),
            .in1(N__69045),
            .in2(N__69021),
            .in3(N__74727),
            .lcout(\c0.n33849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_adj_1391_LC_19_26_7 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_adj_1391_LC_19_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_adj_1391_LC_19_26_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_3_lut_4_lut_adj_1391_LC_19_26_7  (
            .in0(N__68973),
            .in1(N__68955),
            .in2(N__68939),
            .in3(N__68913),
            .lcout(\c0.n8_adj_4540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1689_LC_19_27_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1689_LC_19_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1689_LC_19_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1689_LC_19_27_0  (
            .in0(N__73977),
            .in1(N__69129),
            .in2(_gnd_net_),
            .in3(N__74515),
            .lcout(\c0.n20_adj_4698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1691_LC_19_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1691_LC_19_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1691_LC_19_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1691_LC_19_27_1  (
            .in0(_gnd_net_),
            .in1(N__73347),
            .in2(_gnd_net_),
            .in3(N__68821),
            .lcout(\c0.n18596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1925_LC_19_27_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1925_LC_19_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1925_LC_19_27_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1925_LC_19_27_2  (
            .in0(N__73978),
            .in1(N__69130),
            .in2(_gnd_net_),
            .in3(N__68847),
            .lcout(\c0.n6_adj_4756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i240_LC_19_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i240_LC_19_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i240_LC_19_27_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i240_LC_19_27_3  (
            .in0(N__80100),
            .in1(N__78560),
            .in2(N__69315),
            .in3(N__74457),
            .lcout(\c0.data_in_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97763),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1915_LC_19_27_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1915_LC_19_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1915_LC_19_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1915_LC_19_27_4  (
            .in0(N__74152),
            .in1(N__73351),
            .in2(N__68826),
            .in3(N__69351),
            .lcout(),
            .ltout(\c0.n4_adj_4751_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1919_LC_19_27_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1919_LC_19_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1919_LC_19_27_5 .LUT_INIT=16'b1011011111101101;
    LogicCell40 \c0.i2_4_lut_adj_1919_LC_19_27_5  (
            .in0(N__74366),
            .in1(N__69333),
            .in2(N__69327),
            .in3(N__69144),
            .lcout(\c0.n20_adj_4754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1918_LC_19_27_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1918_LC_19_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1918_LC_19_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1918_LC_19_27_6  (
            .in0(N__73979),
            .in1(N__69311),
            .in2(N__69303),
            .in3(N__69279),
            .lcout(\c0.n35250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i209_LC_19_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i209_LC_19_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i209_LC_19_28_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i209_LC_19_28_0  (
            .in0(N__79848),
            .in1(N__80321),
            .in2(N__69248),
            .in3(N__80925),
            .lcout(\c0.data_in_frame_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i203_LC_19_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i203_LC_19_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i203_LC_19_28_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i203_LC_19_28_1  (
            .in0(N__80684),
            .in1(N__87148),
            .in2(N__74043),
            .in3(N__79850),
            .lcout(\c0.data_in_frame_25_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97777),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1627_LC_19_28_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1627_LC_19_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1627_LC_19_28_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1627_LC_19_28_2  (
            .in0(N__73132),
            .in1(N__74038),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n33846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1914_LC_19_28_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1914_LC_19_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1914_LC_19_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1914_LC_19_28_4  (
            .in0(N__69195),
            .in1(N__69186),
            .in2(N__69179),
            .in3(N__69162),
            .lcout(),
            .ltout(\c0.n16_adj_4750_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_adj_1916_LC_19_28_5 .C_ON=1'b0;
    defparam \c0.i8_3_lut_adj_1916_LC_19_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_adj_1916_LC_19_28_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i8_3_lut_adj_1916_LC_19_28_5  (
            .in0(_gnd_net_),
            .in1(N__73133),
            .in2(N__69147),
            .in3(N__74151),
            .lcout(\c0.n18_adj_4752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i221_LC_19_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i221_LC_19_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i221_LC_19_28_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i221_LC_19_28_6  (
            .in0(N__79849),
            .in1(N__78255),
            .in2(N__84255),
            .in3(N__69134),
            .lcout(\c0.data_in_frame_27_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97777),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30704_1_lut_LC_20_2_2 .C_ON=1'b0;
    defparam \quad_counter1.i30704_1_lut_LC_20_2_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30704_1_lut_LC_20_2_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter1.i30704_1_lut_LC_20_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69476),
            .lcout(\quad_counter1.n36131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i8_4_lut_adj_1285_LC_20_3_1 .C_ON=1'b0;
    defparam \quad_counter1.i8_4_lut_adj_1285_LC_20_3_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i8_4_lut_adj_1285_LC_20_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i8_4_lut_adj_1285_LC_20_3_1  (
            .in0(N__69592),
            .in1(N__69774),
            .in2(N__69809),
            .in3(N__69646),
            .lcout(),
            .ltout(\quad_counter1.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1286_LC_20_3_2 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1286_LC_20_3_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1286_LC_20_3_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1286_LC_20_3_2  (
            .in0(N__74574),
            .in1(N__69432),
            .in2(N__69528),
            .in3(N__69835),
            .lcout(\quad_counter1.n2837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23551_2_lut_LC_20_3_3 .C_ON=1'b0;
    defparam \quad_counter1.i23551_2_lut_LC_20_3_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23551_2_lut_LC_20_3_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter1.i23551_2_lut_LC_20_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69424),
            .in3(N__81841),
            .lcout(),
            .ltout(\quad_counter1.n28267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1282_LC_20_3_4 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1282_LC_20_3_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1282_LC_20_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1282_LC_20_3_4  (
            .in0(N__69391),
            .in1(N__69670),
            .in2(N__69438),
            .in3(N__69367),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_4_lut_adj_1283_LC_20_3_5 .C_ON=1'b0;
    defparam \quad_counter1.i1_4_lut_adj_1283_LC_20_3_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_4_lut_adj_1283_LC_20_3_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i1_4_lut_adj_1283_LC_20_3_5  (
            .in0(N__69697),
            .in1(N__69619),
            .in2(N__69435),
            .in3(N__69724),
            .lcout(\quad_counter1.n12_adj_4456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_2_lut_LC_20_4_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_2_lut_LC_20_4_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_2_lut_LC_20_4_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1884_2_lut_LC_20_4_0  (
            .in0(N__81804),
            .in1(N__81803),
            .in2(N__75565),
            .in3(N__69402),
            .lcout(\quad_counter1.n2819 ),
            .ltout(),
            .carryin(bfn_20_4_0_),
            .carryout(\quad_counter1.n30549 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_3_lut_LC_20_4_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_3_lut_LC_20_4_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_3_lut_LC_20_4_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_3_lut_LC_20_4_1  (
            .in0(N__75527),
            .in1(N__75526),
            .in2(N__81632),
            .in3(N__69378),
            .lcout(\quad_counter1.n2818 ),
            .ltout(),
            .carryin(\quad_counter1.n30549 ),
            .carryout(\quad_counter1.n30550 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_4_lut_LC_20_4_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_4_lut_LC_20_4_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_4_lut_LC_20_4_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1884_4_lut_LC_20_4_2  (
            .in0(N__75503),
            .in1(N__75504),
            .in2(N__75566),
            .in3(N__69354),
            .lcout(\quad_counter1.n2817 ),
            .ltout(),
            .carryin(\quad_counter1.n30550 ),
            .carryout(\quad_counter1.n30551 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_5_lut_LC_20_4_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_5_lut_LC_20_4_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_5_lut_LC_20_4_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1884_5_lut_LC_20_4_3  (
            .in0(N__75480),
            .in1(N__75479),
            .in2(N__75569),
            .in3(N__69708),
            .lcout(\quad_counter1.n2816 ),
            .ltout(),
            .carryin(\quad_counter1.n30551 ),
            .carryout(\quad_counter1.n30552 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_6_lut_LC_20_4_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_6_lut_LC_20_4_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_6_lut_LC_20_4_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1884_6_lut_LC_20_4_4  (
            .in0(N__75459),
            .in1(N__75458),
            .in2(N__75567),
            .in3(N__69684),
            .lcout(\quad_counter1.n2815 ),
            .ltout(),
            .carryin(\quad_counter1.n30552 ),
            .carryout(\quad_counter1.n30553 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_7_lut_LC_20_4_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_7_lut_LC_20_4_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_7_lut_LC_20_4_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1884_7_lut_LC_20_4_5  (
            .in0(N__75438),
            .in1(N__75437),
            .in2(N__75570),
            .in3(N__69654),
            .lcout(\quad_counter1.n2814 ),
            .ltout(),
            .carryin(\quad_counter1.n30553 ),
            .carryout(\quad_counter1.n30554 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_8_lut_LC_20_4_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_8_lut_LC_20_4_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_8_lut_LC_20_4_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1884_8_lut_LC_20_4_6  (
            .in0(N__75417),
            .in1(N__75416),
            .in2(N__75568),
            .in3(N__69651),
            .lcout(\quad_counter1.n2813 ),
            .ltout(),
            .carryin(\quad_counter1.n30554 ),
            .carryout(\quad_counter1.n30555 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_9_lut_LC_20_4_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_9_lut_LC_20_4_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_9_lut_LC_20_4_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_9_lut_LC_20_4_7  (
            .in0(N__79362),
            .in1(N__79361),
            .in2(N__81633),
            .in3(N__69630),
            .lcout(\quad_counter1.n2812 ),
            .ltout(),
            .carryin(\quad_counter1.n30555 ),
            .carryout(\quad_counter1.n30556 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_10_lut_LC_20_5_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_10_lut_LC_20_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_10_lut_LC_20_5_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_10_lut_LC_20_5_0  (
            .in0(N__75615),
            .in1(N__75614),
            .in2(N__81624),
            .in3(N__69627),
            .lcout(\quad_counter1.n2811 ),
            .ltout(),
            .carryin(bfn_20_5_0_),
            .carryout(\quad_counter1.n30557 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_11_lut_LC_20_5_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_11_lut_LC_20_5_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_11_lut_LC_20_5_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_11_lut_LC_20_5_1  (
            .in0(N__79266),
            .in1(N__79265),
            .in2(N__81628),
            .in3(N__69624),
            .lcout(\quad_counter1.n2810 ),
            .ltout(),
            .carryin(\quad_counter1.n30557 ),
            .carryout(\quad_counter1.n30558 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_12_lut_LC_20_5_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_12_lut_LC_20_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_12_lut_LC_20_5_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_12_lut_LC_20_5_2  (
            .in0(N__81651),
            .in1(N__81650),
            .in2(N__81625),
            .in3(N__69597),
            .lcout(\quad_counter1.n2809 ),
            .ltout(),
            .carryin(\quad_counter1.n30558 ),
            .carryout(\quad_counter1.n30559 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_13_lut_LC_20_5_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_13_lut_LC_20_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_13_lut_LC_20_5_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_13_lut_LC_20_5_3  (
            .in0(N__79305),
            .in1(N__79304),
            .in2(N__81629),
            .in3(N__69846),
            .lcout(\quad_counter1.n2808 ),
            .ltout(),
            .carryin(\quad_counter1.n30559 ),
            .carryout(\quad_counter1.n30560 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_14_lut_LC_20_5_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_14_lut_LC_20_5_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_14_lut_LC_20_5_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_14_lut_LC_20_5_4  (
            .in0(N__79287),
            .in1(N__79286),
            .in2(N__81626),
            .in3(N__69843),
            .lcout(\quad_counter1.n2807 ),
            .ltout(),
            .carryin(\quad_counter1.n30560 ),
            .carryout(\quad_counter1.n30561 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_15_lut_LC_20_5_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_15_lut_LC_20_5_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_15_lut_LC_20_5_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_15_lut_LC_20_5_5  (
            .in0(N__79325),
            .in1(N__79324),
            .in2(N__81630),
            .in3(N__69813),
            .lcout(\quad_counter1.n2806 ),
            .ltout(),
            .carryin(\quad_counter1.n30561 ),
            .carryout(\quad_counter1.n30562 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_16_lut_LC_20_5_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1884_16_lut_LC_20_5_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_16_lut_LC_20_5_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_16_lut_LC_20_5_6  (
            .in0(N__81678),
            .in1(N__81677),
            .in2(N__81627),
            .in3(N__69780),
            .lcout(\quad_counter1.n2805 ),
            .ltout(),
            .carryin(\quad_counter1.n30562 ),
            .carryout(\quad_counter1.n30563 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1884_17_lut_LC_20_5_7 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1884_17_lut_LC_20_5_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1884_17_lut_LC_20_5_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1884_17_lut_LC_20_5_7  (
            .in0(N__79343),
            .in1(N__79344),
            .in2(N__81631),
            .in3(N__69777),
            .lcout(\quad_counter1.n2804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_3_lut_adj_1312_LC_20_6_5 .C_ON=1'b0;
    defparam \quad_counter1.i1_3_lut_adj_1312_LC_20_6_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_3_lut_adj_1312_LC_20_6_5 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \quad_counter1.i1_3_lut_adj_1312_LC_20_6_5  (
            .in0(_gnd_net_),
            .in1(N__81970),
            .in2(N__70144),
            .in3(N__70168),
            .lcout(\quad_counter1.n7_adj_4478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i13_4_lut_adj_1317_LC_20_7_0 .C_ON=1'b0;
    defparam \quad_counter1.i13_4_lut_adj_1317_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i13_4_lut_adj_1317_LC_20_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i13_4_lut_adj_1317_LC_20_7_0  (
            .in0(N__70552),
            .in1(N__70194),
            .in2(N__70447),
            .in3(N__69753),
            .lcout(\quad_counter1.n3134 ),
            .ltout(\quad_counter1.n3134_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30725_1_lut_LC_20_7_1 .C_ON=1'b0;
    defparam \quad_counter1.i30725_1_lut_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30725_1_lut_LC_20_7_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30725_1_lut_LC_20_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69747),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1313_LC_20_7_3 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1313_LC_20_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1313_LC_20_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1313_LC_20_7_3  (
            .in0(N__70069),
            .in1(N__69744),
            .in2(N__70021),
            .in3(N__69738),
            .lcout(),
            .ltout(\quad_counter1.n34587_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i8_4_lut_adj_1315_LC_20_7_4 .C_ON=1'b0;
    defparam \quad_counter1.i8_4_lut_adj_1315_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i8_4_lut_adj_1315_LC_20_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i8_4_lut_adj_1315_LC_20_7_4  (
            .in0(N__71062),
            .in1(N__70849),
            .in2(N__70197),
            .in3(N__69895),
            .lcout(\quad_counter1.n22_adj_4481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_2_lut_LC_20_8_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_2_lut_LC_20_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_2_lut_LC_20_8_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2152_2_lut_LC_20_8_0  (
            .in0(N__81972),
            .in1(N__81971),
            .in2(N__69967),
            .in3(N__70188),
            .lcout(\quad_counter1.n3219 ),
            .ltout(),
            .carryin(bfn_20_8_0_),
            .carryout(\quad_counter1.n30615 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_3_lut_LC_20_8_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_3_lut_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_3_lut_LC_20_8_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_3_lut_LC_20_8_1  (
            .in0(N__70185),
            .in1(N__70181),
            .in2(N__70777),
            .in3(N__70155),
            .lcout(\quad_counter1.n3218 ),
            .ltout(),
            .carryin(\quad_counter1.n30615 ),
            .carryout(\quad_counter1.n30616 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_4_lut_LC_20_8_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_4_lut_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_4_lut_LC_20_8_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2152_4_lut_LC_20_8_2  (
            .in0(N__70152),
            .in1(N__70151),
            .in2(N__69968),
            .in3(N__70125),
            .lcout(\quad_counter1.n3217 ),
            .ltout(),
            .carryin(\quad_counter1.n30616 ),
            .carryout(\quad_counter1.n30617 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_5_lut_LC_20_8_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_5_lut_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_5_lut_LC_20_8_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2152_5_lut_LC_20_8_3  (
            .in0(N__70122),
            .in1(N__70121),
            .in2(N__69971),
            .in3(N__70074),
            .lcout(\quad_counter1.n3216 ),
            .ltout(),
            .carryin(\quad_counter1.n30617 ),
            .carryout(\quad_counter1.n30618 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_6_lut_LC_20_8_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_6_lut_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_6_lut_LC_20_8_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2152_6_lut_LC_20_8_4  (
            .in0(N__70071),
            .in1(N__70070),
            .in2(N__69969),
            .in3(N__70026),
            .lcout(\quad_counter1.n3215 ),
            .ltout(),
            .carryin(\quad_counter1.n30618 ),
            .carryout(\quad_counter1.n30619 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_7_lut_LC_20_8_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_7_lut_LC_20_8_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_7_lut_LC_20_8_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2152_7_lut_LC_20_8_5  (
            .in0(N__70022),
            .in1(N__70023),
            .in2(N__69972),
            .in3(N__69996),
            .lcout(\quad_counter1.n3214 ),
            .ltout(),
            .carryin(\quad_counter1.n30619 ),
            .carryout(\quad_counter1.n30620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_8_lut_LC_20_8_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_8_lut_LC_20_8_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_8_lut_LC_20_8_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2152_8_lut_LC_20_8_6  (
            .in0(N__69993),
            .in1(N__69992),
            .in2(N__69970),
            .in3(N__69906),
            .lcout(\quad_counter1.n3213 ),
            .ltout(),
            .carryin(\quad_counter1.n30620 ),
            .carryout(\quad_counter1.n30621 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_9_lut_LC_20_8_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_9_lut_LC_20_8_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_9_lut_LC_20_8_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_9_lut_LC_20_8_7  (
            .in0(N__69903),
            .in1(N__69902),
            .in2(N__70778),
            .in3(N__70563),
            .lcout(\quad_counter1.n3212 ),
            .ltout(),
            .carryin(\quad_counter1.n30621 ),
            .carryout(\quad_counter1.n30622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_10_lut_LC_20_9_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_10_lut_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_10_lut_LC_20_9_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_10_lut_LC_20_9_0  (
            .in0(N__70560),
            .in1(N__70559),
            .in2(N__70813),
            .in3(N__70512),
            .lcout(\quad_counter1.n3211 ),
            .ltout(),
            .carryin(bfn_20_9_0_),
            .carryout(\quad_counter1.n30623 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_11_lut_LC_20_9_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_11_lut_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_11_lut_LC_20_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_11_lut_LC_20_9_1  (
            .in0(N__70509),
            .in1(N__70508),
            .in2(N__70817),
            .in3(N__70458),
            .lcout(\quad_counter1.n3210 ),
            .ltout(),
            .carryin(\quad_counter1.n30623 ),
            .carryout(\quad_counter1.n30624 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_12_lut_LC_20_9_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_12_lut_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_12_lut_LC_20_9_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_12_lut_LC_20_9_2  (
            .in0(N__70455),
            .in1(N__70454),
            .in2(N__70814),
            .in3(N__70404),
            .lcout(\quad_counter1.n3209 ),
            .ltout(),
            .carryin(\quad_counter1.n30624 ),
            .carryout(\quad_counter1.n30625 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_13_lut_LC_20_9_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_13_lut_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_13_lut_LC_20_9_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_13_lut_LC_20_9_3  (
            .in0(N__70401),
            .in1(N__70400),
            .in2(N__70818),
            .in3(N__70350),
            .lcout(\quad_counter1.n3208 ),
            .ltout(),
            .carryin(\quad_counter1.n30625 ),
            .carryout(\quad_counter1.n30626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_14_lut_LC_20_9_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_14_lut_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_14_lut_LC_20_9_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_14_lut_LC_20_9_4  (
            .in0(N__70347),
            .in1(N__70346),
            .in2(N__70815),
            .in3(N__70302),
            .lcout(\quad_counter1.n3207 ),
            .ltout(),
            .carryin(\quad_counter1.n30626 ),
            .carryout(\quad_counter1.n30627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_15_lut_LC_20_9_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_15_lut_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_15_lut_LC_20_9_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_15_lut_LC_20_9_5  (
            .in0(N__70299),
            .in1(N__70298),
            .in2(N__70819),
            .in3(N__70251),
            .lcout(\quad_counter1.n3206 ),
            .ltout(),
            .carryin(\quad_counter1.n30627 ),
            .carryout(\quad_counter1.n30628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_16_lut_LC_20_9_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_16_lut_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_16_lut_LC_20_9_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_16_lut_LC_20_9_6  (
            .in0(N__70248),
            .in1(N__70247),
            .in2(N__70816),
            .in3(N__70200),
            .lcout(\quad_counter1.n3205 ),
            .ltout(),
            .carryin(\quad_counter1.n30628 ),
            .carryout(\quad_counter1.n30629 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_17_lut_LC_20_9_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_17_lut_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_17_lut_LC_20_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_17_lut_LC_20_9_7  (
            .in0(N__71070),
            .in1(N__71069),
            .in2(N__70820),
            .in3(N__71022),
            .lcout(\quad_counter1.n3204 ),
            .ltout(),
            .carryin(\quad_counter1.n30629 ),
            .carryout(\quad_counter1.n30630 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_18_lut_LC_20_10_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_18_lut_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_18_lut_LC_20_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_18_lut_LC_20_10_0  (
            .in0(N__71019),
            .in1(N__71015),
            .in2(N__70833),
            .in3(N__70968),
            .lcout(\quad_counter1.n3203 ),
            .ltout(),
            .carryin(bfn_20_10_0_),
            .carryout(\quad_counter1.n30631 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_19_lut_LC_20_10_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_19_lut_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_19_lut_LC_20_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_19_lut_LC_20_10_1  (
            .in0(N__70965),
            .in1(N__70961),
            .in2(N__70835),
            .in3(N__70914),
            .lcout(\quad_counter1.n3202 ),
            .ltout(),
            .carryin(\quad_counter1.n30631 ),
            .carryout(\quad_counter1.n30632 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_20_lut_LC_20_10_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2152_20_lut_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_20_lut_LC_20_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_20_lut_LC_20_10_2  (
            .in0(N__70911),
            .in1(N__70910),
            .in2(N__70834),
            .in3(N__70860),
            .lcout(\quad_counter1.n3201 ),
            .ltout(),
            .carryin(\quad_counter1.n30632 ),
            .carryout(\quad_counter1.n30633 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2152_21_lut_LC_20_10_3 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_2152_21_lut_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2152_21_lut_LC_20_10_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2152_21_lut_LC_20_10_3  (
            .in0(N__70856),
            .in1(N__70857),
            .in2(N__70836),
            .in3(N__70731),
            .lcout(\quad_counter1.n3200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_2_lut_LC_20_11_0 .C_ON=1'b0;
    defparam \quad_counter0.i2_2_lut_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_2_lut_LC_20_11_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter0.i2_2_lut_LC_20_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__70704),
            .in3(N__70677),
            .lcout(\quad_counter0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i2_2_lut_adj_1209_LC_20_11_1 .C_ON=1'b0;
    defparam \quad_counter0.i2_2_lut_adj_1209_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i2_2_lut_adj_1209_LC_20_11_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter0.i2_2_lut_adj_1209_LC_20_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__70629),
            .in3(N__70594),
            .lcout(\quad_counter0.n8_adj_4394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_adj_1268_LC_20_11_4 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_adj_1268_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_adj_1268_LC_20_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \quad_counter1.i2_2_lut_adj_1268_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__87747),
            .in2(_gnd_net_),
            .in3(N__87834),
            .lcout(\quad_counter1.n8_adj_4444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i3_LC_20_11_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_20_11_7 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_20_11_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_20_11_7  (
            .in0(N__71410),
            .in1(N__71233),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97564),
            .ce(),
            .sr(N__71211));
    defparam \quad_counter1.i5_4_lut_LC_20_12_0 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_LC_20_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i5_4_lut_LC_20_12_0  (
            .in0(N__82256),
            .in1(N__71196),
            .in2(N__71181),
            .in3(N__82283),
            .lcout(\quad_counter1.n35603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_LC_20_12_1 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_LC_20_12_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter1.i2_2_lut_LC_20_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__82234),
            .in3(N__82310),
            .lcout(\quad_counter1.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1270_LC_20_12_2 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1270_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1270_LC_20_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1270_LC_20_12_2  (
            .in0(N__87777),
            .in1(N__71190),
            .in2(N__88050),
            .in3(N__87807),
            .lcout(),
            .ltout(\quad_counter1.n35309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1271_LC_20_12_3 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1271_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1271_LC_20_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1271_LC_20_12_3  (
            .in0(N__88179),
            .in1(N__88149),
            .in2(N__71184),
            .in3(N__88242),
            .lcout(\quad_counter1.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_3_lut_LC_20_12_6 .C_ON=1'b0;
    defparam \quad_counter1.i1_3_lut_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_3_lut_LC_20_12_6 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \quad_counter1.i1_3_lut_LC_20_12_6  (
            .in0(N__82417),
            .in1(_gnd_net_),
            .in2(N__82345),
            .in3(N__82367),
            .lcout(\quad_counter1.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_LC_20_13_3 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_LC_20_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i12_4_lut_LC_20_13_3  (
            .in0(N__82916),
            .in1(N__82889),
            .in2(N__82552),
            .in3(N__82693),
            .lcout(\quad_counter1.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_LC_20_13_4 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_LC_20_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_LC_20_13_4  (
            .in0(N__82487),
            .in1(N__83000),
            .in2(N__82609),
            .in3(N__82631),
            .lcout(\quad_counter1.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_LC_20_13_5 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_LC_20_13_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_LC_20_13_5  (
            .in0(N__82574),
            .in1(N__82862),
            .in2(N__82666),
            .in3(N__82720),
            .lcout(\quad_counter1.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_20_14_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_20_14_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_20_14_4 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_20_14_4  (
            .in0(N__71609),
            .in1(N__71172),
            .in2(N__71155),
            .in3(N__71694),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97589),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_LC_20_14_6 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_LC_20_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i9_4_lut_LC_20_14_6  (
            .in0(N__82943),
            .in1(N__71595),
            .in2(N__82978),
            .in3(N__82522),
            .lcout(\quad_counter1.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_20_15_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_20_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_20_15_6  (
            .in0(N__76176),
            .in1(N__90420),
            .in2(_gnd_net_),
            .in3(N__96112),
            .lcout(),
            .ltout(\c0.n26_adj_4625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30399_4_lut_LC_20_15_7 .C_ON=1'b0;
    defparam \c0.i30399_4_lut_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30399_4_lut_LC_20_15_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.i30399_4_lut_LC_20_15_7  (
            .in0(N__90870),
            .in1(N__71586),
            .in2(N__71571),
            .in3(N__90759),
            .lcout(n35826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_7__1__5468_LC_20_16_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_7__1__5468_LC_20_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_7__1__5468_LC_20_16_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.data_out_frame_7__1__5468_LC_20_16_0  (
            .in0(N__84697),
            .in1(N__85151),
            .in2(N__71541),
            .in3(N__83272),
            .lcout(data_out_frame_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97608),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i5_LC_20_16_2 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i5_LC_20_16_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i5_LC_20_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i5_LC_20_16_2  (
            .in0(N__76543),
            .in1(N__71550),
            .in2(_gnd_net_),
            .in3(N__85716),
            .lcout(encoder1_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_20_16_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_20_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_20_16_4  (
            .in0(N__71537),
            .in1(N__72222),
            .in2(_gnd_net_),
            .in3(N__96113),
            .lcout(),
            .ltout(\c0.n5_adj_4505_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30403_4_lut_LC_20_16_5 .C_ON=1'b0;
    defparam \c0.i30403_4_lut_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i30403_4_lut_LC_20_16_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.i30403_4_lut_LC_20_16_5  (
            .in0(N__71829),
            .in1(N__90100),
            .in2(N__71529),
            .in3(N__90344),
            .lcout(),
            .ltout(\c0.n35830_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30405_4_lut_LC_20_16_6 .C_ON=1'b0;
    defparam \c0.i30405_4_lut_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30405_4_lut_LC_20_16_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.i30405_4_lut_LC_20_16_6  (
            .in0(N__90872),
            .in1(N__90760),
            .in2(N__71526),
            .in3(N__93861),
            .lcout(n35832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_10__5__5440_LC_20_16_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_10__5__5440_LC_20_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_10__5__5440_LC_20_16_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_10__5__5440_LC_20_16_7  (
            .in0(N__85150),
            .in1(N__84698),
            .in2(N__77952),
            .in3(N__71757),
            .lcout(data_out_frame_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30589_3_lut_LC_20_17_0 .C_ON=1'b0;
    defparam \c0.i30589_3_lut_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i30589_3_lut_LC_20_17_0 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \c0.i30589_3_lut_LC_20_17_0  (
            .in0(N__96114),
            .in1(N__71852),
            .in2(_gnd_net_),
            .in3(N__90101),
            .lcout(),
            .ltout(\c0.n36016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30400_4_lut_LC_20_17_1 .C_ON=1'b0;
    defparam \c0.i30400_4_lut_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i30400_4_lut_LC_20_17_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i30400_4_lut_LC_20_17_1  (
            .in0(N__90102),
            .in1(N__71901),
            .in2(N__71745),
            .in3(N__90376),
            .lcout(),
            .ltout(\c0.n35827_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30402_4_lut_LC_20_17_2 .C_ON=1'b0;
    defparam \c0.i30402_4_lut_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i30402_4_lut_LC_20_17_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.i30402_4_lut_LC_20_17_2  (
            .in0(N__90767),
            .in1(N__90873),
            .in2(N__71742),
            .in3(N__83553),
            .lcout(n35829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_12__2__5427_LC_20_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_12__2__5427_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_12__2__5427_LC_20_17_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_12__2__5427_LC_20_17_3  (
            .in0(N__85278),
            .in1(N__84692),
            .in2(N__83137),
            .in3(N__89180),
            .lcout(data_out_frame_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__1__5484_LC_20_17_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__1__5484_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__1__5484_LC_20_17_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__1__5484_LC_20_17_4  (
            .in0(N__84691),
            .in1(N__85280),
            .in2(N__72315),
            .in3(N__71841),
            .lcout(data_out_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97620),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i8_LC_20_17_6 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i8_LC_20_17_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i8_LC_20_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i8_LC_20_17_6  (
            .in0(N__76579),
            .in1(N__71727),
            .in2(_gnd_net_),
            .in3(N__75873),
            .lcout(encoder1_position_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__0__5485_LC_20_17_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__0__5485_LC_20_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__0__5485_LC_20_17_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__0__5485_LC_20_17_7  (
            .in0(N__85279),
            .in1(N__84693),
            .in2(N__83190),
            .in3(N__71717),
            .lcout(data_out_frame_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97620),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i20_LC_20_18_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i20_LC_20_18_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i20_LC_20_18_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \quad_counter1.count_i0_i20_LC_20_18_0  (
            .in0(N__76644),
            .in1(N__71703),
            .in2(N__76590),
            .in3(_gnd_net_),
            .lcout(encoder1_position_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97634),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1485_LC_20_18_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1485_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1485_LC_20_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1485_LC_20_18_1  (
            .in0(N__75863),
            .in1(N__77901),
            .in2(_gnd_net_),
            .in3(N__76235),
            .lcout(\c0.n33795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_20_18_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_20_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_20_18_3  (
            .in0(N__96160),
            .in1(N__71919),
            .in2(_gnd_net_),
            .in3(N__71816),
            .lcout(\c0.n5_adj_4653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_20_18_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_20_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_LC_20_18_4  (
            .in0(N__85391),
            .in1(N__71891),
            .in2(_gnd_net_),
            .in3(N__72009),
            .lcout(\c0.n14_adj_4562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_5__7__5478_LC_20_18_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_5__7__5478_LC_20_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_5__7__5478_LC_20_18_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_5__7__5478_LC_20_18_5  (
            .in0(N__85228),
            .in1(N__84701),
            .in2(N__72468),
            .in3(N__71853),
            .lcout(data_out_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97634),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30661_3_lut_LC_20_18_6 .C_ON=1'b0;
    defparam \c0.i30661_3_lut_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30661_3_lut_LC_20_18_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \c0.i30661_3_lut_LC_20_18_6  (
            .in0(N__90075),
            .in1(N__96159),
            .in2(_gnd_net_),
            .in3(N__71840),
            .lcout(\c0.n36090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__7__5470_LC_20_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__7__5470_LC_20_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__7__5470_LC_20_18_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_6__7__5470_LC_20_18_7  (
            .in0(N__85229),
            .in1(N__84702),
            .in2(N__76914),
            .in3(N__71817),
            .lcout(data_out_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97634),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1468_LC_20_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1468_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1468_LC_20_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1468_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(N__71800),
            .in2(_gnd_net_),
            .in3(N__76904),
            .lcout(\c0.n33892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1469_LC_20_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1469_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1469_LC_20_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1469_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(N__85455),
            .in2(_gnd_net_),
            .in3(N__85490),
            .lcout(),
            .ltout(\c0.n33503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_20_19_3 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_20_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_LC_20_19_3  (
            .in0(N__76635),
            .in1(N__86515),
            .in2(N__71769),
            .in3(N__76738),
            .lcout(),
            .ltout(\c0.n41_adj_4571_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_LC_20_19_4 .C_ON=1'b0;
    defparam \c0.i24_4_lut_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_LC_20_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i24_4_lut_LC_20_19_4  (
            .in0(N__72108),
            .in1(N__71766),
            .in2(N__71760),
            .in3(N__76314),
            .lcout(\c0.n31401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1483_LC_20_19_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1483_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1483_LC_20_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1483_LC_20_19_5  (
            .in0(N__72379),
            .in1(N__79243),
            .in2(_gnd_net_),
            .in3(N__86292),
            .lcout(),
            .ltout(\c0.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_20_19_6 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_20_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_LC_20_19_6  (
            .in0(N__76058),
            .in1(N__71943),
            .in2(N__72117),
            .in3(N__72114),
            .lcout(\c0.n45_adj_4572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1460_LC_20_19_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1460_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1460_LC_20_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1460_LC_20_19_7  (
            .in0(N__72330),
            .in1(N__83271),
            .in2(N__72078),
            .in3(N__76905),
            .lcout(\c0.n18218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1467_LC_20_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1467_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1467_LC_20_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1467_LC_20_20_0  (
            .in0(_gnd_net_),
            .in1(N__77677),
            .in2(_gnd_net_),
            .in3(N__72001),
            .lcout(),
            .ltout(\c0.n33314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_20_20_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_20_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_20_20_1  (
            .in0(N__76352),
            .in1(N__72153),
            .in2(N__72102),
            .in3(N__72098),
            .lcout(),
            .ltout(\c0.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_20_20_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_20_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_20_20_2  (
            .in0(N__76673),
            .in1(N__72464),
            .in2(N__72081),
            .in3(N__72015),
            .lcout(\c0.n26_adj_4559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_LC_20_20_3 .C_ON=1'b0;
    defparam \c0.i4_2_lut_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_LC_20_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i4_2_lut_LC_20_20_3  (
            .in0(_gnd_net_),
            .in1(N__72073),
            .in2(_gnd_net_),
            .in3(N__77409),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1750_LC_20_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1750_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1750_LC_20_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1750_LC_20_20_4  (
            .in0(N__72152),
            .in1(N__77678),
            .in2(_gnd_net_),
            .in3(N__72002),
            .lcout(\c0.n33765 ),
            .ltout(\c0.n33765_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_20_20_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_20_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_20_20_5  (
            .in0(N__72329),
            .in1(N__72486),
            .in2(N__71937),
            .in3(N__71934),
            .lcout(\c0.n33493 ),
            .ltout(\c0.n33493_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_20_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1752_LC_20_20_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1752_LC_20_20_6  (
            .in0(N__72154),
            .in1(_gnd_net_),
            .in2(N__72333),
            .in3(N__72203),
            .lcout(\c0.n6_adj_4560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1711_LC_20_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1711_LC_20_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1711_LC_20_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1711_LC_20_20_7  (
            .in0(N__79065),
            .in1(N__72660),
            .in2(_gnd_net_),
            .in3(N__78037),
            .lcout(\c0.n33389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1458_LC_20_21_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1458_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1458_LC_20_21_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1458_LC_20_21_0  (
            .in0(N__72303),
            .in1(_gnd_net_),
            .in2(N__83186),
            .in3(N__72201),
            .lcout(\c0.n33749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_1__I_0_2_lut_LC_20_21_1 .C_ON=1'b0;
    defparam \c0.control_mode_1__I_0_2_lut_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.control_mode_1__I_0_2_lut_LC_20_21_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.control_mode_1__I_0_2_lut_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(N__83179),
            .in2(_gnd_net_),
            .in3(N__72302),
            .lcout(\c0.data_out_frame_29__7__N_734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1446_LC_20_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1446_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1446_LC_20_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1446_LC_20_21_2  (
            .in0(_gnd_net_),
            .in1(N__76791),
            .in2(_gnd_net_),
            .in3(N__72460),
            .lcout(),
            .ltout(\c0.n33432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1451_LC_20_21_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1451_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1451_LC_20_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1451_LC_20_21_3  (
            .in0(N__76334),
            .in1(N__72279),
            .in2(N__72237),
            .in3(N__72624),
            .lcout(\c0.n18523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i31_LC_20_21_4 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i31_LC_20_21_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i31_LC_20_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i31_LC_20_21_4  (
            .in0(N__76572),
            .in1(N__72234),
            .in2(_gnd_net_),
            .in3(N__85674),
            .lcout(encoder1_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_6__1__5476_LC_20_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_6__1__5476_LC_20_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_6__1__5476_LC_20_21_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_6__1__5476_LC_20_21_5  (
            .in0(N__85274),
            .in1(N__84709),
            .in2(N__73098),
            .in3(N__72221),
            .lcout(data_out_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_3__I_0_2_lut_LC_20_21_6 .C_ON=1'b0;
    defparam \c0.control_mode_3__I_0_2_lut_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.control_mode_3__I_0_2_lut_LC_20_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.control_mode_3__I_0_2_lut_LC_20_21_6  (
            .in0(_gnd_net_),
            .in1(N__72202),
            .in2(_gnd_net_),
            .in3(N__72159),
            .lcout(\c0.data_out_frame_29__7__N_738 ),
            .ltout(\c0.data_out_frame_29__7__N_738_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1445_LC_20_21_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1445_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1445_LC_20_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1445_LC_20_21_7  (
            .in0(N__73231),
            .in1(N__72623),
            .in2(N__72495),
            .in3(N__72492),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1464_LC_20_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1464_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1464_LC_20_22_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1464_LC_20_22_0  (
            .in0(N__86352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86412),
            .lcout(\c0.n33579 ),
            .ltout(\c0.n33579_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1416_LC_20_22_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1416_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1416_LC_20_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1416_LC_20_22_1  (
            .in0(N__86525),
            .in1(N__77781),
            .in2(N__72480),
            .in3(N__83533),
            .lcout(\c0.n10_adj_4547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1754_LC_20_22_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1754_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1754_LC_20_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1754_LC_20_22_2  (
            .in0(N__76788),
            .in1(N__72454),
            .in2(N__72588),
            .in3(N__78036),
            .lcout(\c0.n17510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i7_LC_20_22_4 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i7_LC_20_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i7_LC_20_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.control_mode_i0_i7_LC_20_22_4  (
            .in0(N__77628),
            .in1(N__72456),
            .in2(_gnd_net_),
            .in3(N__77184),
            .lcout(control_mode_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97695),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i2_LC_20_22_5 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i2_LC_20_22_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i2_LC_20_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i2_LC_20_22_5  (
            .in0(N__86113),
            .in1(N__72477),
            .in2(_gnd_net_),
            .in3(N__83316),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97695),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1463_LC_20_22_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1463_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1463_LC_20_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1463_LC_20_22_6  (
            .in0(N__77121),
            .in1(N__72455),
            .in2(N__85922),
            .in3(N__73080),
            .lcout(\c0.n18181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i5_LC_20_22_7 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i5_LC_20_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i5_LC_20_22_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.control_mode_i0_i5_LC_20_22_7  (
            .in0(N__72429),
            .in1(N__76789),
            .in2(_gnd_net_),
            .in3(N__77629),
            .lcout(control_mode_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97695),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1710_LC_20_23_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1710_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1710_LC_20_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1710_LC_20_23_0  (
            .in0(N__78025),
            .in1(N__72362),
            .in2(N__73090),
            .in3(N__72663),
            .lcout(\c0.n33280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i17_LC_20_23_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i17_LC_20_23_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i17_LC_20_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i17_LC_20_23_2  (
            .in0(N__86109),
            .in1(N__72684),
            .in2(_gnd_net_),
            .in3(N__83267),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97711),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1758_LC_20_23_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1758_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1758_LC_20_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1758_LC_20_23_3  (
            .in0(N__79152),
            .in1(N__85783),
            .in2(N__72672),
            .in3(N__85676),
            .lcout(\c0.n31423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1392_LC_20_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1392_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1392_LC_20_23_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1392_LC_20_23_4  (
            .in0(_gnd_net_),
            .in1(N__77948),
            .in2(_gnd_net_),
            .in3(N__86272),
            .lcout(\c0.n6_adj_4541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1712_LC_20_23_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1712_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1712_LC_20_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1712_LC_20_23_6  (
            .in0(N__78024),
            .in1(N__72662),
            .in2(N__76746),
            .in3(N__77553),
            .lcout(\c0.n33414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1470_LC_20_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1470_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1470_LC_20_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1470_LC_20_23_7  (
            .in0(_gnd_net_),
            .in1(N__85782),
            .in2(_gnd_net_),
            .in3(N__85675),
            .lcout(\c0.n33807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i23_LC_20_24_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i23_LC_20_24_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i23_LC_20_24_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i23_LC_20_24_0  (
            .in0(N__86104),
            .in1(N__72612),
            .in2(_gnd_net_),
            .in3(N__72575),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i9_LC_20_24_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i9_LC_20_24_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i9_LC_20_24_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter0.count_i0_i9_LC_20_24_1  (
            .in0(N__77428),
            .in1(N__86106),
            .in2(_gnd_net_),
            .in3(N__72543),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i16_LC_20_24_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i16_LC_20_24_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i16_LC_20_24_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i16_LC_20_24_2  (
            .in0(N__86103),
            .in1(N__72531),
            .in2(_gnd_net_),
            .in3(N__86407),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i181_LC_20_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i181_LC_20_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i181_LC_20_24_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i181_LC_20_24_3  (
            .in0(N__89712),
            .in1(N__84236),
            .in2(N__72515),
            .in3(N__73036),
            .lcout(\c0.data_in_frame_22_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i235_LC_20_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i235_LC_20_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i235_LC_20_24_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i235_LC_20_24_4  (
            .in0(N__78505),
            .in1(N__80718),
            .in2(N__74455),
            .in3(N__73269),
            .lcout(\c0.data_in_frame_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i234_LC_20_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i234_LC_20_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i234_LC_20_24_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i234_LC_20_24_5  (
            .in0(N__75369),
            .in1(N__74441),
            .in2(N__73256),
            .in3(N__78506),
            .lcout(\c0.data_in_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1480_LC_20_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1480_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1480_LC_20_24_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1480_LC_20_24_6  (
            .in0(_gnd_net_),
            .in1(N__77427),
            .in2(_gnd_net_),
            .in3(N__73211),
            .lcout(\c0.n33772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i4_LC_20_24_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i4_LC_20_24_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i4_LC_20_24_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i4_LC_20_24_7  (
            .in0(N__73185),
            .in1(N__86105),
            .in2(_gnd_net_),
            .in3(N__85361),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97729),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i201_LC_20_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i201_LC_20_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i201_LC_20_25_0 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i201_LC_20_25_0  (
            .in0(N__80876),
            .in1(N__74173),
            .in2(N__87303),
            .in3(N__79862),
            .lcout(\c0.data_in_frame_25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i212_LC_20_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i212_LC_20_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i212_LC_20_25_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i212_LC_20_25_1  (
            .in0(N__79859),
            .in1(N__80265),
            .in2(N__78996),
            .in3(N__73162),
            .lcout(\c0.data_in_frame_26_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i204_LC_20_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i204_LC_20_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i204_LC_20_25_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i204_LC_20_25_2  (
            .in0(N__73131),
            .in1(N__78991),
            .in2(N__87304),
            .in3(N__79863),
            .lcout(\c0.data_in_frame_25_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i25_LC_20_25_3 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i25_LC_20_25_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i25_LC_20_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter0.count_i0_i25_LC_20_25_3  (
            .in0(N__73110),
            .in1(N__86115),
            .in2(_gnd_net_),
            .in3(N__73079),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i180_LC_20_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i180_LC_20_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i180_LC_20_25_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i180_LC_20_25_4  (
            .in0(N__89774),
            .in1(N__78990),
            .in2(N__73046),
            .in3(N__72704),
            .lcout(\c0.data_in_frame_22_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i227_LC_20_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i227_LC_20_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i227_LC_20_25_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i227_LC_20_25_5  (
            .in0(N__79861),
            .in1(N__80719),
            .in2(N__74000),
            .in3(N__73930),
            .lcout(\c0.data_in_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i222_LC_20_25_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i222_LC_20_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i222_LC_20_25_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i222_LC_20_25_6  (
            .in0(N__78139),
            .in1(N__75011),
            .in2(N__73980),
            .in3(N__79864),
            .lcout(\c0.data_in_frame_27_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i225_LC_20_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i225_LC_20_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i225_LC_20_25_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i225_LC_20_25_7  (
            .in0(N__79860),
            .in1(N__73688),
            .in2(N__73948),
            .in3(N__80877),
            .lcout(\c0.data_in_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97747),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1531_LC_20_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1531_LC_20_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1531_LC_20_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1531_LC_20_26_0  (
            .in0(N__74290),
            .in1(N__74354),
            .in2(_gnd_net_),
            .in3(N__79469),
            .lcout(\c0.n17627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i199_LC_20_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i199_LC_20_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i199_LC_20_26_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i199_LC_20_26_1  (
            .in0(N__81026),
            .in1(N__73672),
            .in2(N__79878),
            .in3(N__79422),
            .lcout(\c0.data_in_frame_24_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1656_LC_20_26_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1656_LC_20_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1656_LC_20_26_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1656_LC_20_26_2  (
            .in0(N__79421),
            .in1(N__73404),
            .in2(_gnd_net_),
            .in3(N__74807),
            .lcout(\c0.n33933 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i218_LC_20_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i218_LC_20_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i218_LC_20_26_3 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0__i218_LC_20_26_3  (
            .in0(N__75362),
            .in1(N__73352),
            .in2(N__78289),
            .in3(N__79871),
            .lcout(\c0.data_in_frame_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i171_LC_20_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i171_LC_20_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i171_LC_20_26_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i171_LC_20_26_5  (
            .in0(N__78422),
            .in1(N__80700),
            .in2(N__73292),
            .in3(N__78504),
            .lcout(\c0.data_in_frame_21_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i170_LC_20_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i170_LC_20_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i170_LC_20_26_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i170_LC_20_26_6  (
            .in0(N__78503),
            .in1(N__78423),
            .in2(N__73326),
            .in3(N__75363),
            .lcout(\c0.data_in_frame_21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1681_LC_20_26_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1681_LC_20_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1681_LC_20_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1681_LC_20_26_7  (
            .in0(N__73312),
            .in1(N__79002),
            .in2(N__73291),
            .in3(N__74565),
            .lcout(\c0.n33467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i220_LC_20_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i220_LC_20_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i220_LC_20_27_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i220_LC_20_27_0  (
            .in0(N__78240),
            .in1(N__78988),
            .in2(N__74523),
            .in3(N__79845),
            .lcout(\c0.data_in_frame_27_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1655_LC_20_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1655_LC_20_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1655_LC_20_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1655_LC_20_27_2  (
            .in0(_gnd_net_),
            .in1(N__74174),
            .in2(_gnd_net_),
            .in3(N__75110),
            .lcout(\c0.n33678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i238_LC_20_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i238_LC_20_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i238_LC_20_27_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i238_LC_20_27_3  (
            .in0(N__74453),
            .in1(N__75085),
            .in2(N__74475),
            .in3(N__78516),
            .lcout(\c0.data_in_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i236_LC_20_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i236_LC_20_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i236_LC_20_27_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i236_LC_20_27_4  (
            .in0(N__78515),
            .in1(N__78989),
            .in2(N__74370),
            .in3(N__74454),
            .lcout(\c0.data_in_frame_29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97778),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1573_LC_20_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1573_LC_20_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1573_LC_20_27_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1573_LC_20_27_5  (
            .in0(N__79485),
            .in1(N__74355),
            .in2(N__74291),
            .in3(N__74226),
            .lcout(\c0.n33762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1660_LC_20_27_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1660_LC_20_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1660_LC_20_27_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_1660_LC_20_27_7  (
            .in0(N__74175),
            .in1(N__74673),
            .in2(_gnd_net_),
            .in3(N__79395),
            .lcout(\c0.n32259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1648_LC_20_28_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1648_LC_20_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1648_LC_20_28_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1648_LC_20_28_0  (
            .in0(N__74127),
            .in1(N__74092),
            .in2(N__75393),
            .in3(N__74061),
            .lcout(\c0.n33988 ),
            .ltout(\c0.n33988_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1646_LC_20_28_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1646_LC_20_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1646_LC_20_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1646_LC_20_28_1  (
            .in0(_gnd_net_),
            .in1(N__74042),
            .in2(N__74025),
            .in3(N__75106),
            .lcout(\c0.n33536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i200_LC_20_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i200_LC_20_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i200_LC_20_28_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0__i200_LC_20_28_3  (
            .in0(N__80135),
            .in1(N__81104),
            .in2(N__79879),
            .in3(N__75391),
            .lcout(\c0.data_in_frame_24_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i202_LC_20_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i202_LC_20_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i202_LC_20_28_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i202_LC_20_28_4  (
            .in0(N__79854),
            .in1(N__75372),
            .in2(N__75111),
            .in3(N__87263),
            .lcout(\c0.data_in_frame_25_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i198_LC_20_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i198_LC_20_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i198_LC_20_28_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i198_LC_20_28_5  (
            .in0(N__75010),
            .in1(N__81103),
            .in2(N__74759),
            .in3(N__79855),
            .lcout(\c0.data_in_frame_24_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97790),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1665_LC_20_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1665_LC_20_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1665_LC_20_28_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_1665_LC_20_28_6  (
            .in0(N__74808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74752),
            .lcout(),
            .ltout(\c0.n33930_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1659_LC_20_28_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1659_LC_20_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1659_LC_20_28_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1659_LC_20_28_7  (
            .in0(N__79623),
            .in1(N__74736),
            .in2(N__74730),
            .in3(N__74726),
            .lcout(\c0.n10_adj_4674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i7_4_lut_adj_1284_LC_21_4_1 .C_ON=1'b0;
    defparam \quad_counter1.i7_4_lut_adj_1284_LC_21_4_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i7_4_lut_adj_1284_LC_21_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i7_4_lut_adj_1284_LC_21_4_1  (
            .in0(N__74659),
            .in1(N__74638),
            .in2(N__74623),
            .in3(N__74590),
            .lcout(\quad_counter1.n18_adj_4457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23553_2_lut_LC_21_4_3 .C_ON=1'b0;
    defparam \quad_counter1.i23553_2_lut_LC_21_4_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23553_2_lut_LC_21_4_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter1.i23553_2_lut_LC_21_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__75528),
            .in3(N__81796),
            .lcout(),
            .ltout(\quad_counter1.n28269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1302_LC_21_4_4 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1302_LC_21_4_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1302_LC_21_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1302_LC_21_4_4  (
            .in0(N__75499),
            .in1(N__75415),
            .in2(N__74568),
            .in3(N__75478),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4468_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1304_LC_21_4_5 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1304_LC_21_4_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1304_LC_21_4_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1304_LC_21_4_5  (
            .in0(N__75436),
            .in1(N__75613),
            .in2(N__75573),
            .in3(N__75457),
            .lcout(\quad_counter1.n14_adj_4470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30703_1_lut_LC_21_4_7 .C_ON=1'b0;
    defparam \quad_counter1.i30703_1_lut_LC_21_4_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30703_1_lut_LC_21_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter1.i30703_1_lut_LC_21_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81567),
            .lcout(\quad_counter1.n36130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_2_lut_LC_21_5_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_2_lut_LC_21_5_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_2_lut_LC_21_5_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1817_2_lut_LC_21_5_0  (
            .in0(N__86955),
            .in1(N__86954),
            .in2(N__81340),
            .in3(N__75507),
            .lcout(\quad_counter1.n2719 ),
            .ltout(),
            .carryin(bfn_21_5_0_),
            .carryout(\quad_counter1.n30535 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_3_lut_LC_21_5_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_3_lut_LC_21_5_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_3_lut_LC_21_5_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_3_lut_LC_21_5_1  (
            .in0(N__86883),
            .in1(N__86882),
            .in2(N__81403),
            .in3(N__75483),
            .lcout(\quad_counter1.n2718 ),
            .ltout(),
            .carryin(\quad_counter1.n30535 ),
            .carryout(\quad_counter1.n30536 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_4_lut_LC_21_5_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_4_lut_LC_21_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_4_lut_LC_21_5_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1817_4_lut_LC_21_5_2  (
            .in0(N__86826),
            .in1(N__86825),
            .in2(N__81341),
            .in3(N__75462),
            .lcout(\quad_counter1.n2717 ),
            .ltout(),
            .carryin(\quad_counter1.n30536 ),
            .carryout(\quad_counter1.n30537 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_5_lut_LC_21_5_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_5_lut_LC_21_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_5_lut_LC_21_5_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1817_5_lut_LC_21_5_3  (
            .in0(N__86775),
            .in1(N__86774),
            .in2(N__81344),
            .in3(N__75441),
            .lcout(\quad_counter1.n2716 ),
            .ltout(),
            .carryin(\quad_counter1.n30537 ),
            .carryout(\quad_counter1.n30538 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_6_lut_LC_21_5_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_6_lut_LC_21_5_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_6_lut_LC_21_5_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1817_6_lut_LC_21_5_4  (
            .in0(N__86724),
            .in1(N__86723),
            .in2(N__81342),
            .in3(N__75420),
            .lcout(\quad_counter1.n2715 ),
            .ltout(),
            .carryin(\quad_counter1.n30538 ),
            .carryout(\quad_counter1.n30539 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_7_lut_LC_21_5_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_7_lut_LC_21_5_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_7_lut_LC_21_5_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1817_7_lut_LC_21_5_5  (
            .in0(N__86673),
            .in1(N__86672),
            .in2(N__81345),
            .in3(N__75399),
            .lcout(\quad_counter1.n2714 ),
            .ltout(),
            .carryin(\quad_counter1.n30539 ),
            .carryout(\quad_counter1.n30540 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_8_lut_LC_21_5_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_8_lut_LC_21_5_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_8_lut_LC_21_5_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1817_8_lut_LC_21_5_6  (
            .in0(N__87693),
            .in1(N__87692),
            .in2(N__81343),
            .in3(N__75396),
            .lcout(\quad_counter1.n2713 ),
            .ltout(),
            .carryin(\quad_counter1.n30540 ),
            .carryout(\quad_counter1.n30541 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_9_lut_LC_21_5_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_9_lut_LC_21_5_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_9_lut_LC_21_5_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_9_lut_LC_21_5_7  (
            .in0(N__87642),
            .in1(N__87641),
            .in2(N__81404),
            .in3(N__75597),
            .lcout(\quad_counter1.n2712 ),
            .ltout(),
            .carryin(\quad_counter1.n30541 ),
            .carryout(\quad_counter1.n30542 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_10_lut_LC_21_6_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_10_lut_LC_21_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_10_lut_LC_21_6_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_10_lut_LC_21_6_0  (
            .in0(N__87591),
            .in1(N__87590),
            .in2(N__81405),
            .in3(N__75594),
            .lcout(\quad_counter1.n2711 ),
            .ltout(),
            .carryin(bfn_21_6_0_),
            .carryout(\quad_counter1.n30543 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_11_lut_LC_21_6_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_11_lut_LC_21_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_11_lut_LC_21_6_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_11_lut_LC_21_6_1  (
            .in0(N__87540),
            .in1(N__87539),
            .in2(N__81409),
            .in3(N__75591),
            .lcout(\quad_counter1.n2710 ),
            .ltout(),
            .carryin(\quad_counter1.n30543 ),
            .carryout(\quad_counter1.n30544 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_12_lut_LC_21_6_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_12_lut_LC_21_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_12_lut_LC_21_6_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_12_lut_LC_21_6_2  (
            .in0(N__87480),
            .in1(N__87479),
            .in2(N__81406),
            .in3(N__75588),
            .lcout(\quad_counter1.n2709 ),
            .ltout(),
            .carryin(\quad_counter1.n30544 ),
            .carryout(\quad_counter1.n30545 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_13_lut_LC_21_6_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_13_lut_LC_21_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_13_lut_LC_21_6_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_13_lut_LC_21_6_3  (
            .in0(N__87423),
            .in1(N__87422),
            .in2(N__81410),
            .in3(N__75585),
            .lcout(\quad_counter1.n2708 ),
            .ltout(),
            .carryin(\quad_counter1.n30545 ),
            .carryout(\quad_counter1.n30546 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_14_lut_LC_21_6_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_14_lut_LC_21_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_14_lut_LC_21_6_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_14_lut_LC_21_6_4  (
            .in0(N__87363),
            .in1(N__87362),
            .in2(N__81407),
            .in3(N__75582),
            .lcout(\quad_counter1.n2707 ),
            .ltout(),
            .carryin(\quad_counter1.n30546 ),
            .carryout(\quad_counter1.n30547 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_15_lut_LC_21_6_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1817_15_lut_LC_21_6_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_15_lut_LC_21_6_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_15_lut_LC_21_6_5  (
            .in0(N__88035),
            .in1(N__88034),
            .in2(N__81411),
            .in3(N__75579),
            .lcout(\quad_counter1.n2706 ),
            .ltout(),
            .carryin(\quad_counter1.n30547 ),
            .carryout(\quad_counter1.n30548 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1817_16_lut_LC_21_6_6 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1817_16_lut_LC_21_6_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1817_16_lut_LC_21_6_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1817_16_lut_LC_21_6_6  (
            .in0(N__87974),
            .in1(N__87975),
            .in2(N__81408),
            .in3(N__75576),
            .lcout(\quad_counter1.n2705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i6_4_lut_adj_1278_LC_21_8_0 .C_ON=1'b0;
    defparam \quad_counter1.i6_4_lut_adj_1278_LC_21_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i6_4_lut_adj_1278_LC_21_8_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i6_4_lut_adj_1278_LC_21_8_0  (
            .in0(N__87551),
            .in1(N__87385),
            .in2(N__87508),
            .in3(N__87602),
            .lcout(),
            .ltout(\quad_counter1.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i7_4_lut_LC_21_8_1 .C_ON=1'b0;
    defparam \quad_counter1.i7_4_lut_LC_21_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i7_4_lut_LC_21_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i7_4_lut_LC_21_8_1  (
            .in0(N__87325),
            .in1(N__75633),
            .in2(N__75642),
            .in3(N__87997),
            .lcout(\quad_counter1.n2540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23557_2_lut_LC_21_8_2 .C_ON=1'b0;
    defparam \quad_counter1.i23557_2_lut_LC_21_8_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23557_2_lut_LC_21_8_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \quad_counter1.i23557_2_lut_LC_21_8_2  (
            .in0(N__86899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86837),
            .lcout(),
            .ltout(\quad_counter1.n28273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1277_LC_21_8_3 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1277_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1277_LC_21_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1277_LC_21_8_3  (
            .in0(N__86735),
            .in1(N__87653),
            .in2(N__75639),
            .in3(N__86786),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_4_lut_adj_1279_LC_21_8_4 .C_ON=1'b0;
    defparam \quad_counter1.i1_4_lut_adj_1279_LC_21_8_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_4_lut_adj_1279_LC_21_8_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i1_4_lut_adj_1279_LC_21_8_4  (
            .in0(N__86684),
            .in1(N__87442),
            .in2(N__75636),
            .in3(N__87704),
            .lcout(\quad_counter1.n9_adj_4451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_5_i3_2_lut_LC_21_8_5 .C_ON=1'b0;
    defparam \c0.select_369_Select_5_i3_2_lut_LC_21_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_5_i3_2_lut_LC_21_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_5_i3_2_lut_LC_21_8_5  (
            .in0(N__91519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94800),
            .lcout(\c0.n3_adj_4584 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_2_lut_LC_21_9_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_2_lut_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_2_lut_LC_21_9_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1683_2_lut_LC_21_9_0  (
            .in0(N__88124),
            .in1(N__88123),
            .in2(N__75790),
            .in3(N__75627),
            .lcout(\quad_counter1.n2519 ),
            .ltout(),
            .carryin(bfn_21_9_0_),
            .carryout(\quad_counter1.n30510 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_3_lut_LC_21_9_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_3_lut_LC_21_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_3_lut_LC_21_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_3_lut_LC_21_9_1  (
            .in0(N__88074),
            .in1(N__88073),
            .in2(N__75746),
            .in3(N__75624),
            .lcout(\quad_counter1.n2518 ),
            .ltout(),
            .carryin(\quad_counter1.n30510 ),
            .carryout(\quad_counter1.n30511 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_4_lut_LC_21_9_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_4_lut_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_4_lut_LC_21_9_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1683_4_lut_LC_21_9_2  (
            .in0(N__88101),
            .in1(N__88100),
            .in2(N__75791),
            .in3(N__75621),
            .lcout(\quad_counter1.n2517 ),
            .ltout(),
            .carryin(\quad_counter1.n30511 ),
            .carryout(\quad_counter1.n30512 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_5_lut_LC_21_9_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_5_lut_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_5_lut_LC_21_9_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1683_5_lut_LC_21_9_3  (
            .in0(N__87833),
            .in1(N__87832),
            .in2(N__75794),
            .in3(N__75618),
            .lcout(\quad_counter1.n2516 ),
            .ltout(),
            .carryin(\quad_counter1.n30512 ),
            .carryout(\quad_counter1.n30513 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_6_lut_LC_21_9_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_6_lut_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_6_lut_LC_21_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1683_6_lut_LC_21_9_4  (
            .in0(N__87806),
            .in1(N__87805),
            .in2(N__75792),
            .in3(N__75669),
            .lcout(\quad_counter1.n2515 ),
            .ltout(),
            .carryin(\quad_counter1.n30513 ),
            .carryout(\quad_counter1.n30514 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_7_lut_LC_21_9_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_7_lut_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_7_lut_LC_21_9_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1683_7_lut_LC_21_9_5  (
            .in0(N__87776),
            .in1(N__87775),
            .in2(N__75795),
            .in3(N__75666),
            .lcout(\quad_counter1.n2514 ),
            .ltout(),
            .carryin(\quad_counter1.n30514 ),
            .carryout(\quad_counter1.n30515 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_8_lut_LC_21_9_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_8_lut_LC_21_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_8_lut_LC_21_9_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1683_8_lut_LC_21_9_6  (
            .in0(N__87746),
            .in1(N__87745),
            .in2(N__75793),
            .in3(N__75663),
            .lcout(\quad_counter1.n2513 ),
            .ltout(),
            .carryin(\quad_counter1.n30515 ),
            .carryout(\quad_counter1.n30516 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_9_lut_LC_21_9_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_9_lut_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_9_lut_LC_21_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_9_lut_LC_21_9_7  (
            .in0(N__88308),
            .in1(N__88307),
            .in2(N__75747),
            .in3(N__75660),
            .lcout(\quad_counter1.n2512 ),
            .ltout(),
            .carryin(\quad_counter1.n30516 ),
            .carryout(\quad_counter1.n30517 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_10_lut_LC_21_10_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_10_lut_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_10_lut_LC_21_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_10_lut_LC_21_10_0  (
            .in0(N__88275),
            .in1(N__88274),
            .in2(N__75735),
            .in3(N__75657),
            .lcout(\quad_counter1.n2511 ),
            .ltout(),
            .carryin(bfn_21_10_0_),
            .carryout(\quad_counter1.n30518 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_11_lut_LC_21_10_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_11_lut_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_11_lut_LC_21_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_11_lut_LC_21_10_1  (
            .in0(N__88240),
            .in1(N__88241),
            .in2(N__75744),
            .in3(N__75654),
            .lcout(\quad_counter1.n2510 ),
            .ltout(),
            .carryin(\quad_counter1.n30518 ),
            .carryout(\quad_counter1.n30519 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_12_lut_LC_21_10_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_12_lut_LC_21_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_12_lut_LC_21_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_12_lut_LC_21_10_2  (
            .in0(N__88207),
            .in1(N__88208),
            .in2(N__75736),
            .in3(N__75651),
            .lcout(\quad_counter1.n2509 ),
            .ltout(),
            .carryin(\quad_counter1.n30519 ),
            .carryout(\quad_counter1.n30520 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_13_lut_LC_21_10_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1683_13_lut_LC_21_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_13_lut_LC_21_10_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_13_lut_LC_21_10_3  (
            .in0(N__88178),
            .in1(N__88177),
            .in2(N__75745),
            .in3(N__75648),
            .lcout(\quad_counter1.n2508 ),
            .ltout(),
            .carryin(\quad_counter1.n30520 ),
            .carryout(\quad_counter1.n30521 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1683_14_lut_LC_21_10_4 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1683_14_lut_LC_21_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1683_14_lut_LC_21_10_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1683_14_lut_LC_21_10_4  (
            .in0(N__88147),
            .in1(N__88148),
            .in2(N__75737),
            .in3(N__75645),
            .lcout(\quad_counter1.n2507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30707_1_lut_LC_21_10_7 .C_ON=1'b0;
    defparam \quad_counter1.i30707_1_lut_LC_21_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30707_1_lut_LC_21_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter1.i30707_1_lut_LC_21_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75714),
            .lcout(\quad_counter1.n36134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i6_4_lut_LC_21_11_1 .C_ON=1'b0;
    defparam \quad_counter1.i6_4_lut_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i6_4_lut_LC_21_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i6_4_lut_LC_21_11_1  (
            .in0(N__88273),
            .in1(N__88306),
            .in2(N__88212),
            .in3(N__75753),
            .lcout(\quad_counter1.n2441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_prev__i1_LC_21_11_3 .C_ON=1'b0;
    defparam \quad_counter1.count_prev__i1_LC_21_11_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_prev__i1_LC_21_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \quad_counter1.count_prev__i1_LC_21_11_3  (
            .in0(N__75683),
            .in1(N__101335),
            .in2(_gnd_net_),
            .in3(N__75690),
            .lcout(count_prev_0_adj_4815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97573),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i6_4_lut_adj_1301_LC_21_11_4 .C_ON=1'b0;
    defparam \quad_counter1.i6_4_lut_adj_1301_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i6_4_lut_adj_1301_LC_21_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i6_4_lut_adj_1301_LC_21_11_4  (
            .in0(N__81756),
            .in1(N__81705),
            .in2(N__81732),
            .in3(N__82425),
            .lcout(n34871),
            .ltout(n34871_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_per_millisecond_i0_i0_LC_21_11_5 .C_ON=1'b0;
    defparam \quad_counter1.count_per_millisecond_i0_i0_LC_21_11_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_per_millisecond_i0_i0_LC_21_11_5 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \quad_counter1.count_per_millisecond_i0_i0_LC_21_11_5  (
            .in0(N__75684),
            .in1(N__97843),
            .in2(N__75675),
            .in3(N__101336),
            .lcout(data_out_frame_29__7__N_1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97573),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_21__0__5357_LC_21_11_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_21__0__5357_LC_21_11_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_21__0__5357_LC_21_11_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.data_out_frame_21__0__5357_LC_21_11_6  (
            .in0(N__97844),
            .in1(N__85277),
            .in2(N__89867),
            .in3(N__84678),
            .lcout(data_out_frame_21_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97573),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_3_lut_adj_1246_LC_21_13_1 .C_ON=1'b0;
    defparam \quad_counter1.i1_3_lut_adj_1246_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_3_lut_adj_1246_LC_21_13_1 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \quad_counter1.i1_3_lut_adj_1246_LC_21_13_1  (
            .in0(_gnd_net_),
            .in1(N__88390),
            .in2(N__88353),
            .in3(N__88327),
            .lcout(\quad_counter1.n7_adj_4425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_2_lut_adj_1244_LC_21_13_2 .C_ON=1'b0;
    defparam \quad_counter1.i1_2_lut_adj_1244_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_2_lut_adj_1244_LC_21_13_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter1.i1_2_lut_adj_1244_LC_21_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__88875),
            .in3(N__88567),
            .lcout(),
            .ltout(\quad_counter1.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i13_4_lut_LC_21_13_3 .C_ON=1'b0;
    defparam \quad_counter1.i13_4_lut_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i13_4_lut_LC_21_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i13_4_lut_LC_21_13_3  (
            .in0(N__88906),
            .in1(N__88776),
            .in2(N__75672),
            .in3(N__88837),
            .lcout(\quad_counter1.n30_adj_4426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_adj_1245_LC_21_13_4 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_adj_1245_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_adj_1245_LC_21_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \quad_counter1.i2_2_lut_adj_1245_LC_21_13_4  (
            .in0(_gnd_net_),
            .in1(N__88648),
            .in2(_gnd_net_),
            .in3(N__88714),
            .lcout(),
            .ltout(\quad_counter1.n8_adj_4424_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1247_LC_21_13_5 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1247_LC_21_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1247_LC_21_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1247_LC_21_13_5  (
            .in0(N__88669),
            .in1(N__76014),
            .in2(N__76008),
            .in3(N__88687),
            .lcout(\quad_counter1.n35050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_LC_21_14_6 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_LC_21_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_LC_21_14_6  (
            .in0(N__76005),
            .in1(N__75999),
            .in2(N__75993),
            .in3(N__75984),
            .lcout(\quad_counter1.n3332 ),
            .ltout(\quad_counter1.n3332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30719_1_lut_LC_21_14_7 .C_ON=1'b0;
    defparam \quad_counter1.i30719_1_lut_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30719_1_lut_LC_21_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30719_1_lut_LC_21_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__75978),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__2__5419_LC_21_15_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__2__5419_LC_21_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__2__5419_LC_21_15_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_13__2__5419_LC_21_15_3  (
            .in0(N__85284),
            .in1(N__89198),
            .in2(N__86599),
            .in3(N__84454),
            .lcout(data_out_frame_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97609),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i4_LC_21_16_0 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i4_LC_21_16_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i4_LC_21_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.count_i0_i4_LC_21_16_0  (
            .in0(N__85817),
            .in1(N__75975),
            .in2(_gnd_net_),
            .in3(N__76545),
            .lcout(encoder1_position_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97621),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i2_LC_21_16_1 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i2_LC_21_16_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i2_LC_21_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i2_LC_21_16_1  (
            .in0(N__76544),
            .in1(N__75966),
            .in2(_gnd_net_),
            .in3(N__86583),
            .lcout(encoder1_position_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97621),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_21_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_21_16_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_21_16_2  (
            .in0(N__95601),
            .in1(N__83342),
            .in2(_gnd_net_),
            .in3(N__96145),
            .lcout(\c0.n26_adj_4516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1615_LC_21_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1615_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1615_LC_21_16_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i1_2_lut_adj_1615_LC_21_16_5  (
            .in0(_gnd_net_),
            .in1(N__90096),
            .in2(_gnd_net_),
            .in3(N__90343),
            .lcout(\c0.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_21_17_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_21_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_21_17_2  (
            .in0(N__76677),
            .in1(N__75943),
            .in2(N__75874),
            .in3(N__75837),
            .lcout(),
            .ltout(\c0.n12_adj_4553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1427_LC_21_17_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1427_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1427_LC_21_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1427_LC_21_17_3  (
            .in0(N__83059),
            .in1(N__76221),
            .in2(N__76197),
            .in3(N__77692),
            .lcout(\c0.n15711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_17__0__5389_LC_21_17_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_17__0__5389_LC_21_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_17__0__5389_LC_21_17_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.data_out_frame_17__0__5389_LC_21_17_4  (
            .in0(N__84694),
            .in1(N__85282),
            .in2(N__100780),
            .in3(N__89840),
            .lcout(data_out_frame_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__3__5418_LC_21_17_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__3__5418_LC_21_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__3__5418_LC_21_17_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_13__3__5418_LC_21_17_5  (
            .in0(N__85281),
            .in1(N__76190),
            .in2(N__83541),
            .in3(N__84696),
            .lcout(data_out_frame_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__6__5287_LC_21_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__6__5287_LC_21_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__6__5287_LC_21_17_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \c0.data_out_frame_29__6__5287_LC_21_17_6  (
            .in0(N__84695),
            .in1(N__76175),
            .in2(N__95652),
            .in3(N__85283),
            .lcout(data_out_frame_29_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97635),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i12_LC_21_17_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i12_LC_21_17_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i12_LC_21_17_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter1.count_i0_i12_LC_21_17_7  (
            .in0(N__76589),
            .in1(N__76161),
            .in2(_gnd_net_),
            .in3(N__76050),
            .lcout(encoder1_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1387_LC_21_18_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1387_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1387_LC_21_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1387_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__76100),
            .in2(N__77394),
            .in3(N__77312),
            .lcout(\c0.n31280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i0_LC_21_18_2 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i0_LC_21_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i0_LC_21_18_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i0_LC_21_18_2  (
            .in0(N__83178),
            .in1(N__76152),
            .in2(_gnd_net_),
            .in3(N__77631),
            .lcout(control_mode_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97649),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1760_LC_21_18_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1760_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1760_LC_21_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1760_LC_21_18_3  (
            .in0(N__77903),
            .in1(N__77286),
            .in2(N__76101),
            .in3(N__77390),
            .lcout(\c0.n32304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1408_LC_21_18_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1408_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1408_LC_21_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1408_LC_21_18_4  (
            .in0(N__77389),
            .in1(N__76043),
            .in2(_gnd_net_),
            .in3(N__76266),
            .lcout(\c0.n18232 ),
            .ltout(\c0.n18232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1719_LC_21_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1719_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1719_LC_21_18_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1719_LC_21_18_5  (
            .in0(_gnd_net_),
            .in1(N__83482),
            .in2(N__76605),
            .in3(N__83423),
            .lcout(\c0.n32275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1433_LC_21_18_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1433_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1433_LC_21_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1433_LC_21_18_6  (
            .in0(N__77287),
            .in1(N__77313),
            .in2(N__98158),
            .in3(N__77904),
            .lcout(\c0.n17515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.count_i0_i6_LC_21_18_7 .C_ON=1'b0;
    defparam \quad_counter1.count_i0_i6_LC_21_18_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.count_i0_i6_LC_21_18_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \quad_counter1.count_i0_i6_LC_21_18_7  (
            .in0(N__76602),
            .in1(N__76585),
            .in2(_gnd_net_),
            .in3(N__94295),
            .lcout(encoder1_position_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97649),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_5__I_0_2_lut_LC_21_19_1 .C_ON=1'b0;
    defparam \c0.control_mode_5__I_0_2_lut_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.control_mode_5__I_0_2_lut_LC_21_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.control_mode_5__I_0_2_lut_LC_21_19_1  (
            .in0(_gnd_net_),
            .in1(N__76808),
            .in2(_gnd_net_),
            .in3(N__77554),
            .lcout(\c0.data_out_frame_29__7__N_740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1481_LC_21_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1481_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1481_LC_21_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1481_LC_21_19_3  (
            .in0(_gnd_net_),
            .in1(N__86638),
            .in2(_gnd_net_),
            .in3(N__85542),
            .lcout(),
            .ltout(\c0.data_out_frame_29__7__N_976_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_21_19_4 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_21_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_LC_21_19_4  (
            .in0(N__76356),
            .in1(N__77500),
            .in2(N__76338),
            .in3(N__76335),
            .lcout(\c0.n42_adj_4570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1450_LC_21_19_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1450_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1450_LC_21_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1450_LC_21_19_5  (
            .in0(N__76308),
            .in1(N__76290),
            .in2(N__76284),
            .in3(N__76272),
            .lcout(\c0.n35113 ),
            .ltout(\c0.n35113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1452_LC_21_19_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1452_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1452_LC_21_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i5_4_lut_adj_1452_LC_21_19_6  (
            .in0(N__76262),
            .in1(N__77902),
            .in2(N__76239),
            .in3(N__76236),
            .lcout(),
            .ltout(\c0.n12_adj_4561_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1453_LC_21_19_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1453_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1453_LC_21_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1453_LC_21_19_7  (
            .in0(N__83081),
            .in1(N__97976),
            .in2(N__76224),
            .in3(N__83422),
            .lcout(\c0.n17684 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_21_20_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_21_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_21_20_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_21_20_0  (
            .in0(N__77103),
            .in1(N__77058),
            .in2(_gnd_net_),
            .in3(N__77031),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97679),
            .ce(),
            .sr(N__76932));
    defparam \c0.encoder0_position_31__I_0_2_lut_LC_21_20_1 .C_ON=1'b0;
    defparam \c0.encoder0_position_31__I_0_2_lut_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.encoder0_position_31__I_0_2_lut_LC_21_20_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.encoder0_position_31__I_0_2_lut_LC_21_20_1  (
            .in0(N__76856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76906),
            .lcout(\c0.data_out_frame_29__7__N_756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1475_LC_21_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1475_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1475_LC_21_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1475_LC_21_20_2  (
            .in0(_gnd_net_),
            .in1(N__76855),
            .in2(_gnd_net_),
            .in3(N__79064),
            .lcout(\c0.n33732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_2_lut_LC_21_20_3 .C_ON=1'b0;
    defparam \c0.i13_2_lut_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_2_lut_LC_21_20_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i13_2_lut_LC_21_20_3  (
            .in0(_gnd_net_),
            .in1(N__92397),
            .in2(_gnd_net_),
            .in3(N__91746),
            .lcout(\c0.n39_adj_4644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_1_i3_2_lut_LC_21_20_6 .C_ON=1'b0;
    defparam \c0.select_369_Select_1_i3_2_lut_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_1_i3_2_lut_LC_21_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_1_i3_2_lut_LC_21_20_6  (
            .in0(_gnd_net_),
            .in1(N__91115),
            .in2(_gnd_net_),
            .in3(N__94750),
            .lcout(\c0.n3_adj_4579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1753_LC_21_21_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1753_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1753_LC_21_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1753_LC_21_21_0  (
            .in0(N__77711),
            .in1(N__76790),
            .in2(N__76751),
            .in3(N__77542),
            .lcout(\c0.n18199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_89_i9_2_lut_3_lut_LC_21_21_1 .C_ON=1'b0;
    defparam \c0.equal_89_i9_2_lut_3_lut_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.equal_89_i9_2_lut_3_lut_LC_21_21_1 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \c0.equal_89_i9_2_lut_3_lut_LC_21_21_1  (
            .in0(_gnd_net_),
            .in1(N__91251),
            .in2(N__91116),
            .in3(N__93227),
            .lcout(\c0.n9_adj_4530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1459_LC_21_21_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1459_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1459_LC_21_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1459_LC_21_21_3  (
            .in0(N__76652),
            .in1(N__86411),
            .in2(N__76614),
            .in3(N__83309),
            .lcout(\c0.n33425 ),
            .ltout(\c0.n33425_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1457_LC_21_21_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1457_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1457_LC_21_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1457_LC_21_21_4  (
            .in0(N__77712),
            .in1(N__85459),
            .in2(N__77703),
            .in3(N__77691),
            .lcout(\c0.n18901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.control_mode_i0_i4_LC_21_21_5 .C_ON=1'b0;
    defparam \c0.control_mode_i0_i4_LC_21_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.control_mode_i0_i4_LC_21_21_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.control_mode_i0_i4_LC_21_21_5  (
            .in0(N__77543),
            .in1(N__83594),
            .in2(_gnd_net_),
            .in3(N__77626),
            .lcout(control_mode_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97696),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1414_LC_21_21_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1414_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1414_LC_21_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1414_LC_21_21_6  (
            .in0(N__77508),
            .in1(N__77435),
            .in2(N__77373),
            .in3(N__77408),
            .lcout(\c0.n33393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1400_LC_21_22_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1400_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1400_LC_21_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1400_LC_21_22_1  (
            .in0(N__77366),
            .in1(N__77351),
            .in2(_gnd_net_),
            .in3(N__77733),
            .lcout(\c0.n33496 ),
            .ltout(\c0.n33496_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1706_LC_21_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1706_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1706_LC_21_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1706_LC_21_22_2  (
            .in0(_gnd_net_),
            .in1(N__79226),
            .in2(N__77298),
            .in3(N__85921),
            .lcout(),
            .ltout(\c0.n6_adj_4544_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1402_LC_21_22_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1402_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1402_LC_21_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1402_LC_21_22_3  (
            .in0(N__77760),
            .in1(N__77294),
            .in2(N__77241),
            .in3(N__86226),
            .lcout(\c0.n17536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i30672_3_lut_LC_21_22_4.C_ON=1'b0;
    defparam i30672_3_lut_LC_21_22_4.SEQ_MODE=4'b0000;
    defparam i30672_3_lut_LC_21_22_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i30672_3_lut_LC_21_22_4 (
            .in0(N__77238),
            .in1(N__77226),
            .in2(_gnd_net_),
            .in3(N__95791),
            .lcout(n36101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_21_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_21_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_21_22_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i16_LC_21_22_6  (
            .in0(N__87187),
            .in1(N__77185),
            .in2(N__83954),
            .in3(N__80119),
            .lcout(data_in_frame_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97712),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i11_LC_21_22_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i11_LC_21_22_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i11_LC_21_22_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i11_LC_21_22_7  (
            .in0(N__77128),
            .in1(N__77157),
            .in2(_gnd_net_),
            .in3(N__86140),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97712),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i5_LC_21_23_0 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i5_LC_21_23_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i5_LC_21_23_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter0.count_i0_i5_LC_21_23_0  (
            .in0(N__96601),
            .in1(N__77976),
            .in2(_gnd_net_),
            .in3(N__86138),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97730),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i12_LC_21_23_1 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i12_LC_21_23_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i12_LC_21_23_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i12_LC_21_23_1  (
            .in0(N__86137),
            .in1(N__77961),
            .in2(_gnd_net_),
            .in3(N__79233),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97730),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1484_LC_21_23_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1484_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1484_LC_21_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1484_LC_21_23_2  (
            .in0(N__77947),
            .in1(N__77718),
            .in2(_gnd_net_),
            .in3(N__77731),
            .lcout(\c0.n18214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1476_LC_21_23_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1476_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1476_LC_21_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_1476_LC_21_23_3  (
            .in0(N__86489),
            .in1(N__77866),
            .in2(_gnd_net_),
            .in3(N__77820),
            .lcout(\c0.n33896 ),
            .ltout(\c0.n33896_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1749_LC_21_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1749_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1749_LC_21_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1749_LC_21_23_4  (
            .in0(_gnd_net_),
            .in1(N__79148),
            .in2(N__77772),
            .in3(N__86182),
            .lcout(\c0.n6_adj_4565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1477_LC_21_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1477_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1477_LC_21_23_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_1477_LC_21_23_5  (
            .in0(N__86183),
            .in1(_gnd_net_),
            .in2(N__79155),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n33360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1393_LC_21_23_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1393_LC_21_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1393_LC_21_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1393_LC_21_23_6  (
            .in0(N__77769),
            .in1(N__77759),
            .in2(N__77736),
            .in3(N__77732),
            .lcout(\c0.n33681 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1707_LC_21_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1707_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1707_LC_21_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1707_LC_21_24_1  (
            .in0(N__79222),
            .in1(N__85896),
            .in2(_gnd_net_),
            .in3(N__79154),
            .lcout(\c0.n18740 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1747_LC_21_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1747_LC_21_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1747_LC_21_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1747_LC_21_24_3  (
            .in0(N__79221),
            .in1(N__79191),
            .in2(N__85901),
            .in3(N__79153),
            .lcout(),
            .ltout(\c0.n6_adj_4566_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1479_LC_21_24_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1479_LC_21_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1479_LC_21_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1479_LC_21_24_4  (
            .in0(N__86225),
            .in1(N__79080),
            .in2(N__79074),
            .in3(N__79071),
            .lcout(\c0.n31429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1764_LC_21_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1764_LC_21_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1764_LC_21_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1764_LC_21_25_0  (
            .in0(_gnd_net_),
            .in1(N__78706),
            .in2(_gnd_net_),
            .in3(N__78349),
            .lcout(\c0.n18572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i172_LC_21_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i172_LC_21_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i172_LC_21_25_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i172_LC_21_25_1  (
            .in0(N__78978),
            .in1(N__78425),
            .in2(N__78715),
            .in3(N__78536),
            .lcout(\c0.data_in_frame_21_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1748_LC_21_25_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1748_LC_21_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1748_LC_21_25_3 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1748_LC_21_25_3  (
            .in0(N__93226),
            .in1(N__91103),
            .in2(N__91258),
            .in3(N__78693),
            .lcout(\c0.n33224 ),
            .ltout(\c0.n33224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i173_LC_21_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i173_LC_21_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i173_LC_21_25_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i173_LC_21_25_4  (
            .in0(N__78424),
            .in1(N__84244),
            .in2(N__78360),
            .in3(N__78350),
            .lcout(\c0.data_in_frame_21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_91_i9_2_lut_3_lut_LC_21_25_5 .C_ON=1'b0;
    defparam \c0.equal_91_i9_2_lut_3_lut_LC_21_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.equal_91_i9_2_lut_3_lut_LC_21_25_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.equal_91_i9_2_lut_3_lut_LC_21_25_5  (
            .in0(N__93224),
            .in1(N__91246),
            .in2(_gnd_net_),
            .in3(N__91101),
            .lcout(\c0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_88_i9_2_lut_3_lut_LC_21_25_6 .C_ON=1'b0;
    defparam \c0.equal_88_i9_2_lut_3_lut_LC_21_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.equal_88_i9_2_lut_3_lut_LC_21_25_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.equal_88_i9_2_lut_3_lut_LC_21_25_6  (
            .in0(N__91102),
            .in1(N__91250),
            .in2(_gnd_net_),
            .in3(N__93225),
            .lcout(\c0.n9_adj_4628 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i24_LC_21_25_7 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i24_LC_21_25_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i24_LC_21_25_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i24_LC_21_25_7  (
            .in0(N__86139),
            .in1(N__78060),
            .in2(_gnd_net_),
            .in3(N__78020),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97765),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i193_LC_21_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i193_LC_21_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i193_LC_21_26_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i193_LC_21_26_1  (
            .in0(N__81025),
            .in1(N__80975),
            .in2(N__79577),
            .in3(N__79869),
            .lcout(\c0.data_in_frame_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i211_LC_21_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i211_LC_21_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i211_LC_21_26_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i211_LC_21_26_6  (
            .in0(N__79868),
            .in1(N__80267),
            .in2(N__79593),
            .in3(N__80701),
            .lcout(\c0.data_in_frame_26_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i216_LC_21_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i216_LC_21_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i216_LC_21_26_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i216_LC_21_26_7  (
            .in0(N__80266),
            .in1(N__80136),
            .in2(N__79628),
            .in3(N__79870),
            .lcout(\c0.data_in_frame_26_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97779),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1778_LC_21_27_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1778_LC_21_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1778_LC_21_27_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1778_LC_21_27_1  (
            .in0(N__79589),
            .in1(N__79563),
            .in2(_gnd_net_),
            .in3(N__79525),
            .lcout(\c0.n31545 ),
            .ltout(\c0.n31545_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1690_LC_21_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1690_LC_21_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1690_LC_21_27_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1690_LC_21_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__79488),
            .in3(N__79484),
            .lcout(),
            .ltout(\c0.n19_adj_4699_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1700_LC_21_27_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1700_LC_21_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1700_LC_21_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_1700_LC_21_27_3  (
            .in0(N__79420),
            .in1(N__79407),
            .in2(N__79398),
            .in3(N__79394),
            .lcout(\c0.n32_adj_4705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i6_4_lut_adj_1303_LC_22_5_1 .C_ON=1'b0;
    defparam \quad_counter1.i6_4_lut_adj_1303_LC_22_5_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i6_4_lut_adj_1303_LC_22_5_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i6_4_lut_adj_1303_LC_22_5_1  (
            .in0(N__79360),
            .in1(N__79342),
            .in2(N__79326),
            .in3(N__79303),
            .lcout(),
            .ltout(\quad_counter1.n16_adj_4469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i8_3_lut_LC_22_5_2 .C_ON=1'b0;
    defparam \quad_counter1.i8_3_lut_LC_22_5_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i8_3_lut_LC_22_5_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter1.i8_3_lut_LC_22_5_2  (
            .in0(_gnd_net_),
            .in1(N__79285),
            .in2(N__79269),
            .in3(N__79264),
            .lcout(),
            .ltout(\quad_counter1.n18_adj_4471_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i9_4_lut_adj_1305_LC_22_5_3 .C_ON=1'b0;
    defparam \quad_counter1.i9_4_lut_adj_1305_LC_22_5_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i9_4_lut_adj_1305_LC_22_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i9_4_lut_adj_1305_LC_22_5_3  (
            .in0(N__81676),
            .in1(N__81660),
            .in2(N__81654),
            .in3(N__81649),
            .lcout(\quad_counter1.n2738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23531_2_lut_LC_22_5_4 .C_ON=1'b0;
    defparam \quad_counter1.i23531_2_lut_LC_22_5_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23531_2_lut_LC_22_5_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \quad_counter1.i23531_2_lut_LC_22_5_4  (
            .in0(N__82000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81547),
            .lcout(),
            .ltout(\quad_counter1.n28243_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1318_LC_22_5_5 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1318_LC_22_5_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1318_LC_22_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1318_LC_22_5_5  (
            .in0(N__81520),
            .in1(N__81491),
            .in2(N__81462),
            .in3(N__81458),
            .lcout(\quad_counter1.n10_adj_4483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_2_lut_LC_22_6_0 .C_ON=1'b0;
    defparam \quad_counter1.i1_2_lut_LC_22_6_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_2_lut_LC_22_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i1_2_lut_LC_22_6_0  (
            .in0(_gnd_net_),
            .in1(N__87532),
            .in2(_gnd_net_),
            .in3(N__87578),
            .lcout(),
            .ltout(\quad_counter1.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i7_4_lut_adj_1280_LC_22_6_1 .C_ON=1'b0;
    defparam \quad_counter1.i7_4_lut_adj_1280_LC_22_6_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i7_4_lut_adj_1280_LC_22_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i7_4_lut_adj_1280_LC_22_6_1  (
            .in0(N__87415),
            .in1(N__87355),
            .in2(N__81417),
            .in3(N__87472),
            .lcout(),
            .ltout(\quad_counter1.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i8_4_lut_LC_22_6_2 .C_ON=1'b0;
    defparam \quad_counter1.i8_4_lut_LC_22_6_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i8_4_lut_LC_22_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i8_4_lut_LC_22_6_2  (
            .in0(N__88027),
            .in1(N__86919),
            .in2(N__81414),
            .in3(N__87629),
            .lcout(\quad_counter1.n2639 ),
            .ltout(\quad_counter1.n2639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30705_1_lut_LC_22_6_3 .C_ON=1'b0;
    defparam \quad_counter1.i30705_1_lut_LC_22_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30705_1_lut_LC_22_6_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30705_1_lut_LC_22_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__81348),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_11__3__5434_LC_22_6_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_11__3__5434_LC_22_6_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_11__3__5434_LC_22_6_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_11__3__5434_LC_22_6_7  (
            .in0(N__81293),
            .in1(N__85251),
            .in2(N__83232),
            .in3(N__84558),
            .lcout(data_out_frame_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97550),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i0_LC_22_7_0 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i0_LC_22_7_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i0_LC_22_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i0_LC_22_7_0  (
            .in0(_gnd_net_),
            .in1(N__82091),
            .in2(_gnd_net_),
            .in3(N__81762),
            .lcout(\quad_counter1.millisecond_counter_0 ),
            .ltout(),
            .carryin(bfn_22_7_0_),
            .carryout(\quad_counter1.n30171 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i1_LC_22_7_1 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i1_LC_22_7_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i1_LC_22_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i1_LC_22_7_1  (
            .in0(_gnd_net_),
            .in1(N__82472),
            .in2(_gnd_net_),
            .in3(N__81759),
            .lcout(\quad_counter1.millisecond_counter_1 ),
            .ltout(),
            .carryin(\quad_counter1.n30171 ),
            .carryout(\quad_counter1.n30172 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i2_LC_22_7_2 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i2_LC_22_7_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i2_LC_22_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i2_LC_22_7_2  (
            .in0(_gnd_net_),
            .in1(N__81749),
            .in2(_gnd_net_),
            .in3(N__81738),
            .lcout(\quad_counter1.millisecond_counter_2 ),
            .ltout(),
            .carryin(\quad_counter1.n30172 ),
            .carryout(\quad_counter1.n30173 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i3_LC_22_7_3 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i3_LC_22_7_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i3_LC_22_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i3_LC_22_7_3  (
            .in0(_gnd_net_),
            .in1(N__82112),
            .in2(_gnd_net_),
            .in3(N__81735),
            .lcout(\quad_counter1.millisecond_counter_3 ),
            .ltout(),
            .carryin(\quad_counter1.n30173 ),
            .carryout(\quad_counter1.n30174 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i4_LC_22_7_4 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i4_LC_22_7_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i4_LC_22_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i4_LC_22_7_4  (
            .in0(_gnd_net_),
            .in1(N__81722),
            .in2(_gnd_net_),
            .in3(N__81711),
            .lcout(\quad_counter1.millisecond_counter_4 ),
            .ltout(),
            .carryin(\quad_counter1.n30174 ),
            .carryout(\quad_counter1.n30175 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i5_LC_22_7_5 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i5_LC_22_7_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i5_LC_22_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i5_LC_22_7_5  (
            .in0(_gnd_net_),
            .in1(N__82439),
            .in2(_gnd_net_),
            .in3(N__81708),
            .lcout(\quad_counter1.millisecond_counter_5 ),
            .ltout(),
            .carryin(\quad_counter1.n30175 ),
            .carryout(\quad_counter1.n30176 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i6_LC_22_7_6 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i6_LC_22_7_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i6_LC_22_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i6_LC_22_7_6  (
            .in0(_gnd_net_),
            .in1(N__81698),
            .in2(_gnd_net_),
            .in3(N__81687),
            .lcout(\quad_counter1.millisecond_counter_6 ),
            .ltout(),
            .carryin(\quad_counter1.n30176 ),
            .carryout(\quad_counter1.n30177 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i7_LC_22_7_7 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i7_LC_22_7_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i7_LC_22_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i7_LC_22_7_7  (
            .in0(_gnd_net_),
            .in1(N__82457),
            .in2(_gnd_net_),
            .in3(N__81684),
            .lcout(\quad_counter1.millisecond_counter_7 ),
            .ltout(),
            .carryin(\quad_counter1.n30177 ),
            .carryout(\quad_counter1.n30178 ),
            .clk(N__97555),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i8_LC_22_8_0 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i8_LC_22_8_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i8_LC_22_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i8_LC_22_8_0  (
            .in0(_gnd_net_),
            .in1(N__89394),
            .in2(_gnd_net_),
            .in3(N__81681),
            .lcout(\quad_counter1.millisecond_counter_8 ),
            .ltout(),
            .carryin(bfn_22_8_0_),
            .carryout(\quad_counter1.n30179 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i9_LC_22_8_1 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i9_LC_22_8_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i9_LC_22_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i9_LC_22_8_1  (
            .in0(_gnd_net_),
            .in1(N__88380),
            .in2(_gnd_net_),
            .in3(N__82014),
            .lcout(\quad_counter1.millisecond_counter_9 ),
            .ltout(),
            .carryin(\quad_counter1.n30179 ),
            .carryout(\quad_counter1.n30180 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i10_LC_22_8_2 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i10_LC_22_8_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i10_LC_22_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i10_LC_22_8_2  (
            .in0(_gnd_net_),
            .in1(N__82410),
            .in2(_gnd_net_),
            .in3(N__82011),
            .lcout(\quad_counter1.millisecond_counter_10 ),
            .ltout(),
            .carryin(\quad_counter1.n30180 ),
            .carryout(\quad_counter1.n30181 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i11_LC_22_8_3 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i11_LC_22_8_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i11_LC_22_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i11_LC_22_8_3  (
            .in0(_gnd_net_),
            .in1(N__81999),
            .in2(_gnd_net_),
            .in3(N__81975),
            .lcout(\quad_counter1.millisecond_counter_11 ),
            .ltout(),
            .carryin(\quad_counter1.n30181 ),
            .carryout(\quad_counter1.n30182 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i12_LC_22_8_4 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i12_LC_22_8_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i12_LC_22_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i12_LC_22_8_4  (
            .in0(_gnd_net_),
            .in1(N__81960),
            .in2(_gnd_net_),
            .in3(N__81933),
            .lcout(\quad_counter1.millisecond_counter_12 ),
            .ltout(),
            .carryin(\quad_counter1.n30182 ),
            .carryout(\quad_counter1.n30183 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i13_LC_22_8_5 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i13_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i13_LC_22_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i13_LC_22_8_5  (
            .in0(_gnd_net_),
            .in1(N__81909),
            .in2(_gnd_net_),
            .in3(N__81882),
            .lcout(\quad_counter1.millisecond_counter_13 ),
            .ltout(),
            .carryin(\quad_counter1.n30183 ),
            .carryout(\quad_counter1.n30184 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i14_LC_22_8_6 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i14_LC_22_8_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i14_LC_22_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i14_LC_22_8_6  (
            .in0(_gnd_net_),
            .in1(N__81860),
            .in2(_gnd_net_),
            .in3(N__81846),
            .lcout(\quad_counter1.millisecond_counter_14 ),
            .ltout(),
            .carryin(\quad_counter1.n30184 ),
            .carryout(\quad_counter1.n30185 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i15_LC_22_8_7 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i15_LC_22_8_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i15_LC_22_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i15_LC_22_8_7  (
            .in0(_gnd_net_),
            .in1(N__81831),
            .in2(_gnd_net_),
            .in3(N__81807),
            .lcout(\quad_counter1.millisecond_counter_15 ),
            .ltout(),
            .carryin(\quad_counter1.n30185 ),
            .carryout(\quad_counter1.n30186 ),
            .clk(N__97558),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i16_LC_22_9_0 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i16_LC_22_9_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i16_LC_22_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i16_LC_22_9_0  (
            .in0(_gnd_net_),
            .in1(N__81787),
            .in2(_gnd_net_),
            .in3(N__81765),
            .lcout(\quad_counter1.millisecond_counter_16 ),
            .ltout(),
            .carryin(bfn_22_9_0_),
            .carryout(\quad_counter1.n30187 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i17_LC_22_9_1 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i17_LC_22_9_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i17_LC_22_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i17_LC_22_9_1  (
            .in0(_gnd_net_),
            .in1(N__86946),
            .in2(_gnd_net_),
            .in3(N__82044),
            .lcout(\quad_counter1.millisecond_counter_17 ),
            .ltout(),
            .carryin(\quad_counter1.n30187 ),
            .carryout(\quad_counter1.n30188 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i18_LC_22_9_2 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i18_LC_22_9_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i18_LC_22_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i18_LC_22_9_2  (
            .in0(_gnd_net_),
            .in1(N__86905),
            .in2(_gnd_net_),
            .in3(N__82041),
            .lcout(\quad_counter1.millisecond_counter_18 ),
            .ltout(),
            .carryin(\quad_counter1.n30188 ),
            .carryout(\quad_counter1.n30189 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i19_LC_22_9_3 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i19_LC_22_9_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i19_LC_22_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i19_LC_22_9_3  (
            .in0(_gnd_net_),
            .in1(N__88125),
            .in2(_gnd_net_),
            .in3(N__82038),
            .lcout(\quad_counter1.millisecond_counter_19 ),
            .ltout(),
            .carryin(\quad_counter1.n30189 ),
            .carryout(\quad_counter1.n30190 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i20_LC_22_9_4 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i20_LC_22_9_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i20_LC_22_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i20_LC_22_9_4  (
            .in0(_gnd_net_),
            .in1(N__88478),
            .in2(_gnd_net_),
            .in3(N__82035),
            .lcout(\quad_counter1.millisecond_counter_20 ),
            .ltout(),
            .carryin(\quad_counter1.n30190 ),
            .carryout(\quad_counter1.n30191 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i21_LC_22_9_5 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i21_LC_22_9_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i21_LC_22_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i21_LC_22_9_5  (
            .in0(_gnd_net_),
            .in1(N__93485),
            .in2(_gnd_net_),
            .in3(N__82032),
            .lcout(\quad_counter1.millisecond_counter_21 ),
            .ltout(),
            .carryin(\quad_counter1.n30191 ),
            .carryout(\quad_counter1.n30192 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i22_LC_22_9_6 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i22_LC_22_9_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i22_LC_22_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i22_LC_22_9_6  (
            .in0(_gnd_net_),
            .in1(N__95202),
            .in2(_gnd_net_),
            .in3(N__82029),
            .lcout(\quad_counter1.millisecond_counter_22 ),
            .ltout(),
            .carryin(\quad_counter1.n30192 ),
            .carryout(\quad_counter1.n30193 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i23_LC_22_9_7 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i23_LC_22_9_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i23_LC_22_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i23_LC_22_9_7  (
            .in0(_gnd_net_),
            .in1(N__99916),
            .in2(_gnd_net_),
            .in3(N__82026),
            .lcout(\quad_counter1.millisecond_counter_23 ),
            .ltout(),
            .carryin(\quad_counter1.n30193 ),
            .carryout(\quad_counter1.n30194 ),
            .clk(N__97565),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i24_LC_22_10_0 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i24_LC_22_10_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i24_LC_22_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i24_LC_22_10_0  (
            .in0(_gnd_net_),
            .in1(N__95307),
            .in2(_gnd_net_),
            .in3(N__82023),
            .lcout(\quad_counter1.millisecond_counter_24 ),
            .ltout(),
            .carryin(bfn_22_10_0_),
            .carryout(\quad_counter1.n30195 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i25_LC_22_10_1 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i25_LC_22_10_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i25_LC_22_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i25_LC_22_10_1  (
            .in0(_gnd_net_),
            .in1(N__93093),
            .in2(_gnd_net_),
            .in3(N__82020),
            .lcout(\quad_counter1.millisecond_counter_25 ),
            .ltout(),
            .carryin(\quad_counter1.n30195 ),
            .carryout(\quad_counter1.n30196 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i26_LC_22_10_2 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i26_LC_22_10_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i26_LC_22_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i26_LC_22_10_2  (
            .in0(_gnd_net_),
            .in1(N__93054),
            .in2(_gnd_net_),
            .in3(N__82017),
            .lcout(\quad_counter1.millisecond_counter_26 ),
            .ltout(),
            .carryin(\quad_counter1.n30196 ),
            .carryout(\quad_counter1.n30197 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i27_LC_22_10_3 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i27_LC_22_10_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i27_LC_22_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i27_LC_22_10_3  (
            .in0(_gnd_net_),
            .in1(N__93012),
            .in2(_gnd_net_),
            .in3(N__82077),
            .lcout(\quad_counter1.millisecond_counter_27 ),
            .ltout(),
            .carryin(\quad_counter1.n30197 ),
            .carryout(\quad_counter1.n30198 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i28_LC_22_10_4 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i28_LC_22_10_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i28_LC_22_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i28_LC_22_10_4  (
            .in0(_gnd_net_),
            .in1(N__92973),
            .in2(_gnd_net_),
            .in3(N__82074),
            .lcout(\quad_counter1.millisecond_counter_28 ),
            .ltout(),
            .carryin(\quad_counter1.n30198 ),
            .carryout(\quad_counter1.n30199 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i29_LC_22_10_5 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i29_LC_22_10_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i29_LC_22_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i29_LC_22_10_5  (
            .in0(_gnd_net_),
            .in1(N__92937),
            .in2(_gnd_net_),
            .in3(N__82071),
            .lcout(\quad_counter1.millisecond_counter_29 ),
            .ltout(),
            .carryin(\quad_counter1.n30199 ),
            .carryout(\quad_counter1.n30200 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i30_LC_22_10_6 .C_ON=1'b1;
    defparam \quad_counter1.millisecond_counter_1426__i30_LC_22_10_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i30_LC_22_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i30_LC_22_10_6  (
            .in0(_gnd_net_),
            .in1(N__93369),
            .in2(_gnd_net_),
            .in3(N__82068),
            .lcout(\quad_counter1.millisecond_counter_30 ),
            .ltout(),
            .carryin(\quad_counter1.n30200 ),
            .carryout(\quad_counter1.n30201 ),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.millisecond_counter_1426__i31_LC_22_10_7 .C_ON=1'b0;
    defparam \quad_counter1.millisecond_counter_1426__i31_LC_22_10_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter1.millisecond_counter_1426__i31_LC_22_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.millisecond_counter_1426__i31_LC_22_10_7  (
            .in0(_gnd_net_),
            .in1(N__93330),
            .in2(_gnd_net_),
            .in3(N__82065),
            .lcout(\quad_counter1.millisecond_counter_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97574),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_2_lut_LC_22_11_0 .C_ON=1'b1;
    defparam \quad_counter1.add_8377_2_lut_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_2_lut_LC_22_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_8377_2_lut_LC_22_11_0  (
            .in0(_gnd_net_),
            .in1(N__89395),
            .in2(_gnd_net_),
            .in3(N__82062),
            .lcout(\quad_counter1.n12936 ),
            .ltout(),
            .carryin(bfn_22_11_0_),
            .carryout(\quad_counter1.n30447 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_3_lut_LC_22_11_1 .C_ON=1'b1;
    defparam \quad_counter1.add_8377_3_lut_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_3_lut_LC_22_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_8377_3_lut_LC_22_11_1  (
            .in0(_gnd_net_),
            .in1(N__98965),
            .in2(N__89365),
            .in3(N__82059),
            .lcout(\quad_counter1.n12935 ),
            .ltout(),
            .carryin(\quad_counter1.n30447 ),
            .carryout(\quad_counter1.n30448 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_4_lut_LC_22_11_2 .C_ON=1'b1;
    defparam \quad_counter1.add_8377_4_lut_LC_22_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_4_lut_LC_22_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.add_8377_4_lut_LC_22_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__89290),
            .in3(N__82056),
            .lcout(\quad_counter1.n12934 ),
            .ltout(),
            .carryin(\quad_counter1.n30448 ),
            .carryout(\quad_counter1.n30449 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_5_lut_LC_22_11_3 .C_ON=1'b1;
    defparam \quad_counter1.add_8377_5_lut_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_5_lut_LC_22_11_3 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter1.add_8377_5_lut_LC_22_11_3  (
            .in0(N__82053),
            .in1(_gnd_net_),
            .in2(N__89317),
            .in3(N__82047),
            .lcout(\quad_counter1.n10_adj_4454 ),
            .ltout(),
            .carryin(\quad_counter1.n30449 ),
            .carryout(\quad_counter1.n30450 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_6_lut_LC_22_11_4 .C_ON=1'b1;
    defparam \quad_counter1.add_8377_6_lut_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_6_lut_LC_22_11_4 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter1.add_8377_6_lut_LC_22_11_4  (
            .in0(N__82161),
            .in1(_gnd_net_),
            .in2(N__89230),
            .in3(N__82170),
            .lcout(\quad_counter1.n35987 ),
            .ltout(),
            .carryin(\quad_counter1.n30450 ),
            .carryout(\quad_counter1.n30451 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_7_lut_LC_22_11_5 .C_ON=1'b1;
    defparam \quad_counter1.add_8377_7_lut_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_7_lut_LC_22_11_5 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter1.add_8377_7_lut_LC_22_11_5  (
            .in0(N__82167),
            .in1(N__89263),
            .in2(_gnd_net_),
            .in3(N__82155),
            .lcout(\quad_counter1.n8_adj_4453 ),
            .ltout(),
            .carryin(\quad_counter1.n30451 ),
            .carryout(\quad_counter1.n30452 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.add_8377_8_lut_LC_22_11_6 .C_ON=1'b0;
    defparam \quad_counter1.add_8377_8_lut_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.add_8377_8_lut_LC_22_11_6 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \quad_counter1.add_8377_8_lut_LC_22_11_6  (
            .in0(N__82152),
            .in1(N__89338),
            .in2(_gnd_net_),
            .in3(N__82146),
            .lcout(\quad_counter1.n9_adj_4452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30644_3_lut_LC_22_11_7 .C_ON=1'b0;
    defparam \quad_counter1.i30644_3_lut_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30644_3_lut_LC_22_11_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \quad_counter1.i30644_3_lut_LC_22_11_7  (
            .in0(N__82143),
            .in1(N__82137),
            .in2(_gnd_net_),
            .in3(N__82131),
            .lcout(\quad_counter1.n35986 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i13_4_lut_adj_1293_LC_22_12_0 .C_ON=1'b0;
    defparam \quad_counter1.i13_4_lut_adj_1293_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i13_4_lut_adj_1293_LC_22_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i13_4_lut_adj_1293_LC_22_12_0  (
            .in0(N__88755),
            .in1(N__89124),
            .in2(N__88851),
            .in3(N__88920),
            .lcout(),
            .ltout(\quad_counter1.n31_adj_4461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i16_4_lut_adj_1298_LC_22_12_1 .C_ON=1'b0;
    defparam \quad_counter1.i16_4_lut_adj_1298_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i16_4_lut_adj_1298_LC_22_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i16_4_lut_adj_1298_LC_22_12_1  (
            .in0(N__89094),
            .in1(N__88488),
            .in2(N__82125),
            .in3(N__88788),
            .lcout(),
            .ltout(\quad_counter1.n34_adj_4465_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i47_4_lut_LC_22_12_2 .C_ON=1'b0;
    defparam \quad_counter1.i47_4_lut_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i47_4_lut_LC_22_12_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \quad_counter1.i47_4_lut_LC_22_12_2  (
            .in0(N__83376),
            .in1(N__82122),
            .in2(N__82116),
            .in3(N__89028),
            .lcout(),
            .ltout(\quad_counter1.n34207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_3_lut_LC_22_12_3 .C_ON=1'b0;
    defparam \quad_counter1.i2_3_lut_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_3_lut_LC_22_12_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \quad_counter1.i2_3_lut_LC_22_12_3  (
            .in0(_gnd_net_),
            .in1(N__82113),
            .in2(N__82098),
            .in3(N__82095),
            .lcout(),
            .ltout(\quad_counter1.n34519_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1300_LC_22_12_4 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1300_LC_22_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1300_LC_22_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1300_LC_22_12_4  (
            .in0(N__82473),
            .in1(N__82458),
            .in2(N__82443),
            .in3(N__82440),
            .lcout(\quad_counter1.n12_adj_4467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_2_lut_LC_22_13_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_2_lut_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_2_lut_LC_22_13_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2286_2_lut_LC_22_13_0  (
            .in0(N__82419),
            .in1(N__82418),
            .in2(N__82210),
            .in3(N__82383),
            .lcout(\quad_counter1.n3419 ),
            .ltout(),
            .carryin(bfn_22_13_0_),
            .carryout(\quad_counter1.n30654 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_3_lut_LC_22_13_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_3_lut_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_3_lut_LC_22_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_3_lut_LC_22_13_1  (
            .in0(N__82380),
            .in1(N__82379),
            .in2(N__82836),
            .in3(N__82356),
            .lcout(\quad_counter1.n3418 ),
            .ltout(),
            .carryin(\quad_counter1.n30654 ),
            .carryout(\quad_counter1.n30655 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_4_lut_LC_22_13_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_4_lut_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_4_lut_LC_22_13_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2286_4_lut_LC_22_13_2  (
            .in0(N__82353),
            .in1(N__82352),
            .in2(N__82211),
            .in3(N__82326),
            .lcout(\quad_counter1.n3417 ),
            .ltout(),
            .carryin(\quad_counter1.n30655 ),
            .carryout(\quad_counter1.n30656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_5_lut_LC_22_13_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_5_lut_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_5_lut_LC_22_13_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2286_5_lut_LC_22_13_3  (
            .in0(N__82323),
            .in1(N__82322),
            .in2(N__82214),
            .in3(N__82299),
            .lcout(\quad_counter1.n3416 ),
            .ltout(),
            .carryin(\quad_counter1.n30656 ),
            .carryout(\quad_counter1.n30657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_6_lut_LC_22_13_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_6_lut_LC_22_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_6_lut_LC_22_13_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2286_6_lut_LC_22_13_4  (
            .in0(N__82296),
            .in1(N__82295),
            .in2(N__82212),
            .in3(N__82272),
            .lcout(\quad_counter1.n3415 ),
            .ltout(),
            .carryin(\quad_counter1.n30657 ),
            .carryout(\quad_counter1.n30658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_7_lut_LC_22_13_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_7_lut_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_7_lut_LC_22_13_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2286_7_lut_LC_22_13_5  (
            .in0(N__82269),
            .in1(N__82268),
            .in2(N__82215),
            .in3(N__82245),
            .lcout(\quad_counter1.n3414 ),
            .ltout(),
            .carryin(\quad_counter1.n30658 ),
            .carryout(\quad_counter1.n30659 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_8_lut_LC_22_13_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_8_lut_LC_22_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_8_lut_LC_22_13_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2286_8_lut_LC_22_13_6  (
            .in0(N__82242),
            .in1(N__82241),
            .in2(N__82213),
            .in3(N__82173),
            .lcout(\quad_counter1.n3413 ),
            .ltout(),
            .carryin(\quad_counter1.n30659 ),
            .carryout(\quad_counter1.n30660 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_9_lut_LC_22_13_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_9_lut_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_9_lut_LC_22_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_9_lut_LC_22_13_7  (
            .in0(N__82728),
            .in1(N__82727),
            .in2(N__82837),
            .in3(N__82704),
            .lcout(\quad_counter1.n3412 ),
            .ltout(),
            .carryin(\quad_counter1.n30660 ),
            .carryout(\quad_counter1.n30661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_10_lut_LC_22_14_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_10_lut_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_10_lut_LC_22_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_10_lut_LC_22_14_0  (
            .in0(N__82701),
            .in1(N__82700),
            .in2(N__82838),
            .in3(N__82677),
            .lcout(\quad_counter1.n3411 ),
            .ltout(),
            .carryin(bfn_22_14_0_),
            .carryout(\quad_counter1.n30662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_11_lut_LC_22_14_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_11_lut_LC_22_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_11_lut_LC_22_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_11_lut_LC_22_14_1  (
            .in0(N__82674),
            .in1(N__82673),
            .in2(N__82842),
            .in3(N__82647),
            .lcout(\quad_counter1.n3410 ),
            .ltout(),
            .carryin(\quad_counter1.n30662 ),
            .carryout(\quad_counter1.n30663 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_12_lut_LC_22_14_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_12_lut_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_12_lut_LC_22_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_12_lut_LC_22_14_2  (
            .in0(N__82644),
            .in1(N__82643),
            .in2(N__82839),
            .in3(N__82620),
            .lcout(\quad_counter1.n3409 ),
            .ltout(),
            .carryin(\quad_counter1.n30663 ),
            .carryout(\quad_counter1.n30664 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_13_lut_LC_22_14_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_13_lut_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_13_lut_LC_22_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_13_lut_LC_22_14_3  (
            .in0(N__82617),
            .in1(N__82616),
            .in2(N__82843),
            .in3(N__82590),
            .lcout(\quad_counter1.n3408 ),
            .ltout(),
            .carryin(\quad_counter1.n30664 ),
            .carryout(\quad_counter1.n30665 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_14_lut_LC_22_14_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_14_lut_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_14_lut_LC_22_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_14_lut_LC_22_14_4  (
            .in0(N__82587),
            .in1(N__82586),
            .in2(N__82840),
            .in3(N__82563),
            .lcout(\quad_counter1.n3407 ),
            .ltout(),
            .carryin(\quad_counter1.n30665 ),
            .carryout(\quad_counter1.n30666 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_15_lut_LC_22_14_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_15_lut_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_15_lut_LC_22_14_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_15_lut_LC_22_14_5  (
            .in0(N__82560),
            .in1(N__82559),
            .in2(N__82844),
            .in3(N__82533),
            .lcout(\quad_counter1.n3406 ),
            .ltout(),
            .carryin(\quad_counter1.n30666 ),
            .carryout(\quad_counter1.n30667 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_16_lut_LC_22_14_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_16_lut_LC_22_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_16_lut_LC_22_14_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_16_lut_LC_22_14_6  (
            .in0(N__82530),
            .in1(N__82529),
            .in2(N__82841),
            .in3(N__82503),
            .lcout(\quad_counter1.n3405 ),
            .ltout(),
            .carryin(\quad_counter1.n30667 ),
            .carryout(\quad_counter1.n30668 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_17_lut_LC_22_14_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_17_lut_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_17_lut_LC_22_14_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_17_lut_LC_22_14_7  (
            .in0(N__82500),
            .in1(N__82499),
            .in2(N__82845),
            .in3(N__82476),
            .lcout(\quad_counter1.n3404 ),
            .ltout(),
            .carryin(\quad_counter1.n30668 ),
            .carryout(\quad_counter1.n30669 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_18_lut_LC_22_15_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_18_lut_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_18_lut_LC_22_15_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_18_lut_LC_22_15_0  (
            .in0(N__83013),
            .in1(N__83012),
            .in2(N__82846),
            .in3(N__82989),
            .lcout(\quad_counter1.n3403 ),
            .ltout(),
            .carryin(bfn_22_15_0_),
            .carryout(\quad_counter1.n30670 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_19_lut_LC_22_15_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_19_lut_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_19_lut_LC_22_15_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_19_lut_LC_22_15_1  (
            .in0(N__82985),
            .in1(N__82986),
            .in2(N__82849),
            .in3(N__82959),
            .lcout(\quad_counter1.n3402 ),
            .ltout(),
            .carryin(\quad_counter1.n30670 ),
            .carryout(\quad_counter1.n30671 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_20_lut_LC_22_15_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_20_lut_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_20_lut_LC_22_15_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_20_lut_LC_22_15_2  (
            .in0(N__82956),
            .in1(N__82955),
            .in2(N__82847),
            .in3(N__82932),
            .lcout(\quad_counter1.n3401 ),
            .ltout(),
            .carryin(\quad_counter1.n30671 ),
            .carryout(\quad_counter1.n30672 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_21_lut_LC_22_15_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_21_lut_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_21_lut_LC_22_15_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_21_lut_LC_22_15_3  (
            .in0(N__82929),
            .in1(N__82928),
            .in2(N__82850),
            .in3(N__82905),
            .lcout(\quad_counter1.n3400 ),
            .ltout(),
            .carryin(\quad_counter1.n30672 ),
            .carryout(\quad_counter1.n30673 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_22_lut_LC_22_15_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2286_22_lut_LC_22_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_22_lut_LC_22_15_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_22_lut_LC_22_15_4  (
            .in0(N__82902),
            .in1(N__82901),
            .in2(N__82848),
            .in3(N__82878),
            .lcout(\quad_counter1.n3399 ),
            .ltout(),
            .carryin(\quad_counter1.n30673 ),
            .carryout(\quad_counter1.n30674 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2286_23_lut_LC_22_15_5 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_2286_23_lut_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2286_23_lut_LC_22_15_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2286_23_lut_LC_22_15_5  (
            .in0(N__82874),
            .in1(N__82875),
            .in2(N__82851),
            .in3(N__82740),
            .lcout(\quad_counter1.n3398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1250_LC_22_15_6 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1250_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1250_LC_22_15_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1250_LC_22_15_6  (
            .in0(N__88804),
            .in1(N__89080),
            .in2(N__88611),
            .in3(N__88546),
            .lcout(\quad_counter1.n27_adj_4429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i11_4_lut_adj_1248_LC_22_15_7 .C_ON=1'b0;
    defparam \quad_counter1.i11_4_lut_adj_1248_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i11_4_lut_adj_1248_LC_22_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i11_4_lut_adj_1248_LC_22_15_7  (
            .in0(N__89110),
            .in1(N__82737),
            .in2(N__89145),
            .in3(N__88741),
            .lcout(\quad_counter1.n28_adj_4427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i15_4_lut_adj_1299_LC_22_16_2 .C_ON=1'b0;
    defparam \quad_counter1.i15_4_lut_adj_1299_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i15_4_lut_adj_1299_LC_22_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i15_4_lut_adj_1299_LC_22_16_2  (
            .in0(N__89208),
            .in1(N__88584),
            .in2(N__88821),
            .in3(N__89040),
            .lcout(\quad_counter1.n33_adj_4466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_10_i3_2_lut_LC_22_16_3 .C_ON=1'b0;
    defparam \c0.select_369_Select_10_i3_2_lut_LC_22_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_10_i3_2_lut_LC_22_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_10_i3_2_lut_LC_22_16_3  (
            .in0(_gnd_net_),
            .in1(N__91841),
            .in2(_gnd_net_),
            .in3(N__94689),
            .lcout(\c0.n3_adj_4589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30396_4_lut_LC_22_17_0 .C_ON=1'b0;
    defparam \c0.i30396_4_lut_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i30396_4_lut_LC_22_17_0 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.i30396_4_lut_LC_22_17_0  (
            .in0(N__94206),
            .in1(N__83367),
            .in2(N__90871),
            .in3(N__90758),
            .lcout(n35823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__3__5298_LC_22_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__3__5298_LC_22_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__3__5298_LC_22_17_1 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \c0.data_out_frame_28__3__5298_LC_22_17_1  (
            .in0(N__93969),
            .in1(N__83343),
            .in2(N__85276),
            .in3(N__84559),
            .lcout(data_out_frame_28_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1466_LC_22_17_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1466_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1466_LC_22_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1466_LC_22_17_6  (
            .in0(N__83330),
            .in1(N__83280),
            .in2(N__83228),
            .in3(N__83169),
            .lcout(\c0.n33353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1953_LC_22_17_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1953_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1953_LC_22_17_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1953_LC_22_17_7  (
            .in0(N__96758),
            .in1(N__100206),
            .in2(N__93803),
            .in3(N__100806),
            .lcout(\c0.n17570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_22_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_22_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1556_LC_22_18_0  (
            .in0(N__83139),
            .in1(N__83483),
            .in2(N__83151),
            .in3(N__83424),
            .lcout(\c0.n15729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1431_LC_22_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1431_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1431_LC_22_18_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1431_LC_22_18_1  (
            .in0(_gnd_net_),
            .in1(N__83147),
            .in2(_gnd_net_),
            .in3(N__83138),
            .lcout(\c0.n31446 ),
            .ltout(\c0.n31446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1432_LC_22_18_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1432_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1432_LC_22_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1432_LC_22_18_2  (
            .in0(_gnd_net_),
            .in1(N__83085),
            .in2(N__83067),
            .in3(N__83064),
            .lcout(\c0.n31928 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_2054_LC_22_18_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_2054_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_2054_LC_22_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_2054_LC_22_18_6  (
            .in0(N__84759),
            .in1(N__85322),
            .in2(N__86600),
            .in3(N__85541),
            .lcout(\c0.n32372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_22_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_22_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_22_19_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i13_LC_22_19_1  (
            .in0(N__84245),
            .in1(N__83868),
            .in2(N__83595),
            .in3(N__87126),
            .lcout(data_in_frame_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_22_19_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_22_19_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_3_lut_LC_22_19_2  (
            .in0(N__84760),
            .in1(N__85321),
            .in2(_gnd_net_),
            .in3(N__86645),
            .lcout(\c0.n33746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1708_LC_22_19_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1708_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1708_LC_22_19_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1708_LC_22_19_4  (
            .in0(N__90381),
            .in1(N__90095),
            .in2(_gnd_net_),
            .in3(N__95790),
            .lcout(n17453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_22_19_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_22_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_22_19_6  (
            .in0(N__96543),
            .in1(N__97824),
            .in2(_gnd_net_),
            .in3(N__96168),
            .lcout(\c0.n26_adj_4654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1765_LC_22_20_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1765_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1765_LC_22_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1765_LC_22_20_0  (
            .in0(N__83534),
            .in1(N__94311),
            .in2(N__85840),
            .in3(N__97975),
            .lcout(\c0.n33861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1718_LC_22_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1718_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1718_LC_22_20_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1718_LC_22_20_1  (
            .in0(N__94076),
            .in1(N__83481),
            .in2(_gnd_net_),
            .in3(N__83421),
            .lcout(\c0.n32290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.encoder1_position_7__I_0_5546_2_lut_LC_22_20_4 .C_ON=1'b0;
    defparam \c0.encoder1_position_7__I_0_5546_2_lut_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.encoder1_position_7__I_0_5546_2_lut_LC_22_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.encoder1_position_7__I_0_5546_2_lut_LC_22_20_4  (
            .in0(_gnd_net_),
            .in1(N__94310),
            .in2(_gnd_net_),
            .in3(N__97974),
            .lcout(),
            .ltout(\c0.data_out_frame_29__7__N_658_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1461_LC_22_20_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1461_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1461_LC_22_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1461_LC_22_20_5  (
            .in0(N__83385),
            .in1(N__85510),
            .in2(N__83379),
            .in3(N__90573),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1743_LC_22_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1743_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1743_LC_22_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1743_LC_22_20_6  (
            .in0(N__85511),
            .in1(N__85463),
            .in2(N__85401),
            .in3(N__85380),
            .lcout(\c0.n18469 ),
            .ltout(\c0.n18469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1486_LC_22_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1486_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1486_LC_22_20_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1486_LC_22_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__85326),
            .in3(N__90574),
            .lcout(\c0.n31466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1722_LC_22_21_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1722_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1722_LC_22_21_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1722_LC_22_21_0  (
            .in0(N__85323),
            .in1(N__101038),
            .in2(_gnd_net_),
            .in3(N__101101),
            .lcout(\c0.n10_adj_4528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1394_LC_22_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1394_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1394_LC_22_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1394_LC_22_21_1  (
            .in0(N__84769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86607),
            .lcout(),
            .ltout(\c0.n18241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1354_LC_22_21_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1354_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1354_LC_22_21_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1354_LC_22_21_2  (
            .in0(N__98243),
            .in1(N__94955),
            .in2(N__85299),
            .in3(N__96491),
            .lcout(),
            .ltout(\c0.n14_adj_4527_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1355_LC_22_21_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1355_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1355_LC_22_21_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1355_LC_22_21_3  (
            .in0(N__85296),
            .in1(N__94262),
            .in2(N__85290),
            .in3(N__86448),
            .lcout(\c0.n33529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_22_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1751_LC_22_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1751_LC_22_21_4  (
            .in0(N__90929),
            .in1(N__100929),
            .in2(_gnd_net_),
            .in3(N__90578),
            .lcout(\c0.n31511 ),
            .ltout(\c0.n31511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1456_LC_22_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1456_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1456_LC_22_21_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1456_LC_22_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__85287),
            .in3(N__90930),
            .lcout(\c0.n33687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_13__1__5420_LC_22_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame_13__1__5420_LC_22_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_13__1__5420_LC_22_21_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \c0.data_out_frame_13__1__5420_LC_22_21_7  (
            .in0(N__84269),
            .in1(N__85273),
            .in2(N__84774),
            .in3(N__84560),
            .lcout(data_out_frame_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1755_LC_22_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1755_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1755_LC_22_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1755_LC_22_22_1  (
            .in0(N__86186),
            .in1(N__86310),
            .in2(N__85857),
            .in3(N__86491),
            .lcout(),
            .ltout(\c0.n6_adj_4558_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1437_LC_22_22_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1437_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1437_LC_22_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1437_LC_22_22_2  (
            .in0(N__85626),
            .in1(N__85830),
            .in2(N__85791),
            .in3(N__85788),
            .lcout(\c0.n18898 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_LC_22_22_3 .C_ON=1'b0;
    defparam \c0.i15_2_lut_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_LC_22_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i15_2_lut_LC_22_22_3  (
            .in0(_gnd_net_),
            .in1(N__94982),
            .in2(_gnd_net_),
            .in3(N__100165),
            .lcout(\c0.n32424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1741_LC_22_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1741_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1741_LC_22_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1741_LC_22_22_4  (
            .in0(N__85735),
            .in1(N__86443),
            .in2(_gnd_net_),
            .in3(N__94362),
            .lcout(\c0.n18499 ),
            .ltout(\c0.n18499_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1942_LC_22_22_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1942_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1942_LC_22_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1942_LC_22_22_5  (
            .in0(N__90448),
            .in1(N__94513),
            .in2(N__85695),
            .in3(N__94983),
            .lcout(\c0.n35426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1439_LC_22_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1439_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1439_LC_22_22_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1439_LC_22_22_6  (
            .in0(_gnd_net_),
            .in1(N__86444),
            .in2(_gnd_net_),
            .in3(N__94363),
            .lcout(),
            .ltout(\c0.n33569_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1421_LC_22_22_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1421_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1421_LC_22_22_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1421_LC_22_22_7  (
            .in0(N__98247),
            .in1(N__86606),
            .in2(N__85692),
            .in3(N__86646),
            .lcout(\c0.n21_adj_4551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1547_LC_22_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1547_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1547_LC_22_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1547_LC_22_23_1  (
            .in0(N__86637),
            .in1(N__85537),
            .in2(N__94534),
            .in3(N__86610),
            .lcout(\c0.n15775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1478_LC_22_23_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1478_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1478_LC_22_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1478_LC_22_23_2  (
            .in0(N__85688),
            .in1(N__86540),
            .in2(N__85625),
            .in3(N__85548),
            .lcout(\c0.n33897 ),
            .ltout(\c0.n33897_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1543_LC_22_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1543_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1543_LC_22_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1543_LC_22_23_3  (
            .in0(N__86636),
            .in1(N__86609),
            .in2(N__86544),
            .in3(N__98335),
            .lcout(\c0.n32333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1438_LC_22_23_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1438_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1438_LC_22_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1438_LC_22_23_4  (
            .in0(N__86309),
            .in1(N__86541),
            .in2(N__86529),
            .in3(N__86490),
            .lcout(\c0.n18895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1744_LC_22_23_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1744_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1744_LC_22_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1744_LC_22_23_5  (
            .in0(N__86419),
            .in1(N__86185),
            .in2(N__86363),
            .in3(N__86308),
            .lcout(\c0.n33318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1471_LC_22_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1471_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1471_LC_22_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1471_LC_22_23_7  (
            .in0(_gnd_net_),
            .in1(N__86271),
            .in2(_gnd_net_),
            .in3(N__86184),
            .lcout(\c0.n33487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i28_LC_22_25_2 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i28_LC_22_25_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i28_LC_22_25_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i28_LC_22_25_2  (
            .in0(N__86142),
            .in1(N__86214),
            .in2(_gnd_net_),
            .in3(N__86181),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97780),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.count_i0_i26_LC_22_25_6 .C_ON=1'b0;
    defparam \quad_counter0.count_i0_i26_LC_22_25_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.count_i0_i26_LC_22_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \quad_counter0.count_i0_i26_LC_22_25_6  (
            .in0(N__86141),
            .in1(N__85941),
            .in2(_gnd_net_),
            .in3(N__85900),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97780),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_3_i3_2_lut_LC_23_4_3 .C_ON=1'b0;
    defparam \c0.select_369_Select_3_i3_2_lut_LC_23_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_3_i3_2_lut_LC_23_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_3_i3_2_lut_LC_23_4_3  (
            .in0(_gnd_net_),
            .in1(N__91298),
            .in2(_gnd_net_),
            .in3(N__94747),
            .lcout(\c0.n3_adj_4581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_4_i3_2_lut_LC_23_5_1 .C_ON=1'b0;
    defparam \c0.select_369_Select_4_i3_2_lut_LC_23_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_4_i3_2_lut_LC_23_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_4_i3_2_lut_LC_23_5_1  (
            .in0(_gnd_net_),
            .in1(N__91405),
            .in2(_gnd_net_),
            .in3(N__94833),
            .lcout(\c0.n3_adj_4583 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_82_i9_2_lut_3_lut_LC_23_6_0 .C_ON=1'b0;
    defparam \c0.equal_82_i9_2_lut_3_lut_LC_23_6_0 .SEQ_MODE=4'b0000;
    defparam \c0.equal_82_i9_2_lut_3_lut_LC_23_6_0 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.equal_82_i9_2_lut_3_lut_LC_23_6_0  (
            .in0(N__93198),
            .in1(N__91202),
            .in2(_gnd_net_),
            .in3(N__91032),
            .lcout(\c0.n9_adj_4493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23555_2_lut_LC_23_6_3 .C_ON=1'b0;
    defparam \quad_counter1.i23555_2_lut_LC_23_6_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23555_2_lut_LC_23_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23555_2_lut_LC_23_6_3  (
            .in0(_gnd_net_),
            .in1(N__86869),
            .in2(_gnd_net_),
            .in3(N__86947),
            .lcout(),
            .ltout(\quad_counter1.n28271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_LC_23_6_4 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_LC_23_6_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_LC_23_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_LC_23_6_4  (
            .in0(N__86813),
            .in1(N__87680),
            .in2(N__86925),
            .in3(N__86762),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4423_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_4_lut_adj_1281_LC_23_6_5 .C_ON=1'b0;
    defparam \quad_counter1.i2_4_lut_adj_1281_LC_23_6_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_4_lut_adj_1281_LC_23_6_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i2_4_lut_adj_1281_LC_23_6_5  (
            .in0(N__86660),
            .in1(N__87967),
            .in2(N__86922),
            .in3(N__86711),
            .lcout(\quad_counter1.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_2_lut_LC_23_7_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_2_lut_LC_23_7_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_2_lut_LC_23_7_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1750_2_lut_LC_23_7_0  (
            .in0(N__86913),
            .in1(N__86912),
            .in2(N__87877),
            .in3(N__86853),
            .lcout(\quad_counter1.n2619 ),
            .ltout(),
            .carryin(bfn_23_7_0_),
            .carryout(\quad_counter1.n30522 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_3_lut_LC_23_7_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_3_lut_LC_23_7_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_3_lut_LC_23_7_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_3_lut_LC_23_7_1  (
            .in0(N__86850),
            .in1(N__86849),
            .in2(N__87947),
            .in3(N__86802),
            .lcout(\quad_counter1.n2618 ),
            .ltout(),
            .carryin(\quad_counter1.n30522 ),
            .carryout(\quad_counter1.n30523 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_4_lut_LC_23_7_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_4_lut_LC_23_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_4_lut_LC_23_7_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1750_4_lut_LC_23_7_2  (
            .in0(N__86799),
            .in1(N__86798),
            .in2(N__87878),
            .in3(N__86751),
            .lcout(\quad_counter1.n2617 ),
            .ltout(),
            .carryin(\quad_counter1.n30523 ),
            .carryout(\quad_counter1.n30524 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_5_lut_LC_23_7_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_5_lut_LC_23_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_5_lut_LC_23_7_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1750_5_lut_LC_23_7_3  (
            .in0(N__86748),
            .in1(N__86747),
            .in2(N__87881),
            .in3(N__86700),
            .lcout(\quad_counter1.n2616 ),
            .ltout(),
            .carryin(\quad_counter1.n30524 ),
            .carryout(\quad_counter1.n30525 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_6_lut_LC_23_7_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_6_lut_LC_23_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_6_lut_LC_23_7_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1750_6_lut_LC_23_7_4  (
            .in0(N__86697),
            .in1(N__86696),
            .in2(N__87879),
            .in3(N__86649),
            .lcout(\quad_counter1.n2615 ),
            .ltout(),
            .carryin(\quad_counter1.n30525 ),
            .carryout(\quad_counter1.n30526 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_7_lut_LC_23_7_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_7_lut_LC_23_7_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_7_lut_LC_23_7_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1750_7_lut_LC_23_7_5  (
            .in0(N__87717),
            .in1(N__87716),
            .in2(N__87882),
            .in3(N__87669),
            .lcout(\quad_counter1.n2614 ),
            .ltout(),
            .carryin(\quad_counter1.n30526 ),
            .carryout(\quad_counter1.n30527 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_8_lut_LC_23_7_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_8_lut_LC_23_7_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_8_lut_LC_23_7_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1750_8_lut_LC_23_7_6  (
            .in0(N__87666),
            .in1(N__87665),
            .in2(N__87880),
            .in3(N__87618),
            .lcout(\quad_counter1.n2613 ),
            .ltout(),
            .carryin(\quad_counter1.n30527 ),
            .carryout(\quad_counter1.n30528 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_9_lut_LC_23_7_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_9_lut_LC_23_7_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_9_lut_LC_23_7_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_9_lut_LC_23_7_7  (
            .in0(N__87615),
            .in1(N__87614),
            .in2(N__87948),
            .in3(N__87567),
            .lcout(\quad_counter1.n2612 ),
            .ltout(),
            .carryin(\quad_counter1.n30528 ),
            .carryout(\quad_counter1.n30529 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_10_lut_LC_23_8_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_10_lut_LC_23_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_10_lut_LC_23_8_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_10_lut_LC_23_8_0  (
            .in0(N__87564),
            .in1(N__87563),
            .in2(N__87935),
            .in3(N__87513),
            .lcout(\quad_counter1.n2611 ),
            .ltout(),
            .carryin(bfn_23_8_0_),
            .carryout(\quad_counter1.n30530 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_11_lut_LC_23_8_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_11_lut_LC_23_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_11_lut_LC_23_8_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_11_lut_LC_23_8_1  (
            .in0(N__87510),
            .in1(N__87509),
            .in2(N__87944),
            .in3(N__87453),
            .lcout(\quad_counter1.n2610 ),
            .ltout(),
            .carryin(\quad_counter1.n30530 ),
            .carryout(\quad_counter1.n30531 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_12_lut_LC_23_8_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_12_lut_LC_23_8_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_12_lut_LC_23_8_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_12_lut_LC_23_8_2  (
            .in0(N__87450),
            .in1(N__87449),
            .in2(N__87936),
            .in3(N__87396),
            .lcout(\quad_counter1.n2609 ),
            .ltout(),
            .carryin(\quad_counter1.n30531 ),
            .carryout(\quad_counter1.n30532 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_13_lut_LC_23_8_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_13_lut_LC_23_8_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_13_lut_LC_23_8_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_13_lut_LC_23_8_3  (
            .in0(N__87393),
            .in1(N__87392),
            .in2(N__87945),
            .in3(N__87336),
            .lcout(\quad_counter1.n2608 ),
            .ltout(),
            .carryin(\quad_counter1.n30532 ),
            .carryout(\quad_counter1.n30533 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_14_lut_LC_23_8_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1750_14_lut_LC_23_8_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_14_lut_LC_23_8_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_14_lut_LC_23_8_4  (
            .in0(N__87333),
            .in1(N__87332),
            .in2(N__87937),
            .in3(N__88008),
            .lcout(\quad_counter1.n2607 ),
            .ltout(),
            .carryin(\quad_counter1.n30533 ),
            .carryout(\quad_counter1.n30534 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1750_15_lut_LC_23_8_5 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1750_15_lut_LC_23_8_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1750_15_lut_LC_23_8_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1750_15_lut_LC_23_8_5  (
            .in0(N__88004),
            .in1(N__88005),
            .in2(N__87946),
            .in3(N__87978),
            .lcout(\quad_counter1.n2606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30706_1_lut_LC_23_8_7 .C_ON=1'b0;
    defparam \quad_counter1.i30706_1_lut_LC_23_8_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30706_1_lut_LC_23_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter1.i30706_1_lut_LC_23_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87911),
            .lcout(\quad_counter1.n36133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_2_lut_LC_23_9_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_2_lut_LC_23_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_2_lut_LC_23_9_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1616_2_lut_LC_23_9_0  (
            .in0(N__88477),
            .in1(N__88476),
            .in2(N__88525),
            .in3(N__87840),
            .lcout(\quad_counter1.n2419 ),
            .ltout(),
            .carryin(bfn_23_9_0_),
            .carryout(\quad_counter1.n30499 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_3_lut_LC_23_9_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_3_lut_LC_23_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_3_lut_LC_23_9_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1616_3_lut_LC_23_9_1  (
            .in0(N__93471),
            .in1(N__93470),
            .in2(N__88442),
            .in3(N__87837),
            .lcout(\quad_counter1.n2418 ),
            .ltout(),
            .carryin(\quad_counter1.n30499 ),
            .carryout(\quad_counter1.n30500 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_4_lut_LC_23_9_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_4_lut_LC_23_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_4_lut_LC_23_9_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1616_4_lut_LC_23_9_2  (
            .in0(N__93441),
            .in1(N__93440),
            .in2(N__88526),
            .in3(N__87810),
            .lcout(\quad_counter1.n2417 ),
            .ltout(),
            .carryin(\quad_counter1.n30500 ),
            .carryout(\quad_counter1.n30501 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_5_lut_LC_23_9_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_5_lut_LC_23_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_5_lut_LC_23_9_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1616_5_lut_LC_23_9_3  (
            .in0(N__93408),
            .in1(N__93407),
            .in2(N__88529),
            .in3(N__87780),
            .lcout(\quad_counter1.n2416 ),
            .ltout(),
            .carryin(\quad_counter1.n30501 ),
            .carryout(\quad_counter1.n30502 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_6_lut_LC_23_9_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_6_lut_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_6_lut_LC_23_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1616_6_lut_LC_23_9_4  (
            .in0(N__93783),
            .in1(N__93782),
            .in2(N__88527),
            .in3(N__87750),
            .lcout(\quad_counter1.n2415 ),
            .ltout(),
            .carryin(\quad_counter1.n30502 ),
            .carryout(\quad_counter1.n30503 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_7_lut_LC_23_9_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_7_lut_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_7_lut_LC_23_9_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1616_7_lut_LC_23_9_5  (
            .in0(N__93755),
            .in1(N__93756),
            .in2(N__88530),
            .in3(N__87720),
            .lcout(\quad_counter1.n2414 ),
            .ltout(),
            .carryin(\quad_counter1.n30503 ),
            .carryout(\quad_counter1.n30504 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_8_lut_LC_23_9_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_8_lut_LC_23_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_8_lut_LC_23_9_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1616_8_lut_LC_23_9_6  (
            .in0(N__93729),
            .in1(N__93728),
            .in2(N__88528),
            .in3(N__88278),
            .lcout(\quad_counter1.n2413 ),
            .ltout(),
            .carryin(\quad_counter1.n30504 ),
            .carryout(\quad_counter1.n30505 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_9_lut_LC_23_9_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_9_lut_LC_23_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_9_lut_LC_23_9_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1616_9_lut_LC_23_9_7  (
            .in0(N__93660),
            .in1(N__93656),
            .in2(N__88443),
            .in3(N__88245),
            .lcout(\quad_counter1.n2412 ),
            .ltout(),
            .carryin(\quad_counter1.n30505 ),
            .carryout(\quad_counter1.n30506 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_10_lut_LC_23_10_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_10_lut_LC_23_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_10_lut_LC_23_10_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1616_10_lut_LC_23_10_0  (
            .in0(N__93933),
            .in1(N__93932),
            .in2(N__88432),
            .in3(N__88215),
            .lcout(\quad_counter1.n2411 ),
            .ltout(),
            .carryin(bfn_23_10_0_),
            .carryout(\quad_counter1.n30507 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_11_lut_LC_23_10_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_11_lut_LC_23_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_11_lut_LC_23_10_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1616_11_lut_LC_23_10_1  (
            .in0(N__93621),
            .in1(N__93620),
            .in2(N__88440),
            .in3(N__88182),
            .lcout(\quad_counter1.n2410 ),
            .ltout(),
            .carryin(\quad_counter1.n30507 ),
            .carryout(\quad_counter1.n30508 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_12_lut_LC_23_10_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1616_12_lut_LC_23_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_12_lut_LC_23_10_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1616_12_lut_LC_23_10_2  (
            .in0(N__93591),
            .in1(N__93590),
            .in2(N__88433),
            .in3(N__88155),
            .lcout(\quad_counter1.n2409 ),
            .ltout(),
            .carryin(\quad_counter1.n30508 ),
            .carryout(\quad_counter1.n30509 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1616_13_lut_LC_23_10_3 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1616_13_lut_LC_23_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1616_13_lut_LC_23_10_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1616_13_lut_LC_23_10_3  (
            .in0(N__93956),
            .in1(N__93957),
            .in2(N__88441),
            .in3(N__88152),
            .lcout(\quad_counter1.n2408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_9_i3_2_lut_LC_23_10_5 .C_ON=1'b0;
    defparam \c0.select_369_Select_9_i3_2_lut_LC_23_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_9_i3_2_lut_LC_23_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_9_i3_2_lut_LC_23_10_5  (
            .in0(N__91736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94821),
            .lcout(\c0.n3_adj_4588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_3_lut_adj_1269_LC_23_10_6 .C_ON=1'b0;
    defparam \quad_counter1.i1_3_lut_adj_1269_LC_23_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_3_lut_adj_1269_LC_23_10_6 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \quad_counter1.i1_3_lut_adj_1269_LC_23_10_6  (
            .in0(_gnd_net_),
            .in1(N__88122),
            .in2(N__88093),
            .in3(N__88061),
            .lcout(\quad_counter1.n7_adj_4445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30708_1_lut_LC_23_10_7 .C_ON=1'b0;
    defparam \quad_counter1.i30708_1_lut_LC_23_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30708_1_lut_LC_23_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \quad_counter1.i30708_1_lut_LC_23_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__88414),
            .lcout(\quad_counter1.n36135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i10_4_lut_adj_1292_LC_23_11_0 .C_ON=1'b0;
    defparam \quad_counter1.i10_4_lut_adj_1292_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i10_4_lut_adj_1292_LC_23_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i10_4_lut_adj_1292_LC_23_11_0  (
            .in0(N__88632),
            .in1(N__88725),
            .in2(N__88623),
            .in3(N__88890),
            .lcout(\quad_counter1.n28_adj_4460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23561_2_lut_LC_23_11_1 .C_ON=1'b0;
    defparam \quad_counter1.i23561_2_lut_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23561_2_lut_LC_23_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23561_2_lut_LC_23_11_1  (
            .in0(_gnd_net_),
            .in1(N__88482),
            .in2(_gnd_net_),
            .in3(N__93463),
            .lcout(),
            .ltout(\quad_counter1.n28277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1260_LC_23_11_2 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1260_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1260_LC_23_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1260_LC_23_11_2  (
            .in0(N__93439),
            .in1(N__93400),
            .in2(N__88452),
            .in3(N__93721),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_4_lut_LC_23_11_3 .C_ON=1'b0;
    defparam \quad_counter1.i1_4_lut_LC_23_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_4_lut_LC_23_11_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i1_4_lut_LC_23_11_3  (
            .in0(N__93775),
            .in1(N__93649),
            .in2(N__88449),
            .in3(N__93748),
            .lcout(),
            .ltout(\quad_counter1.n7_adj_4439_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1262_LC_23_11_4 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1262_LC_23_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1262_LC_23_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1262_LC_23_11_4  (
            .in0(N__93589),
            .in1(N__93619),
            .in2(N__88446),
            .in3(N__93909),
            .lcout(\quad_counter1.n2342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_2_lut_LC_23_12_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_2_lut_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_2_lut_LC_23_12_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2353_2_lut_LC_23_12_0  (
            .in0(N__88392),
            .in1(N__88391),
            .in2(N__89449),
            .in3(N__88356),
            .lcout(\quad_counter1.n3519 ),
            .ltout(),
            .carryin(bfn_23_12_0_),
            .carryout(\quad_counter1.n30675 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_3_lut_LC_23_12_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_3_lut_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_3_lut_LC_23_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_3_lut_LC_23_12_1  (
            .in0(N__88352),
            .in1(N__88351),
            .in2(N__89568),
            .in3(N__88332),
            .lcout(\quad_counter1.n3518 ),
            .ltout(),
            .carryin(\quad_counter1.n30675 ),
            .carryout(\quad_counter1.n30676 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_4_lut_LC_23_12_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_4_lut_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_4_lut_LC_23_12_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2353_4_lut_LC_23_12_2  (
            .in0(N__88329),
            .in1(N__88328),
            .in2(N__89450),
            .in3(N__88311),
            .lcout(\quad_counter1.n3517 ),
            .ltout(),
            .carryin(\quad_counter1.n30676 ),
            .carryout(\quad_counter1.n30677 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_5_lut_LC_23_12_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_5_lut_LC_23_12_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_5_lut_LC_23_12_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2353_5_lut_LC_23_12_3  (
            .in0(N__88716),
            .in1(N__88715),
            .in2(N__89453),
            .in3(N__88698),
            .lcout(\quad_counter1.n3516 ),
            .ltout(),
            .carryin(\quad_counter1.n30677 ),
            .carryout(\quad_counter1.n30678 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_6_lut_LC_23_12_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_6_lut_LC_23_12_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_6_lut_LC_23_12_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2353_6_lut_LC_23_12_4  (
            .in0(N__88695),
            .in1(N__88694),
            .in2(N__89451),
            .in3(N__88674),
            .lcout(\quad_counter1.n3515 ),
            .ltout(),
            .carryin(\quad_counter1.n30678 ),
            .carryout(\quad_counter1.n30679 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_7_lut_LC_23_12_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_7_lut_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_7_lut_LC_23_12_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2353_7_lut_LC_23_12_5  (
            .in0(N__88671),
            .in1(N__88670),
            .in2(N__89454),
            .in3(N__88653),
            .lcout(\quad_counter1.n3514 ),
            .ltout(),
            .carryin(\quad_counter1.n30679 ),
            .carryout(\quad_counter1.n30680 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_8_lut_LC_23_12_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_8_lut_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_8_lut_LC_23_12_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_2353_8_lut_LC_23_12_6  (
            .in0(N__88650),
            .in1(N__88649),
            .in2(N__89452),
            .in3(N__88626),
            .lcout(\quad_counter1.n3513 ),
            .ltout(),
            .carryin(\quad_counter1.n30680 ),
            .carryout(\quad_counter1.n30681 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_9_lut_LC_23_12_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_9_lut_LC_23_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_9_lut_LC_23_12_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_9_lut_LC_23_12_7  (
            .in0(N__88958),
            .in1(N__88957),
            .in2(N__89569),
            .in3(N__88614),
            .lcout(\quad_counter1.n3512 ),
            .ltout(),
            .carryin(\quad_counter1.n30681 ),
            .carryout(\quad_counter1.n30682 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_10_lut_LC_23_13_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_10_lut_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_10_lut_LC_23_13_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_10_lut_LC_23_13_0  (
            .in0(N__88607),
            .in1(N__88606),
            .in2(N__89570),
            .in3(N__88587),
            .lcout(\quad_counter1.n3511 ),
            .ltout(),
            .carryin(bfn_23_13_0_),
            .carryout(\quad_counter1.n30683 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_11_lut_LC_23_13_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_11_lut_LC_23_13_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_11_lut_LC_23_13_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_11_lut_LC_23_13_1  (
            .in0(N__88982),
            .in1(N__88981),
            .in2(N__89574),
            .in3(N__88572),
            .lcout(\quad_counter1.n3510 ),
            .ltout(),
            .carryin(\quad_counter1.n30683 ),
            .carryout(\quad_counter1.n30684 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_12_lut_LC_23_13_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_12_lut_LC_23_13_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_12_lut_LC_23_13_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_12_lut_LC_23_13_2  (
            .in0(N__88569),
            .in1(N__88568),
            .in2(N__89571),
            .in3(N__88551),
            .lcout(\quad_counter1.n3509 ),
            .ltout(),
            .carryin(\quad_counter1.n30684 ),
            .carryout(\quad_counter1.n30685 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_13_lut_LC_23_13_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_13_lut_LC_23_13_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_13_lut_LC_23_13_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_13_lut_LC_23_13_3  (
            .in0(N__88548),
            .in1(N__88547),
            .in2(N__89575),
            .in3(N__88914),
            .lcout(\quad_counter1.n3508 ),
            .ltout(),
            .carryin(\quad_counter1.n30685 ),
            .carryout(\quad_counter1.n30686 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_14_lut_LC_23_13_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_14_lut_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_14_lut_LC_23_13_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_14_lut_LC_23_13_4  (
            .in0(N__88910),
            .in1(N__88911),
            .in2(N__89572),
            .in3(N__88881),
            .lcout(\quad_counter1.n3507 ),
            .ltout(),
            .carryin(\quad_counter1.n30686 ),
            .carryout(\quad_counter1.n30687 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_15_lut_LC_23_13_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_15_lut_LC_23_13_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_15_lut_LC_23_13_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_15_lut_LC_23_13_5  (
            .in0(N__89019),
            .in1(N__89018),
            .in2(N__89576),
            .in3(N__88878),
            .lcout(\quad_counter1.n3506 ),
            .ltout(),
            .carryin(\quad_counter1.n30687 ),
            .carryout(\quad_counter1.n30688 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_16_lut_LC_23_13_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_16_lut_LC_23_13_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_16_lut_LC_23_13_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_16_lut_LC_23_13_6  (
            .in0(N__88874),
            .in1(N__88873),
            .in2(N__89573),
            .in3(N__88854),
            .lcout(\quad_counter1.n3505 ),
            .ltout(),
            .carryin(\quad_counter1.n30688 ),
            .carryout(\quad_counter1.n30689 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_17_lut_LC_23_13_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_17_lut_LC_23_13_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_17_lut_LC_23_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_17_lut_LC_23_13_7  (
            .in0(N__89001),
            .in1(N__89000),
            .in2(N__89577),
            .in3(N__88842),
            .lcout(\quad_counter1.n3504 ),
            .ltout(),
            .carryin(\quad_counter1.n30689 ),
            .carryout(\quad_counter1.n30690 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_18_lut_LC_23_14_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_18_lut_LC_23_14_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_18_lut_LC_23_14_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_18_lut_LC_23_14_0  (
            .in0(N__88839),
            .in1(N__88838),
            .in2(N__89564),
            .in3(N__88809),
            .lcout(\quad_counter1.n3503 ),
            .ltout(),
            .carryin(bfn_23_14_0_),
            .carryout(\quad_counter1.n30691 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_19_lut_LC_23_14_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_19_lut_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_19_lut_LC_23_14_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_19_lut_LC_23_14_1  (
            .in0(N__88806),
            .in1(N__88805),
            .in2(N__89578),
            .in3(N__88779),
            .lcout(\quad_counter1.n3502 ),
            .ltout(),
            .carryin(\quad_counter1.n30691 ),
            .carryout(\quad_counter1.n30692 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_20_lut_LC_23_14_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_20_lut_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_20_lut_LC_23_14_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_20_lut_LC_23_14_2  (
            .in0(N__88775),
            .in1(N__88774),
            .in2(N__89565),
            .in3(N__88746),
            .lcout(\quad_counter1.n3501 ),
            .ltout(),
            .carryin(\quad_counter1.n30692 ),
            .carryout(\quad_counter1.n30693 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_21_lut_LC_23_14_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_21_lut_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_21_lut_LC_23_14_3 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_21_lut_LC_23_14_3  (
            .in0(N__88743),
            .in1(N__88742),
            .in2(N__89579),
            .in3(N__89148),
            .lcout(\quad_counter1.n3500 ),
            .ltout(),
            .carryin(\quad_counter1.n30693 ),
            .carryout(\quad_counter1.n30694 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_22_lut_LC_23_14_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_22_lut_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_22_lut_LC_23_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_22_lut_LC_23_14_4  (
            .in0(N__89144),
            .in1(N__89143),
            .in2(N__89566),
            .in3(N__89115),
            .lcout(\quad_counter1.n3499 ),
            .ltout(),
            .carryin(\quad_counter1.n30694 ),
            .carryout(\quad_counter1.n30695 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_23_lut_LC_23_14_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_2353_23_lut_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_23_lut_LC_23_14_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_23_lut_LC_23_14_5  (
            .in0(N__89112),
            .in1(N__89111),
            .in2(N__89580),
            .in3(N__89085),
            .lcout(\quad_counter1.n3498 ),
            .ltout(),
            .carryin(\quad_counter1.n30695 ),
            .carryout(\quad_counter1.n30696 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_2353_24_lut_LC_23_14_6 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_2353_24_lut_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_2353_24_lut_LC_23_14_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_2353_24_lut_LC_23_14_6  (
            .in0(N__89081),
            .in1(N__89082),
            .in2(N__89567),
            .in3(N__89064),
            .lcout(),
            .ltout(\quad_counter1.n3497_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1295_LC_23_14_7 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1295_LC_23_14_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1295_LC_23_14_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1295_LC_23_14_7  (
            .in0(N__89061),
            .in1(N__89055),
            .in2(N__89049),
            .in3(N__89046),
            .lcout(\quad_counter1.n30_adj_4463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1297_LC_23_15_0 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1297_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1297_LC_23_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1297_LC_23_15_0  (
            .in0(N__89319),
            .in1(N__89343),
            .in2(N__89409),
            .in3(N__89292),
            .lcout(),
            .ltout(\quad_counter1.n12_adj_4464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30568_4_lut_LC_23_15_1 .C_ON=1'b0;
    defparam \quad_counter1.i30568_4_lut_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30568_4_lut_LC_23_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i30568_4_lut_LC_23_15_1  (
            .in0(N__89232),
            .in1(N__89367),
            .in2(N__89031),
            .in3(N__89268),
            .lcout(\quad_counter1.n35985 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i12_4_lut_adj_1249_LC_23_15_4 .C_ON=1'b0;
    defparam \quad_counter1.i12_4_lut_adj_1249_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i12_4_lut_adj_1249_LC_23_15_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i12_4_lut_adj_1249_LC_23_15_4  (
            .in0(N__89017),
            .in1(N__88999),
            .in2(N__88983),
            .in3(N__88962),
            .lcout(),
            .ltout(\quad_counter1.n29_adj_4428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i16_4_lut_LC_23_15_5 .C_ON=1'b0;
    defparam \quad_counter1.i16_4_lut_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i16_4_lut_LC_23_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i16_4_lut_LC_23_15_5  (
            .in0(N__88938),
            .in1(N__88926),
            .in2(N__89589),
            .in3(N__89586),
            .lcout(\quad_counter1.n3431 ),
            .ltout(\quad_counter1.n3431_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30715_1_lut_LC_23_15_6 .C_ON=1'b0;
    defparam \quad_counter1.i30715_1_lut_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30715_1_lut_LC_23_15_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30715_1_lut_LC_23_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__89457),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_15_i3_2_lut_LC_23_16_1 .C_ON=1'b0;
    defparam \c0.select_369_Select_15_i3_2_lut_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_15_i3_2_lut_LC_23_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_15_i3_2_lut_LC_23_16_1  (
            .in0(_gnd_net_),
            .in1(N__92048),
            .in2(_gnd_net_),
            .in3(N__94690),
            .lcout(\c0.n3_adj_4594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23692_2_lut_LC_23_16_4 .C_ON=1'b0;
    defparam \quad_counter1.i23692_2_lut_LC_23_16_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23692_2_lut_LC_23_16_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23692_2_lut_LC_23_16_4  (
            .in0(_gnd_net_),
            .in1(N__89402),
            .in2(_gnd_net_),
            .in3(N__89366),
            .lcout(),
            .ltout(\quad_counter1.n28415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1294_LC_23_16_5 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1294_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1294_LC_23_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1294_LC_23_16_5  (
            .in0(N__89342),
            .in1(N__89318),
            .in2(N__89295),
            .in3(N__89291),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4462_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_adj_1296_LC_23_16_6 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_adj_1296_LC_23_16_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_adj_1296_LC_23_16_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i3_4_lut_adj_1296_LC_23_16_6  (
            .in0(N__89267),
            .in1(N__89244),
            .in2(N__89235),
            .in3(N__89231),
            .lcout(\quad_counter1.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_23_16_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_23_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_23_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_23_16_7  (
            .in0(N__89202),
            .in1(N__89184),
            .in2(_gnd_net_),
            .in3(N__96182),
            .lcout(\c0.n11_adj_4513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_6_i3_2_lut_LC_23_17_0 .C_ON=1'b0;
    defparam \c0.select_369_Select_6_i3_2_lut_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_6_i3_2_lut_LC_23_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_6_i3_2_lut_LC_23_17_0  (
            .in0(_gnd_net_),
            .in1(N__91638),
            .in2(_gnd_net_),
            .in3(N__94780),
            .lcout(\c0.n3_adj_4585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1376_LC_23_17_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1376_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1376_LC_23_17_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1376_LC_23_17_1  (
            .in0(N__90408),
            .in1(N__90449),
            .in2(N__94929),
            .in3(N__94422),
            .lcout(\c0.n33607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_8_i3_2_lut_LC_23_17_2 .C_ON=1'b0;
    defparam \c0.select_369_Select_8_i3_2_lut_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_8_i3_2_lut_LC_23_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_8_i3_2_lut_LC_23_17_2  (
            .in0(N__91785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94781),
            .lcout(\c0.n3_adj_4587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_4_lut_LC_23_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_4_lut_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_4_lut_LC_23_17_3 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_4_lut_LC_23_17_3  (
            .in0(N__101204),
            .in1(N__101295),
            .in2(N__98043),
            .in3(N__100683),
            .lcout(\c0.n32377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_11_i3_2_lut_LC_23_17_4 .C_ON=1'b0;
    defparam \c0.select_369_Select_11_i3_2_lut_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_11_i3_2_lut_LC_23_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_11_i3_2_lut_LC_23_17_4  (
            .in0(_gnd_net_),
            .in1(N__91887),
            .in2(_gnd_net_),
            .in3(N__94782),
            .lcout(\c0.n3_adj_4590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1403_LC_23_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1403_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1403_LC_23_17_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1403_LC_23_17_5  (
            .in0(N__101203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__101294),
            .lcout(\c0.n33379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_13_i3_2_lut_LC_23_17_6 .C_ON=1'b0;
    defparam \c0.select_369_Select_13_i3_2_lut_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_13_i3_2_lut_LC_23_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_13_i3_2_lut_LC_23_17_6  (
            .in0(N__91968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94783),
            .lcout(\c0.n3_adj_4592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_23_17_7 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_23_17_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_LC_23_17_7  (
            .in0(N__91528),
            .in1(N__92322),
            .in2(N__92127),
            .in3(N__91784),
            .lcout(\c0.n45_adj_4645 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_23_18_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_23_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_LC_23_18_0  (
            .in0(N__90429),
            .in1(N__94389),
            .in2(N__90453),
            .in3(N__90602),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.equal_69_i9_2_lut_3_lut_LC_23_18_3 .C_ON=1'b0;
    defparam \c0.equal_69_i9_2_lut_3_lut_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.equal_69_i9_2_lut_3_lut_LC_23_18_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \c0.equal_69_i9_2_lut_3_lut_LC_23_18_3  (
            .in0(N__93223),
            .in1(N__91221),
            .in2(_gnd_net_),
            .in3(N__91097),
            .lcout(\c0.n9_adj_4552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_14_i3_2_lut_LC_23_18_5 .C_ON=1'b0;
    defparam \c0.select_369_Select_14_i3_2_lut_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_14_i3_2_lut_LC_23_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_14_i3_2_lut_LC_23_18_5  (
            .in0(_gnd_net_),
            .in1(N__92009),
            .in2(_gnd_net_),
            .in3(N__94786),
            .lcout(\c0.n3_adj_4593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1920_LC_23_18_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1920_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1920_LC_23_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1920_LC_23_18_6  (
            .in0(N__101342),
            .in1(N__101197),
            .in2(N__100750),
            .in3(N__101089),
            .lcout(\c0.n15827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_12_i3_2_lut_LC_23_18_7 .C_ON=1'b0;
    defparam \c0.select_369_Select_12_i3_2_lut_LC_23_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_12_i3_2_lut_LC_23_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_12_i3_2_lut_LC_23_18_7  (
            .in0(N__91929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94785),
            .lcout(\c0.n3_adj_4591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1944_LC_23_19_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1944_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1944_LC_23_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1944_LC_23_19_0  (
            .in0(N__98409),
            .in1(N__100104),
            .in2(N__94242),
            .in3(N__96270),
            .lcout(\c0.n31299 ),
            .ltout(\c0.n31299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__6__5295_LC_23_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__6__5295_LC_23_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__6__5295_LC_23_19_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.data_out_frame_28__6__5295_LC_23_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__90423),
            .in3(N__97900),
            .lcout(\c0.data_out_frame_28_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97697),
            .ce(N__96929),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1728_LC_23_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1728_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1728_LC_23_19_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1728_LC_23_19_2  (
            .in0(N__94527),
            .in1(N__98345),
            .in2(_gnd_net_),
            .in3(N__100103),
            .lcout(\c0.n32238 ),
            .ltout(\c0.n32238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__5__5296_LC_23_19_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__5__5296_LC_23_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__5__5296_LC_23_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__5__5296_LC_23_19_3  (
            .in0(N__94893),
            .in1(N__93996),
            .in2(N__90399),
            .in3(N__97901),
            .lcout(\c0.data_out_frame_28_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97697),
            .ce(N__96929),
            .sr(_gnd_net_));
    defparam \c0.i9480_2_lut_LC_23_19_5 .C_ON=1'b0;
    defparam \c0.i9480_2_lut_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9480_2_lut_LC_23_19_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.i9480_2_lut_LC_23_19_5  (
            .in0(N__96180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__90392),
            .lcout(),
            .ltout(\c0.n14078_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30620_4_lut_LC_23_19_6 .C_ON=1'b0;
    defparam \c0.i30620_4_lut_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i30620_4_lut_LC_23_19_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \c0.i30620_4_lut_LC_23_19_6  (
            .in0(N__90105),
            .in1(N__89871),
            .in2(N__89847),
            .in3(N__89844),
            .lcout(\c0.n35983 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_1596_LC_23_20_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_1596_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_1596_LC_23_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_adj_1596_LC_23_20_0  (
            .in0(N__91928),
            .in1(N__92194),
            .in2(N__92010),
            .in3(N__91709),
            .lcout(\c0.n43_adj_4641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_1597_LC_23_20_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_1597_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_1597_LC_23_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_1597_LC_23_20_1  (
            .in0(N__91967),
            .in1(N__92493),
            .in2(N__91842),
            .in3(N__92049),
            .lcout(\c0.n40_adj_4643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_23_20_2 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_23_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_LC_23_20_2  (
            .in0(N__92358),
            .in1(N__91886),
            .in2(N__92093),
            .in3(N__92241),
            .lcout(),
            .ltout(\c0.n41_adj_4642_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i24_4_lut_adj_1598_LC_23_20_3 .C_ON=1'b0;
    defparam \c0.i24_4_lut_adj_1598_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i24_4_lut_adj_1598_LC_23_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i24_4_lut_adj_1598_LC_23_20_3  (
            .in0(N__94125),
            .in1(N__90543),
            .in2(N__90534),
            .in3(N__90531),
            .lcout(),
            .ltout(\c0.n50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_adj_1599_LC_23_20_4 .C_ON=1'b0;
    defparam \c0.i25_4_lut_adj_1599_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_adj_1599_LC_23_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i25_4_lut_adj_1599_LC_23_20_4  (
            .in0(N__90525),
            .in1(N__90519),
            .in2(N__90510),
            .in3(N__90507),
            .lcout(\c0.n18083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_20_i3_2_lut_LC_23_20_7 .C_ON=1'b0;
    defparam \c0.select_369_Select_20_i3_2_lut_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_20_i3_2_lut_LC_23_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_20_i3_2_lut_LC_23_20_7  (
            .in0(N__92195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94784),
            .lcout(\c0.n3_adj_4599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_19_i3_2_lut_LC_23_21_0 .C_ON=1'b0;
    defparam \c0.select_369_Select_19_i3_2_lut_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_19_i3_2_lut_LC_23_21_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_19_i3_2_lut_LC_23_21_0  (
            .in0(N__94817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92120),
            .lcout(\c0.n3_adj_4598 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1552_LC_23_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1552_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1552_LC_23_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1552_LC_23_21_2  (
            .in0(N__100166),
            .in1(N__98026),
            .in2(N__101341),
            .in3(N__101189),
            .lcout(\c0.n17669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_16_i3_2_lut_LC_23_21_4 .C_ON=1'b0;
    defparam \c0.select_369_Select_16_i3_2_lut_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_16_i3_2_lut_LC_23_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_16_i3_2_lut_LC_23_21_4  (
            .in0(N__94816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92094),
            .lcout(\c0.n3_adj_4595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1554_LC_23_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1554_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1554_LC_23_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1554_LC_23_21_5  (
            .in0(N__101190),
            .in1(N__95007),
            .in2(N__98038),
            .in3(N__101321),
            .lcout(\c0.n32337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_23_22_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_23_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_23_22_0  (
            .in0(N__93846),
            .in1(N__90585),
            .in2(_gnd_net_),
            .in3(N__96179),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i30673_4_lut_LC_23_22_1.C_ON=1'b0;
    defparam i30673_4_lut_LC_23_22_1.SEQ_MODE=4'b0000;
    defparam i30673_4_lut_LC_23_22_1.LUT_INIT=16'b0101000011001100;
    LogicCell40 i30673_4_lut_LC_23_22_1 (
            .in0(N__90877),
            .in1(N__90807),
            .in2(N__90798),
            .in3(N__90789),
            .lcout(n36102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1348_LC_23_22_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1348_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1348_LC_23_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1348_LC_23_22_2  (
            .in0(N__94882),
            .in1(N__90609),
            .in2(N__98217),
            .in3(N__96459),
            .lcout(),
            .ltout(\c0.n14_adj_4522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1350_LC_23_22_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1350_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1350_LC_23_22_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_4_lut_adj_1350_LC_23_22_3  (
            .in0(N__96783),
            .in1(N__90942),
            .in2(N__90591),
            .in3(N__98136),
            .lcout(),
            .ltout(\c0.n9_adj_4524_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__4__5289_LC_23_22_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__4__5289_LC_23_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__4__5289_LC_23_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_29__4__5289_LC_23_22_4  (
            .in0(N__94059),
            .in1(N__94341),
            .in2(N__90588),
            .in3(N__94266),
            .lcout(\c0.data_out_frame_29_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97748),
            .ce(N__96997),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_18_i3_2_lut_LC_23_23_0 .C_ON=1'b0;
    defparam \c0.select_369_Select_18_i3_2_lut_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_18_i3_2_lut_LC_23_23_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_18_i3_2_lut_LC_23_23_0  (
            .in0(N__94802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92163),
            .lcout(\c0.n3_adj_4597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_24_i3_2_lut_LC_23_23_1 .C_ON=1'b0;
    defparam \c0.select_369_Select_24_i3_2_lut_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_24_i3_2_lut_LC_23_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_24_i3_2_lut_LC_23_23_1  (
            .in0(_gnd_net_),
            .in1(N__94190),
            .in2(_gnd_net_),
            .in3(N__94803),
            .lcout(\c0.n3_adj_4603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_22_i3_2_lut_LC_23_23_2 .C_ON=1'b0;
    defparam \c0.select_369_Select_22_i3_2_lut_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_22_i3_2_lut_LC_23_23_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_22_i3_2_lut_LC_23_23_2  (
            .in0(N__94804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92240),
            .lcout(\c0.n3_adj_4601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1757_LC_23_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1757_LC_23_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1757_LC_23_23_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1757_LC_23_23_4  (
            .in0(N__90941),
            .in1(N__100884),
            .in2(N__100257),
            .in3(N__90579),
            .lcout(\c0.n35251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_1595_LC_23_23_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_1595_LC_23_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_1595_LC_23_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_1595_LC_23_23_5  (
            .in0(N__92162),
            .in1(N__92423),
            .in2(N__91639),
            .in3(N__92272),
            .lcout(\c0.n42_adj_4640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_23_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1742_LC_23_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1742_LC_23_23_6  (
            .in0(N__94371),
            .in1(N__96492),
            .in2(_gnd_net_),
            .in3(N__90940),
            .lcout(\c0.n32359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_2_i3_2_lut_LC_23_23_7 .C_ON=1'b0;
    defparam \c0.select_369_Select_2_i3_2_lut_LC_23_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_2_i3_2_lut_LC_23_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_2_i3_2_lut_LC_23_23_7  (
            .in0(_gnd_net_),
            .in1(N__91239),
            .in2(_gnd_net_),
            .in3(N__94801),
            .lcout(\c0.n3_adj_4580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_29_i3_2_lut_LC_23_24_0 .C_ON=1'b0;
    defparam \c0.select_369_Select_29_i3_2_lut_LC_23_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_29_i3_2_lut_LC_23_24_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_29_i3_2_lut_LC_23_24_0  (
            .in0(N__94814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__92424),
            .lcout(\c0.n3_adj_4608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_23_i3_2_lut_LC_23_24_7 .C_ON=1'b0;
    defparam \c0.select_369_Select_23_i3_2_lut_LC_23_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_23_i3_2_lut_LC_23_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_23_i3_2_lut_LC_23_24_7  (
            .in0(_gnd_net_),
            .in1(N__92274),
            .in2(_gnd_net_),
            .in3(N__94815),
            .lcout(\c0.n3_adj_4602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_25_i3_2_lut_LC_23_26_4 .C_ON=1'b0;
    defparam \c0.select_369_Select_25_i3_2_lut_LC_23_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_25_i3_2_lut_LC_23_26_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.select_369_Select_25_i3_2_lut_LC_23_26_4  (
            .in0(N__94832),
            .in1(N__92318),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n3_adj_4604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_26_i3_2_lut_LC_23_27_2 .C_ON=1'b0;
    defparam \c0.select_369_Select_26_i3_2_lut_LC_23_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_26_i3_2_lut_LC_23_27_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.select_369_Select_26_i3_2_lut_LC_23_27_2  (
            .in0(N__94831),
            .in1(N__92354),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n3_adj_4605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_30_i3_2_lut_LC_23_28_0 .C_ON=1'b0;
    defparam \c0.select_369_Select_30_i3_2_lut_LC_23_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_30_i3_2_lut_LC_23_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_30_i3_2_lut_LC_23_28_0  (
            .in0(_gnd_net_),
            .in1(N__94151),
            .in2(_gnd_net_),
            .in3(N__94748),
            .lcout(\c0.n3_adj_4609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_27_i3_2_lut_LC_23_28_6 .C_ON=1'b0;
    defparam \c0.select_369_Select_27_i3_2_lut_LC_23_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_27_i3_2_lut_LC_23_28_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_27_i3_2_lut_LC_23_28_6  (
            .in0(_gnd_net_),
            .in1(N__92390),
            .in2(_gnd_net_),
            .in3(N__94749),
            .lcout(\c0.n3_adj_4606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i0_LC_24_1_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i0_LC_24_1_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i0_LC_24_1_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_24_1_0  (
            .in0(_gnd_net_),
            .in1(N__93133),
            .in2(N__90912),
            .in3(N__92877),
            .lcout(\c0.FRAME_MATCHER_i_0 ),
            .ltout(),
            .carryin(bfn_24_1_0_),
            .carryout(\c0.n29970 ),
            .clk(N__97540),
            .ce(),
            .sr(N__93117));
    defparam \c0.add_49_2_THRU_CRY_0_LC_24_1_1 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_0_LC_24_1_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_0_LC_24_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_0_LC_24_1_1  (
            .in0(_gnd_net_),
            .in1(N__99188),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970 ),
            .carryout(\c0.n29970_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_1_LC_24_1_2 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_1_LC_24_1_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_1_LC_24_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_1_LC_24_1_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99338),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29970_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_2_LC_24_1_3 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_2_LC_24_1_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_2_LC_24_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_2_LC_24_1_3  (
            .in0(_gnd_net_),
            .in1(N__99192),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29970_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_3_LC_24_1_4 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_3_LC_24_1_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_3_LC_24_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_3_LC_24_1_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99339),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29970_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_4_LC_24_1_5 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_4_LC_24_1_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_4_LC_24_1_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_4_LC_24_1_5  (
            .in0(_gnd_net_),
            .in1(N__99196),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29970_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_5_LC_24_1_6 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_5_LC_24_1_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_5_LC_24_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_5_LC_24_1_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99340),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29970_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_2_THRU_CRY_6_LC_24_1_7 .C_ON=1'b1;
    defparam \c0.add_49_2_THRU_CRY_6_LC_24_1_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_2_THRU_CRY_6_LC_24_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_2_THRU_CRY_6_LC_24_1_7  (
            .in0(_gnd_net_),
            .in1(N__99200),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29970_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29970_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i1_LC_24_2_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i1_LC_24_2_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_24_2_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_24_2_0  (
            .in0(N__92876),
            .in1(N__90981),
            .in2(_gnd_net_),
            .in3(N__90963),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(bfn_24_2_0_),
            .carryout(\c0.n29971 ),
            .clk(N__97543),
            .ce(),
            .sr(N__90960));
    defparam \c0.add_49_3_THRU_CRY_0_LC_24_2_1 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_0_LC_24_2_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_0_LC_24_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_0_LC_24_2_1  (
            .in0(_gnd_net_),
            .in1(N__99175),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971 ),
            .carryout(\c0.n29971_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_1_LC_24_2_2 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_1_LC_24_2_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_1_LC_24_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_1_LC_24_2_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99335),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29971_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_2_LC_24_2_3 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_2_LC_24_2_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_2_LC_24_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_2_LC_24_2_3  (
            .in0(_gnd_net_),
            .in1(N__99179),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29971_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_3_LC_24_2_4 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_3_LC_24_2_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_3_LC_24_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_3_LC_24_2_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99336),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29971_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_4_LC_24_2_5 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_4_LC_24_2_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_4_LC_24_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_4_LC_24_2_5  (
            .in0(_gnd_net_),
            .in1(N__99183),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29971_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_5_LC_24_2_6 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_5_LC_24_2_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_5_LC_24_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_5_LC_24_2_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99337),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29971_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_3_THRU_CRY_6_LC_24_2_7 .C_ON=1'b1;
    defparam \c0.add_49_3_THRU_CRY_6_LC_24_2_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_3_THRU_CRY_6_LC_24_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_3_THRU_CRY_6_LC_24_2_7  (
            .in0(_gnd_net_),
            .in1(N__99187),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29971_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29971_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_24_3_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i2_LC_24_3_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_24_3_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_24_3_0  (
            .in0(N__92916),
            .in1(N__91155),
            .in2(_gnd_net_),
            .in3(N__91137),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(bfn_24_3_0_),
            .carryout(\c0.n29972 ),
            .clk(N__97546),
            .ce(),
            .sr(N__91134));
    defparam \c0.add_49_4_THRU_CRY_0_LC_24_3_1 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_0_LC_24_3_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_0_LC_24_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_0_LC_24_3_1  (
            .in0(_gnd_net_),
            .in1(N__99162),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972 ),
            .carryout(\c0.n29972_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_1_LC_24_3_2 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_1_LC_24_3_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_1_LC_24_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_1_LC_24_3_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99332),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29972_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_2_LC_24_3_3 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_2_LC_24_3_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_2_LC_24_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_2_LC_24_3_3  (
            .in0(_gnd_net_),
            .in1(N__99166),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29972_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_3_LC_24_3_4 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_3_LC_24_3_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_3_LC_24_3_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_3_LC_24_3_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99333),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29972_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_4_LC_24_3_5 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_4_LC_24_3_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_4_LC_24_3_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_4_LC_24_3_5  (
            .in0(_gnd_net_),
            .in1(N__99170),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29972_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_5_LC_24_3_6 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_5_LC_24_3_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_5_LC_24_3_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_5_LC_24_3_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99334),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29972_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_4_THRU_CRY_6_LC_24_3_7 .C_ON=1'b1;
    defparam \c0.add_49_4_THRU_CRY_6_LC_24_3_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_4_THRU_CRY_6_LC_24_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_4_THRU_CRY_6_LC_24_3_7  (
            .in0(_gnd_net_),
            .in1(N__99174),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29972_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29972_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i3_LC_24_4_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i3_LC_24_4_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_24_4_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_24_4_0  (
            .in0(N__92915),
            .in1(N__91294),
            .in2(_gnd_net_),
            .in3(N__91278),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(bfn_24_4_0_),
            .carryout(\c0.n29973 ),
            .clk(N__97551),
            .ce(),
            .sr(N__91275));
    defparam \c0.add_49_5_THRU_CRY_0_LC_24_4_1 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_0_LC_24_4_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_0_LC_24_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_0_LC_24_4_1  (
            .in0(_gnd_net_),
            .in1(N__98949),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973 ),
            .carryout(\c0.n29973_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_1_LC_24_4_2 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_1_LC_24_4_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_1_LC_24_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_1_LC_24_4_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99152),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29973_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_2_LC_24_4_3 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_2_LC_24_4_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_2_LC_24_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_2_LC_24_4_3  (
            .in0(_gnd_net_),
            .in1(N__98953),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29973_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_3_LC_24_4_4 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_3_LC_24_4_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_3_LC_24_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_3_LC_24_4_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99153),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29973_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_4_LC_24_4_5 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_4_LC_24_4_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_4_LC_24_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_4_LC_24_4_5  (
            .in0(_gnd_net_),
            .in1(N__98957),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29973_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_5_LC_24_4_6 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_5_LC_24_4_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_5_LC_24_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_5_LC_24_4_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99154),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29973_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_5_THRU_CRY_6_LC_24_4_7 .C_ON=1'b1;
    defparam \c0.add_49_5_THRU_CRY_6_LC_24_4_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_5_THRU_CRY_6_LC_24_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_5_THRU_CRY_6_LC_24_4_7  (
            .in0(_gnd_net_),
            .in1(N__98961),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29973_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29973_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i4_LC_24_5_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i4_LC_24_5_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_24_5_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_24_5_0  (
            .in0(N__92914),
            .in1(N__91404),
            .in2(_gnd_net_),
            .in3(N__91383),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(bfn_24_5_0_),
            .carryout(\c0.n29974 ),
            .clk(N__97556),
            .ce(),
            .sr(N__91380));
    defparam \c0.add_49_6_THRU_CRY_0_LC_24_5_1 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_0_LC_24_5_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_0_LC_24_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_0_LC_24_5_1  (
            .in0(_gnd_net_),
            .in1(N__98978),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974 ),
            .carryout(\c0.n29974_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_1_LC_24_5_2 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_1_LC_24_5_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_1_LC_24_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_1_LC_24_5_2  (
            .in0(_gnd_net_),
            .in1(N__98938),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29974_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_2_LC_24_5_3 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_2_LC_24_5_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_2_LC_24_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_2_LC_24_5_3  (
            .in0(_gnd_net_),
            .in1(N__98979),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29974_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_3_LC_24_5_4 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_3_LC_24_5_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_3_LC_24_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_3_LC_24_5_4  (
            .in0(_gnd_net_),
            .in1(N__98939),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29974_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_4_LC_24_5_5 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_4_LC_24_5_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_4_LC_24_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_4_LC_24_5_5  (
            .in0(_gnd_net_),
            .in1(N__98980),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29974_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_5_LC_24_5_6 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_5_LC_24_5_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_5_LC_24_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_5_LC_24_5_6  (
            .in0(_gnd_net_),
            .in1(N__98940),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29974_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_6_THRU_CRY_6_LC_24_5_7 .C_ON=1'b1;
    defparam \c0.add_49_6_THRU_CRY_6_LC_24_5_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_6_THRU_CRY_6_LC_24_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_6_THRU_CRY_6_LC_24_5_7  (
            .in0(_gnd_net_),
            .in1(N__98981),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29974_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29974_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_24_6_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i5_LC_24_6_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_24_6_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_24_6_0  (
            .in0(N__92875),
            .in1(N__91501),
            .in2(_gnd_net_),
            .in3(N__91485),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(bfn_24_6_0_),
            .carryout(\c0.n29975 ),
            .clk(N__97559),
            .ce(),
            .sr(N__91482));
    defparam \c0.add_49_7_THRU_CRY_0_LC_24_6_1 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_0_LC_24_6_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_0_LC_24_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_0_LC_24_6_1  (
            .in0(_gnd_net_),
            .in1(N__98925),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975 ),
            .carryout(\c0.n29975_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_1_LC_24_6_2 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_1_LC_24_6_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_1_LC_24_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_1_LC_24_6_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99146),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29975_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_2_LC_24_6_3 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_2_LC_24_6_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_2_LC_24_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_2_LC_24_6_3  (
            .in0(_gnd_net_),
            .in1(N__98929),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29975_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_3_LC_24_6_4 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_3_LC_24_6_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_3_LC_24_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_3_LC_24_6_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99147),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29975_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_4_LC_24_6_5 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_4_LC_24_6_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_4_LC_24_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_4_LC_24_6_5  (
            .in0(_gnd_net_),
            .in1(N__98933),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29975_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_5_LC_24_6_6 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_5_LC_24_6_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_5_LC_24_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_5_LC_24_6_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29975_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_7_THRU_CRY_6_LC_24_6_7 .C_ON=1'b1;
    defparam \c0.add_49_7_THRU_CRY_6_LC_24_6_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_7_THRU_CRY_6_LC_24_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_7_THRU_CRY_6_LC_24_6_7  (
            .in0(_gnd_net_),
            .in1(N__98937),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29975_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29975_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i6_LC_24_7_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i6_LC_24_7_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_24_7_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_24_7_0  (
            .in0(N__92874),
            .in1(N__91591),
            .in2(_gnd_net_),
            .in3(N__91578),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(bfn_24_7_0_),
            .carryout(\c0.n29976 ),
            .clk(N__97566),
            .ce(),
            .sr(N__91575));
    defparam \c0.add_49_8_THRU_CRY_0_LC_24_7_1 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_0_LC_24_7_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_0_LC_24_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_0_LC_24_7_1  (
            .in0(_gnd_net_),
            .in1(N__98749),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976 ),
            .carryout(\c0.n29976_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_1_LC_24_7_2 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_1_LC_24_7_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_1_LC_24_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_1_LC_24_7_2  (
            .in0(_gnd_net_),
            .in1(N__98753),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29976_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_2_LC_24_7_3 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_2_LC_24_7_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_2_LC_24_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_2_LC_24_7_3  (
            .in0(_gnd_net_),
            .in1(N__98750),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29976_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_3_LC_24_7_4 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_3_LC_24_7_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_3_LC_24_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_3_LC_24_7_4  (
            .in0(_gnd_net_),
            .in1(N__98754),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29976_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_4_LC_24_7_5 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_4_LC_24_7_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_4_LC_24_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_4_LC_24_7_5  (
            .in0(_gnd_net_),
            .in1(N__98751),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29976_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_5_LC_24_7_6 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_5_LC_24_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_5_LC_24_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_5_LC_24_7_6  (
            .in0(_gnd_net_),
            .in1(N__98755),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29976_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_8_THRU_CRY_6_LC_24_7_7 .C_ON=1'b1;
    defparam \c0.add_49_8_THRU_CRY_6_LC_24_7_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_8_THRU_CRY_6_LC_24_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_8_THRU_CRY_6_LC_24_7_7  (
            .in0(_gnd_net_),
            .in1(N__98752),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29976_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29976_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i7_LC_24_8_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i7_LC_24_8_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_24_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_24_8_0  (
            .in0(N__92902),
            .in1(N__91693),
            .in2(_gnd_net_),
            .in3(N__91674),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(bfn_24_8_0_),
            .carryout(\c0.n29977 ),
            .clk(N__97575),
            .ce(),
            .sr(N__91671));
    defparam \c0.add_49_9_THRU_CRY_0_LC_24_8_1 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_0_LC_24_8_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_0_LC_24_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_0_LC_24_8_1  (
            .in0(_gnd_net_),
            .in1(N__98620),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977 ),
            .carryout(\c0.n29977_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_1_LC_24_8_2 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_1_LC_24_8_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_1_LC_24_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_1_LC_24_8_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98779),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29977_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_2_LC_24_8_3 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_2_LC_24_8_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_2_LC_24_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_2_LC_24_8_3  (
            .in0(_gnd_net_),
            .in1(N__98624),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29977_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_3_LC_24_8_4 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_3_LC_24_8_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_3_LC_24_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_3_LC_24_8_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98780),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29977_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_4_LC_24_8_5 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_4_LC_24_8_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_4_LC_24_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_4_LC_24_8_5  (
            .in0(_gnd_net_),
            .in1(N__98628),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29977_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_5_LC_24_8_6 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_5_LC_24_8_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_5_LC_24_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_5_LC_24_8_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98781),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29977_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_9_THRU_CRY_6_LC_24_8_7 .C_ON=1'b1;
    defparam \c0.add_49_9_THRU_CRY_6_LC_24_8_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_9_THRU_CRY_6_LC_24_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_9_THRU_CRY_6_LC_24_8_7  (
            .in0(_gnd_net_),
            .in1(N__98632),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29977_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29977_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i8_LC_24_9_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i8_LC_24_9_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_24_9_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_24_9_0  (
            .in0(N__92873),
            .in1(N__91778),
            .in2(_gnd_net_),
            .in3(N__91764),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(bfn_24_9_0_),
            .carryout(\c0.n29978 ),
            .clk(N__97582),
            .ce(),
            .sr(N__91761));
    defparam \c0.add_49_10_THRU_CRY_0_LC_24_9_1 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_0_LC_24_9_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_0_LC_24_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_0_LC_24_9_1  (
            .in0(_gnd_net_),
            .in1(N__98788),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978 ),
            .carryout(\c0.n29978_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_1_LC_24_9_2 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_1_LC_24_9_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_1_LC_24_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_1_LC_24_9_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98972),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29978_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_2_LC_24_9_3 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_2_LC_24_9_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_2_LC_24_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_2_LC_24_9_3  (
            .in0(_gnd_net_),
            .in1(N__98792),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29978_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_3_LC_24_9_4 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_3_LC_24_9_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_3_LC_24_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_3_LC_24_9_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98973),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29978_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_4_LC_24_9_5 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_4_LC_24_9_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_4_LC_24_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_4_LC_24_9_5  (
            .in0(_gnd_net_),
            .in1(N__98796),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29978_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_5_LC_24_9_6 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_5_LC_24_9_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_5_LC_24_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_5_LC_24_9_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98974),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29978_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_10_THRU_CRY_6_LC_24_9_7 .C_ON=1'b1;
    defparam \c0.add_49_10_THRU_CRY_6_LC_24_9_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_10_THRU_CRY_6_LC_24_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_10_THRU_CRY_6_LC_24_9_7  (
            .in0(_gnd_net_),
            .in1(N__98800),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29978_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29978_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i9_LC_24_10_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i9_LC_24_10_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_24_10_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_24_10_0  (
            .in0(N__92894),
            .in1(N__91735),
            .in2(_gnd_net_),
            .in3(N__91716),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(bfn_24_10_0_),
            .carryout(\c0.n29979 ),
            .clk(N__97590),
            .ce(),
            .sr(N__91848));
    defparam \c0.add_49_11_THRU_CRY_0_LC_24_10_1 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_0_LC_24_10_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_0_LC_24_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_0_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(N__98801),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979 ),
            .carryout(\c0.n29979_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_1_LC_24_10_2 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_1_LC_24_10_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_1_LC_24_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_1_LC_24_10_2  (
            .in0(_gnd_net_),
            .in1(N__98805),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29979_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_2_LC_24_10_3 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_2_LC_24_10_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_2_LC_24_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_2_LC_24_10_3  (
            .in0(_gnd_net_),
            .in1(N__98802),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29979_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_3_LC_24_10_4 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_3_LC_24_10_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_3_LC_24_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_3_LC_24_10_4  (
            .in0(_gnd_net_),
            .in1(N__98806),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29979_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_4_LC_24_10_5 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_4_LC_24_10_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_4_LC_24_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_4_LC_24_10_5  (
            .in0(_gnd_net_),
            .in1(N__98803),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29979_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_5_LC_24_10_6 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_5_LC_24_10_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_5_LC_24_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_5_LC_24_10_6  (
            .in0(_gnd_net_),
            .in1(N__98807),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29979_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_11_THRU_CRY_6_LC_24_10_7 .C_ON=1'b1;
    defparam \c0.add_49_11_THRU_CRY_6_LC_24_10_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_11_THRU_CRY_6_LC_24_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_11_THRU_CRY_6_LC_24_10_7  (
            .in0(_gnd_net_),
            .in1(N__98804),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29979_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29979_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i10_LC_24_11_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i10_LC_24_11_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_24_11_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_24_11_0  (
            .in0(N__92844),
            .in1(N__91822),
            .in2(_gnd_net_),
            .in3(N__91803),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(bfn_24_11_0_),
            .carryout(\c0.n29980 ),
            .clk(N__97598),
            .ce(),
            .sr(N__91800));
    defparam \c0.add_49_12_THRU_CRY_0_LC_24_11_1 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_0_LC_24_11_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_0_LC_24_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_0_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(N__98808),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980 ),
            .carryout(\c0.n29980_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_1_LC_24_11_2 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_1_LC_24_11_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_1_LC_24_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_1_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98975),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29980_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_2_LC_24_11_3 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_2_LC_24_11_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_2_LC_24_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_2_LC_24_11_3  (
            .in0(_gnd_net_),
            .in1(N__98812),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29980_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_3_LC_24_11_4 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_3_LC_24_11_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_3_LC_24_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_3_LC_24_11_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29980_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_4_LC_24_11_5 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_4_LC_24_11_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_4_LC_24_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_4_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(N__98816),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29980_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_5_LC_24_11_6 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_5_LC_24_11_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_5_LC_24_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_5_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__98977),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29980_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_12_THRU_CRY_6_LC_24_11_7 .C_ON=1'b1;
    defparam \c0.add_49_12_THRU_CRY_6_LC_24_11_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_12_THRU_CRY_6_LC_24_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_12_THRU_CRY_6_LC_24_11_7  (
            .in0(_gnd_net_),
            .in1(N__98820),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29980_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29980_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i11_LC_24_12_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i11_LC_24_12_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_24_12_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_24_12_0  (
            .in0(N__92904),
            .in1(N__91879),
            .in2(_gnd_net_),
            .in3(N__91863),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(bfn_24_12_0_),
            .carryout(\c0.n29981 ),
            .clk(N__97610),
            .ce(),
            .sr(N__91860));
    defparam \c0.add_49_13_THRU_CRY_0_LC_24_12_1 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_0_LC_24_12_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_0_LC_24_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_0_LC_24_12_1  (
            .in0(_gnd_net_),
            .in1(N__98837),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981 ),
            .carryout(\c0.n29981_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_1_LC_24_12_2 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_1_LC_24_12_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_1_LC_24_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_1_LC_24_12_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99027),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29981_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_2_LC_24_12_3 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_2_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_2_LC_24_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_2_LC_24_12_3  (
            .in0(_gnd_net_),
            .in1(N__98841),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29981_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_3_LC_24_12_4 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_3_LC_24_12_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_3_LC_24_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_3_LC_24_12_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99028),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29981_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_4_LC_24_12_5 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_4_LC_24_12_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_4_LC_24_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_4_LC_24_12_5  (
            .in0(_gnd_net_),
            .in1(N__98845),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29981_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_5_LC_24_12_6 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_5_LC_24_12_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_5_LC_24_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_5_LC_24_12_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99029),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29981_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_13_THRU_CRY_6_LC_24_12_7 .C_ON=1'b1;
    defparam \c0.add_49_13_THRU_CRY_6_LC_24_12_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_13_THRU_CRY_6_LC_24_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_13_THRU_CRY_6_LC_24_12_7  (
            .in0(_gnd_net_),
            .in1(N__98849),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29981_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29981_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_24_13_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i12_LC_24_13_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_24_13_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_24_13_0  (
            .in0(N__92903),
            .in1(N__91913),
            .in2(_gnd_net_),
            .in3(N__91902),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(bfn_24_13_0_),
            .carryout(\c0.n29982 ),
            .clk(N__97622),
            .ce(),
            .sr(N__91899));
    defparam \c0.add_49_14_THRU_CRY_0_LC_24_13_1 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_0_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_0_LC_24_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_0_LC_24_13_1  (
            .in0(_gnd_net_),
            .in1(N__99030),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982 ),
            .carryout(\c0.n29982_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_1_LC_24_13_2 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_1_LC_24_13_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_1_LC_24_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_1_LC_24_13_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99201),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29982_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_2_LC_24_13_3 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_2_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_2_LC_24_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_2_LC_24_13_3  (
            .in0(_gnd_net_),
            .in1(N__99034),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29982_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_3_LC_24_13_4 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_3_LC_24_13_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_3_LC_24_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_3_LC_24_13_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99202),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29982_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_4_LC_24_13_5 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_4_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_4_LC_24_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_4_LC_24_13_5  (
            .in0(_gnd_net_),
            .in1(N__99038),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29982_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_5_LC_24_13_6 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_5_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_5_LC_24_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_5_LC_24_13_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99203),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29982_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_14_THRU_CRY_6_LC_24_13_7 .C_ON=1'b1;
    defparam \c0.add_49_14_THRU_CRY_6_LC_24_13_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_14_THRU_CRY_6_LC_24_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_14_THRU_CRY_6_LC_24_13_7  (
            .in0(_gnd_net_),
            .in1(N__99042),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29982_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29982_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i13_LC_24_14_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i13_LC_24_14_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_24_14_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_24_14_0  (
            .in0(N__92841),
            .in1(N__91960),
            .in2(_gnd_net_),
            .in3(N__91944),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(bfn_24_14_0_),
            .carryout(\c0.n29983 ),
            .clk(N__97636),
            .ce(),
            .sr(N__91941));
    defparam \c0.add_49_15_THRU_CRY_0_LC_24_14_1 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_0_LC_24_14_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_0_LC_24_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_0_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(N__99043),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983 ),
            .carryout(\c0.n29983_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_1_LC_24_14_2 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_1_LC_24_14_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_1_LC_24_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_1_LC_24_14_2  (
            .in0(_gnd_net_),
            .in1(N__99047),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29983_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_2_LC_24_14_3 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_2_LC_24_14_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_2_LC_24_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_2_LC_24_14_3  (
            .in0(_gnd_net_),
            .in1(N__99044),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29983_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_3_LC_24_14_4 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_3_LC_24_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_3_LC_24_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_3_LC_24_14_4  (
            .in0(_gnd_net_),
            .in1(N__99048),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29983_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_4_LC_24_14_5 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_4_LC_24_14_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_4_LC_24_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_4_LC_24_14_5  (
            .in0(_gnd_net_),
            .in1(N__99045),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29983_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_5_LC_24_14_6 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_5_LC_24_14_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_5_LC_24_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_5_LC_24_14_6  (
            .in0(_gnd_net_),
            .in1(N__99049),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29983_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_15_THRU_CRY_6_LC_24_14_7 .C_ON=1'b1;
    defparam \c0.add_49_15_THRU_CRY_6_LC_24_14_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_15_THRU_CRY_6_LC_24_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_15_THRU_CRY_6_LC_24_14_7  (
            .in0(_gnd_net_),
            .in1(N__99046),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29983_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29983_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i14_LC_24_15_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i14_LC_24_15_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_24_15_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_24_15_0  (
            .in0(N__92839),
            .in1(N__91999),
            .in2(_gnd_net_),
            .in3(N__91983),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(bfn_24_15_0_),
            .carryout(\c0.n29984 ),
            .clk(N__97651),
            .ce(),
            .sr(N__91980));
    defparam \c0.add_49_16_THRU_CRY_0_LC_24_15_1 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_0_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_0_LC_24_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_0_LC_24_15_1  (
            .in0(_gnd_net_),
            .in1(N__99050),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984 ),
            .carryout(\c0.n29984_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_1_LC_24_15_2 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_1_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_1_LC_24_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_1_LC_24_15_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99204),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29984_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_2_LC_24_15_3 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_2_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_2_LC_24_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_2_LC_24_15_3  (
            .in0(_gnd_net_),
            .in1(N__99054),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29984_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_3_LC_24_15_4 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_3_LC_24_15_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_3_LC_24_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_3_LC_24_15_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99205),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29984_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_4_LC_24_15_5 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_4_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_4_LC_24_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_4_LC_24_15_5  (
            .in0(_gnd_net_),
            .in1(N__99058),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29984_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_5_LC_24_15_6 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_5_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_5_LC_24_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_5_LC_24_15_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99206),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29984_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_16_THRU_CRY_6_LC_24_15_7 .C_ON=1'b1;
    defparam \c0.add_49_16_THRU_CRY_6_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_16_THRU_CRY_6_LC_24_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_16_THRU_CRY_6_LC_24_15_7  (
            .in0(_gnd_net_),
            .in1(N__99062),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29984_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29984_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i15_LC_24_16_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i15_LC_24_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_24_16_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_24_16_0  (
            .in0(N__92845),
            .in1(N__92041),
            .in2(_gnd_net_),
            .in3(N__92022),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(bfn_24_16_0_),
            .carryout(\c0.n29985 ),
            .clk(N__97664),
            .ce(),
            .sr(N__92019));
    defparam \c0.add_49_17_THRU_CRY_0_LC_24_16_1 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_0_LC_24_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_0_LC_24_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_0_LC_24_16_1  (
            .in0(_gnd_net_),
            .in1(N__99066),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985 ),
            .carryout(\c0.n29985_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_1_LC_24_16_2 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_1_LC_24_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_1_LC_24_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_1_LC_24_16_2  (
            .in0(_gnd_net_),
            .in1(N__99063),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29985_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_2_LC_24_16_3 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_2_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_2_LC_24_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_2_LC_24_16_3  (
            .in0(_gnd_net_),
            .in1(N__99067),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29985_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_3_LC_24_16_4 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_3_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_3_LC_24_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_3_LC_24_16_4  (
            .in0(_gnd_net_),
            .in1(N__99064),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29985_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_4_LC_24_16_5 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_4_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_4_LC_24_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_4_LC_24_16_5  (
            .in0(_gnd_net_),
            .in1(N__99068),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29985_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_5_LC_24_16_6 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_5_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_5_LC_24_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_5_LC_24_16_6  (
            .in0(_gnd_net_),
            .in1(N__99065),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29985_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_17_THRU_CRY_6_LC_24_16_7 .C_ON=1'b1;
    defparam \c0.add_49_17_THRU_CRY_6_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_17_THRU_CRY_6_LC_24_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_17_THRU_CRY_6_LC_24_16_7  (
            .in0(_gnd_net_),
            .in1(N__99069),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29985_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29985_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_24_17_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i16_LC_24_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_24_17_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_24_17_0  (
            .in0(N__92840),
            .in1(N__92080),
            .in2(_gnd_net_),
            .in3(N__92064),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(bfn_24_17_0_),
            .carryout(\c0.n29986 ),
            .clk(N__97681),
            .ce(),
            .sr(N__92061));
    defparam \c0.add_49_18_THRU_CRY_0_LC_24_17_1 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_0_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_0_LC_24_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_0_LC_24_17_1  (
            .in0(_gnd_net_),
            .in1(N__99207),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986 ),
            .carryout(\c0.n29986_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_1_LC_24_17_2 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_1_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_1_LC_24_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_1_LC_24_17_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99341),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29986_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_2_LC_24_17_3 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_2_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_2_LC_24_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_2_LC_24_17_3  (
            .in0(_gnd_net_),
            .in1(N__99211),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29986_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_3_LC_24_17_4 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_3_LC_24_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_3_LC_24_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_3_LC_24_17_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99342),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29986_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_4_LC_24_17_5 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_4_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_4_LC_24_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_4_LC_24_17_5  (
            .in0(_gnd_net_),
            .in1(N__99215),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29986_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_5_LC_24_17_6 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_5_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_5_LC_24_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_5_LC_24_17_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29986_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_18_THRU_CRY_6_LC_24_17_7 .C_ON=1'b1;
    defparam \c0.add_49_18_THRU_CRY_6_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_18_THRU_CRY_6_LC_24_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_18_THRU_CRY_6_LC_24_17_7  (
            .in0(_gnd_net_),
            .in1(N__99219),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29986_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29986_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i17_LC_24_18_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i17_LC_24_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_24_18_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_24_18_0  (
            .in0(N__92842),
            .in1(N__94463),
            .in2(_gnd_net_),
            .in3(N__92097),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(bfn_24_18_0_),
            .carryout(\c0.n29987 ),
            .clk(N__97698),
            .ce(),
            .sr(N__94449));
    defparam \c0.add_49_19_THRU_CRY_0_LC_24_18_1 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_0_LC_24_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_0_LC_24_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_0_LC_24_18_1  (
            .in0(_gnd_net_),
            .in1(N__99220),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987 ),
            .carryout(\c0.n29987_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_1_LC_24_18_2 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_1_LC_24_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_1_LC_24_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_1_LC_24_18_2  (
            .in0(_gnd_net_),
            .in1(N__99224),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29987_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_2_LC_24_18_3 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_2_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_2_LC_24_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_2_LC_24_18_3  (
            .in0(_gnd_net_),
            .in1(N__99221),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29987_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_3_LC_24_18_4 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_3_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_3_LC_24_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_3_LC_24_18_4  (
            .in0(_gnd_net_),
            .in1(N__99225),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29987_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_4_LC_24_18_5 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_4_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_4_LC_24_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_4_LC_24_18_5  (
            .in0(_gnd_net_),
            .in1(N__99222),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29987_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_5_LC_24_18_6 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_5_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_5_LC_24_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_5_LC_24_18_6  (
            .in0(_gnd_net_),
            .in1(N__99226),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29987_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_19_THRU_CRY_6_LC_24_18_7 .C_ON=1'b1;
    defparam \c0.add_49_19_THRU_CRY_6_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_19_THRU_CRY_6_LC_24_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_19_THRU_CRY_6_LC_24_18_7  (
            .in0(_gnd_net_),
            .in1(N__99223),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29987_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29987_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_24_19_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i18_LC_24_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_24_19_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_24_19_0  (
            .in0(N__92843),
            .in1(N__92156),
            .in2(_gnd_net_),
            .in3(N__92142),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(bfn_24_19_0_),
            .carryout(\c0.n29988 ),
            .clk(N__97714),
            .ce(),
            .sr(N__92139));
    defparam \c0.add_49_20_THRU_CRY_0_LC_24_19_1 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_0_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_0_LC_24_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_0_LC_24_19_1  (
            .in0(_gnd_net_),
            .in1(N__99227),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988 ),
            .carryout(\c0.n29988_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_1_LC_24_19_2 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_1_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_1_LC_24_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_1_LC_24_19_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99344),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29988_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_2_LC_24_19_3 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_2_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_2_LC_24_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_2_LC_24_19_3  (
            .in0(_gnd_net_),
            .in1(N__99231),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29988_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_3_LC_24_19_4 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_3_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_3_LC_24_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_3_LC_24_19_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99345),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29988_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_4_LC_24_19_5 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_4_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_4_LC_24_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_4_LC_24_19_5  (
            .in0(_gnd_net_),
            .in1(N__99235),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29988_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_5_LC_24_19_6 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_5_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_5_LC_24_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_5_LC_24_19_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99346),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29988_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_20_THRU_CRY_6_LC_24_19_7 .C_ON=1'b1;
    defparam \c0.add_49_20_THRU_CRY_6_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_20_THRU_CRY_6_LC_24_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_20_THRU_CRY_6_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(N__99239),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29988_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29988_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i19_LC_24_20_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i19_LC_24_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_24_20_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_24_20_0  (
            .in0(N__92895),
            .in1(N__92119),
            .in2(_gnd_net_),
            .in3(N__92100),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(bfn_24_20_0_),
            .carryout(\c0.n29989 ),
            .clk(N__97731),
            .ce(),
            .sr(N__92205));
    defparam \c0.add_49_21_THRU_CRY_0_LC_24_20_1 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_0_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_0_LC_24_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_0_LC_24_20_1  (
            .in0(_gnd_net_),
            .in1(N__99240),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989 ),
            .carryout(\c0.n29989_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_1_LC_24_20_2 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_1_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_1_LC_24_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_1_LC_24_20_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99347),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29989_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_2_LC_24_20_3 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_2_LC_24_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_2_LC_24_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_2_LC_24_20_3  (
            .in0(_gnd_net_),
            .in1(N__99244),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29989_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_3_LC_24_20_4 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_3_LC_24_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_3_LC_24_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_3_LC_24_20_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29989_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_4_LC_24_20_5 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_4_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_4_LC_24_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_4_LC_24_20_5  (
            .in0(_gnd_net_),
            .in1(N__99248),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29989_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_5_LC_24_20_6 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_5_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_5_LC_24_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_5_LC_24_20_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99349),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29989_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_21_THRU_CRY_6_LC_24_20_7 .C_ON=1'b1;
    defparam \c0.add_49_21_THRU_CRY_6_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_21_THRU_CRY_6_LC_24_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_21_THRU_CRY_6_LC_24_20_7  (
            .in0(_gnd_net_),
            .in1(N__99252),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29989_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29989_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i20_LC_24_21_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i20_LC_24_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_24_21_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_24_21_0  (
            .in0(N__92897),
            .in1(N__92196),
            .in2(_gnd_net_),
            .in3(N__92181),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(bfn_24_21_0_),
            .carryout(\c0.n29990 ),
            .clk(N__97749),
            .ce(),
            .sr(N__92178));
    defparam \c0.add_49_22_THRU_CRY_0_LC_24_21_1 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_0_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_0_LC_24_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_0_LC_24_21_1  (
            .in0(_gnd_net_),
            .in1(N__99350),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990 ),
            .carryout(\c0.n29990_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_1_LC_24_21_2 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_1_LC_24_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_1_LC_24_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_1_LC_24_21_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99467),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29990_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_2_LC_24_21_3 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_2_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_2_LC_24_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_2_LC_24_21_3  (
            .in0(_gnd_net_),
            .in1(N__99354),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29990_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_3_LC_24_21_4 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_3_LC_24_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_3_LC_24_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_3_LC_24_21_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99468),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29990_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_4_LC_24_21_5 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_4_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_4_LC_24_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_4_LC_24_21_5  (
            .in0(_gnd_net_),
            .in1(N__99358),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29990_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_5_LC_24_21_6 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_5_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_5_LC_24_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_5_LC_24_21_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99469),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29990_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_22_THRU_CRY_6_LC_24_21_7 .C_ON=1'b1;
    defparam \c0.add_49_22_THRU_CRY_6_LC_24_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_22_THRU_CRY_6_LC_24_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_22_THRU_CRY_6_LC_24_21_7  (
            .in0(_gnd_net_),
            .in1(N__99362),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29990_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29990_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i21_LC_24_22_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i21_LC_24_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_24_22_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_24_22_0  (
            .in0(N__92898),
            .in1(N__94855),
            .in2(_gnd_net_),
            .in3(N__92208),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(bfn_24_22_0_),
            .carryout(\c0.n29991 ),
            .clk(N__97766),
            .ce(),
            .sr(N__94587));
    defparam \c0.add_49_23_THRU_CRY_0_LC_24_22_1 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_0_LC_24_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_0_LC_24_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_0_LC_24_22_1  (
            .in0(_gnd_net_),
            .in1(N__99363),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991 ),
            .carryout(\c0.n29991_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_1_LC_24_22_2 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_1_LC_24_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_1_LC_24_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_1_LC_24_22_2  (
            .in0(_gnd_net_),
            .in1(N__99367),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29991_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_2_LC_24_22_3 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_2_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_2_LC_24_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_2_LC_24_22_3  (
            .in0(_gnd_net_),
            .in1(N__99364),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29991_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_3_LC_24_22_4 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_3_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_3_LC_24_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_3_LC_24_22_4  (
            .in0(_gnd_net_),
            .in1(N__99368),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29991_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_4_LC_24_22_5 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_4_LC_24_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_4_LC_24_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_4_LC_24_22_5  (
            .in0(_gnd_net_),
            .in1(N__99365),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29991_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_5_LC_24_22_6 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_5_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_5_LC_24_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_5_LC_24_22_6  (
            .in0(_gnd_net_),
            .in1(N__99369),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29991_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_23_THRU_CRY_6_LC_24_22_7 .C_ON=1'b1;
    defparam \c0.add_49_23_THRU_CRY_6_LC_24_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_23_THRU_CRY_6_LC_24_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_23_THRU_CRY_6_LC_24_22_7  (
            .in0(_gnd_net_),
            .in1(N__99366),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29991_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29991_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i22_LC_24_23_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i22_LC_24_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_24_23_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_24_23_0  (
            .in0(N__92899),
            .in1(N__92239),
            .in2(_gnd_net_),
            .in3(N__92220),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(bfn_24_23_0_),
            .carryout(\c0.n29992 ),
            .clk(N__97781),
            .ce(),
            .sr(N__92217));
    defparam \c0.add_49_24_THRU_CRY_0_LC_24_23_1 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_0_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_0_LC_24_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_0_LC_24_23_1  (
            .in0(_gnd_net_),
            .in1(N__99370),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992 ),
            .carryout(\c0.n29992_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_1_LC_24_23_2 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_1_LC_24_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_1_LC_24_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_1_LC_24_23_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99470),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29992_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_2_LC_24_23_3 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_2_LC_24_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_2_LC_24_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_2_LC_24_23_3  (
            .in0(_gnd_net_),
            .in1(N__99374),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29992_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_3_LC_24_23_4 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_3_LC_24_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_3_LC_24_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_3_LC_24_23_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29992_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_4_LC_24_23_5 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_4_LC_24_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_4_LC_24_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_4_LC_24_23_5  (
            .in0(_gnd_net_),
            .in1(N__99378),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29992_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_5_LC_24_23_6 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_5_LC_24_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_5_LC_24_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_5_LC_24_23_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99472),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29992_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_24_THRU_CRY_6_LC_24_23_7 .C_ON=1'b1;
    defparam \c0.add_49_24_THRU_CRY_6_LC_24_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_24_THRU_CRY_6_LC_24_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_24_THRU_CRY_6_LC_24_23_7  (
            .in0(_gnd_net_),
            .in1(N__99382),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29992_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29992_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i23_LC_24_24_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i23_LC_24_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_24_24_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_24_24_0  (
            .in0(N__92900),
            .in1(N__92273),
            .in2(_gnd_net_),
            .in3(N__92256),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(bfn_24_24_0_),
            .carryout(\c0.n29993 ),
            .clk(N__97791),
            .ce(),
            .sr(N__92253));
    defparam \c0.add_49_25_THRU_CRY_0_LC_24_24_1 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_0_LC_24_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_0_LC_24_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_0_LC_24_24_1  (
            .in0(_gnd_net_),
            .in1(N__99383),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993 ),
            .carryout(\c0.n29993_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_1_LC_24_24_2 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_1_LC_24_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_1_LC_24_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_1_LC_24_24_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99473),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29993_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_2_LC_24_24_3 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_2_LC_24_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_2_LC_24_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_2_LC_24_24_3  (
            .in0(_gnd_net_),
            .in1(N__99387),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29993_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_3_LC_24_24_4 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_3_LC_24_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_3_LC_24_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_3_LC_24_24_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99474),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29993_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_4_LC_24_24_5 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_4_LC_24_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_4_LC_24_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_4_LC_24_24_5  (
            .in0(_gnd_net_),
            .in1(N__99391),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29993_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_5_LC_24_24_6 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_5_LC_24_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_5_LC_24_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_5_LC_24_24_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99475),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29993_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_25_THRU_CRY_6_LC_24_24_7 .C_ON=1'b1;
    defparam \c0.add_49_25_THRU_CRY_6_LC_24_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_25_THRU_CRY_6_LC_24_24_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_25_THRU_CRY_6_LC_24_24_7  (
            .in0(_gnd_net_),
            .in1(N__99395),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29993_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29993_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i24_LC_24_25_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i24_LC_24_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_24_25_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_24_25_0  (
            .in0(N__92896),
            .in1(N__94177),
            .in2(_gnd_net_),
            .in3(N__92289),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(bfn_24_25_0_),
            .carryout(\c0.n29994 ),
            .clk(N__97794),
            .ce(),
            .sr(N__92286));
    defparam \c0.add_49_26_THRU_CRY_0_LC_24_25_1 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_0_LC_24_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_0_LC_24_25_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_0_LC_24_25_1  (
            .in0(_gnd_net_),
            .in1(N__99476),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994 ),
            .carryout(\c0.n29994_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_1_LC_24_25_2 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_1_LC_24_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_1_LC_24_25_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_1_LC_24_25_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99562),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29994_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_2_LC_24_25_3 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_2_LC_24_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_2_LC_24_25_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_2_LC_24_25_3  (
            .in0(_gnd_net_),
            .in1(N__99480),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29994_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_3_LC_24_25_4 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_3_LC_24_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_3_LC_24_25_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_3_LC_24_25_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99563),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29994_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_4_LC_24_25_5 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_4_LC_24_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_4_LC_24_25_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_4_LC_24_25_5  (
            .in0(_gnd_net_),
            .in1(N__99484),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29994_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_5_LC_24_25_6 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_5_LC_24_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_5_LC_24_25_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_5_LC_24_25_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29994_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_26_THRU_CRY_6_LC_24_25_7 .C_ON=1'b1;
    defparam \c0.add_49_26_THRU_CRY_6_LC_24_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_26_THRU_CRY_6_LC_24_25_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_26_THRU_CRY_6_LC_24_25_7  (
            .in0(_gnd_net_),
            .in1(N__99488),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29994_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29994_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_24_26_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i25_LC_24_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_24_26_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_24_26_0  (
            .in0(N__92864),
            .in1(N__92317),
            .in2(_gnd_net_),
            .in3(N__92298),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(bfn_24_26_0_),
            .carryout(\c0.n29995 ),
            .clk(N__97796),
            .ce(),
            .sr(N__92295));
    defparam \c0.add_49_27_THRU_CRY_0_LC_24_26_1 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_0_LC_24_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_0_LC_24_26_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_0_LC_24_26_1  (
            .in0(_gnd_net_),
            .in1(N__99489),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995 ),
            .carryout(\c0.n29995_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_1_LC_24_26_2 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_1_LC_24_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_1_LC_24_26_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_1_LC_24_26_2  (
            .in0(_gnd_net_),
            .in1(N__99493),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29995_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_2_LC_24_26_3 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_2_LC_24_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_2_LC_24_26_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_2_LC_24_26_3  (
            .in0(_gnd_net_),
            .in1(N__99490),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29995_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_3_LC_24_26_4 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_3_LC_24_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_3_LC_24_26_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_3_LC_24_26_4  (
            .in0(_gnd_net_),
            .in1(N__99494),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29995_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_4_LC_24_26_5 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_4_LC_24_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_4_LC_24_26_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_4_LC_24_26_5  (
            .in0(_gnd_net_),
            .in1(N__99491),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29995_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_5_LC_24_26_6 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_5_LC_24_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_5_LC_24_26_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_5_LC_24_26_6  (
            .in0(_gnd_net_),
            .in1(N__99495),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29995_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_27_THRU_CRY_6_LC_24_26_7 .C_ON=1'b1;
    defparam \c0.add_49_27_THRU_CRY_6_LC_24_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_27_THRU_CRY_6_LC_24_26_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_27_THRU_CRY_6_LC_24_26_7  (
            .in0(_gnd_net_),
            .in1(N__99492),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29995_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29995_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i26_LC_24_27_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i26_LC_24_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_24_27_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_24_27_0  (
            .in0(N__92865),
            .in1(N__92353),
            .in2(_gnd_net_),
            .in3(N__92334),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(bfn_24_27_0_),
            .carryout(\c0.n29996 ),
            .clk(N__97797),
            .ce(),
            .sr(N__92331));
    defparam \c0.add_49_28_THRU_CRY_0_LC_24_27_1 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_0_LC_24_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_0_LC_24_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_0_LC_24_27_1  (
            .in0(_gnd_net_),
            .in1(N__99496),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996 ),
            .carryout(\c0.n29996_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_1_LC_24_27_2 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_1_LC_24_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_1_LC_24_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_1_LC_24_27_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99565),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29996_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_2_LC_24_27_3 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_2_LC_24_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_2_LC_24_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_2_LC_24_27_3  (
            .in0(_gnd_net_),
            .in1(N__99500),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29996_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_3_LC_24_27_4 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_3_LC_24_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_3_LC_24_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_3_LC_24_27_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99566),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29996_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_4_LC_24_27_5 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_4_LC_24_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_4_LC_24_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_4_LC_24_27_5  (
            .in0(_gnd_net_),
            .in1(N__99504),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29996_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_5_LC_24_27_6 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_5_LC_24_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_5_LC_24_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_5_LC_24_27_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99567),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29996_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_28_THRU_CRY_6_LC_24_27_7 .C_ON=1'b1;
    defparam \c0.add_49_28_THRU_CRY_6_LC_24_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_28_THRU_CRY_6_LC_24_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_28_THRU_CRY_6_LC_24_27_7  (
            .in0(_gnd_net_),
            .in1(N__99508),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29996_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29996_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i27_LC_24_28_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i27_LC_24_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_24_28_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_24_28_0  (
            .in0(N__92866),
            .in1(N__92389),
            .in2(_gnd_net_),
            .in3(N__92370),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(bfn_24_28_0_),
            .carryout(\c0.n29997 ),
            .clk(N__97801),
            .ce(),
            .sr(N__92367));
    defparam \c0.add_49_29_THRU_CRY_0_LC_24_28_1 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_0_LC_24_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_0_LC_24_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_0_LC_24_28_1  (
            .in0(_gnd_net_),
            .in1(N__99558),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997 ),
            .carryout(\c0.n29997_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_1_LC_24_28_2 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_1_LC_24_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_1_LC_24_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_1_LC_24_28_2  (
            .in0(_gnd_net_),
            .in1(N__99509),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29997_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_2_LC_24_28_3 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_2_LC_24_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_2_LC_24_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_2_LC_24_28_3  (
            .in0(_gnd_net_),
            .in1(N__99559),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29997_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_3_LC_24_28_4 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_3_LC_24_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_3_LC_24_28_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_3_LC_24_28_4  (
            .in0(_gnd_net_),
            .in1(N__99510),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29997_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_4_LC_24_28_5 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_4_LC_24_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_4_LC_24_28_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_4_LC_24_28_5  (
            .in0(_gnd_net_),
            .in1(N__99560),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29997_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_5_LC_24_28_6 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_5_LC_24_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_5_LC_24_28_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_5_LC_24_28_6  (
            .in0(_gnd_net_),
            .in1(N__99511),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29997_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_29_THRU_CRY_6_LC_24_28_7 .C_ON=1'b1;
    defparam \c0.add_49_29_THRU_CRY_6_LC_24_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_29_THRU_CRY_6_LC_24_28_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_29_THRU_CRY_6_LC_24_28_7  (
            .in0(_gnd_net_),
            .in1(N__99561),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29997_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29997_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i28_LC_24_29_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i28_LC_24_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_24_29_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_24_29_0  (
            .in0(N__92901),
            .in1(N__92482),
            .in2(_gnd_net_),
            .in3(N__92427),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(bfn_24_29_0_),
            .carryout(\c0.n29998 ),
            .clk(N__97802),
            .ce(),
            .sr(N__92463));
    defparam \c0.add_49_30_THRU_CRY_0_LC_24_29_1 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_0_LC_24_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_0_LC_24_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_0_LC_24_29_1  (
            .in0(_gnd_net_),
            .in1(N__99568),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998 ),
            .carryout(\c0.n29998_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_1_LC_24_29_2 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_1_LC_24_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_1_LC_24_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_1_LC_24_29_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99601),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29998_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_2_LC_24_29_3 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_2_LC_24_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_2_LC_24_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_2_LC_24_29_3  (
            .in0(_gnd_net_),
            .in1(N__99572),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29998_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_3_LC_24_29_4 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_3_LC_24_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_3_LC_24_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_3_LC_24_29_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99602),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29998_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_4_LC_24_29_5 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_4_LC_24_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_4_LC_24_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_4_LC_24_29_5  (
            .in0(_gnd_net_),
            .in1(N__99576),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29998_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_5_LC_24_29_6 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_5_LC_24_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_5_LC_24_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_5_LC_24_29_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99603),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29998_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_30_THRU_CRY_6_LC_24_29_7 .C_ON=1'b1;
    defparam \c0.add_49_30_THRU_CRY_6_LC_24_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_30_THRU_CRY_6_LC_24_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_30_THRU_CRY_6_LC_24_29_7  (
            .in0(_gnd_net_),
            .in1(N__99580),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29998_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29998_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i29_LC_24_30_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i29_LC_24_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_24_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_24_30_0  (
            .in0(N__92870),
            .in1(N__92416),
            .in2(_gnd_net_),
            .in3(N__92400),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(bfn_24_30_0_),
            .carryout(\c0.n29999 ),
            .clk(N__97803),
            .ce(),
            .sr(N__92454));
    defparam \c0.add_49_31_THRU_CRY_0_LC_24_30_1 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_0_LC_24_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_0_LC_24_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_0_LC_24_30_1  (
            .in0(_gnd_net_),
            .in1(N__99581),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999 ),
            .carryout(\c0.n29999_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_1_LC_24_30_2 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_1_LC_24_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_1_LC_24_30_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_1_LC_24_30_2  (
            .in0(_gnd_net_),
            .in1(N__99585),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n29999_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_2_LC_24_30_3 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_2_LC_24_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_2_LC_24_30_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_2_LC_24_30_3  (
            .in0(_gnd_net_),
            .in1(N__99582),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n29999_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_3_LC_24_30_4 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_3_LC_24_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_3_LC_24_30_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_3_LC_24_30_4  (
            .in0(_gnd_net_),
            .in1(N__99586),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n29999_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_4_LC_24_30_5 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_4_LC_24_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_4_LC_24_30_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_4_LC_24_30_5  (
            .in0(_gnd_net_),
            .in1(N__99583),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n29999_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_5_LC_24_30_6 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_5_LC_24_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_5_LC_24_30_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_5_LC_24_30_6  (
            .in0(_gnd_net_),
            .in1(N__99587),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n29999_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_31_THRU_CRY_6_LC_24_30_7 .C_ON=1'b1;
    defparam \c0.add_49_31_THRU_CRY_6_LC_24_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_31_THRU_CRY_6_LC_24_30_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_31_THRU_CRY_6_LC_24_30_7  (
            .in0(_gnd_net_),
            .in1(N__99584),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n29999_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n29999_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i30_LC_24_31_0 .C_ON=1'b1;
    defparam \c0.FRAME_MATCHER_i_i30_LC_24_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_24_31_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_24_31_0  (
            .in0(N__92871),
            .in1(N__94144),
            .in2(_gnd_net_),
            .in3(N__92442),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(bfn_24_31_0_),
            .carryout(\c0.n30000 ),
            .clk(N__97804),
            .ce(),
            .sr(N__92439));
    defparam \c0.add_49_32_THRU_CRY_0_LC_24_31_1 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_0_LC_24_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_0_LC_24_31_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_0_LC_24_31_1  (
            .in0(_gnd_net_),
            .in1(N__99588),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000 ),
            .carryout(\c0.n30000_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_1_LC_24_31_2 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_1_LC_24_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_1_LC_24_31_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_1_LC_24_31_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99604),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000_THRU_CRY_0_THRU_CO ),
            .carryout(\c0.n30000_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_2_LC_24_31_3 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_2_LC_24_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_2_LC_24_31_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_2_LC_24_31_3  (
            .in0(_gnd_net_),
            .in1(N__99592),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000_THRU_CRY_1_THRU_CO ),
            .carryout(\c0.n30000_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_3_LC_24_31_4 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_3_LC_24_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_3_LC_24_31_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_3_LC_24_31_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99605),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000_THRU_CRY_2_THRU_CO ),
            .carryout(\c0.n30000_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_4_LC_24_31_5 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_4_LC_24_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_4_LC_24_31_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_4_LC_24_31_5  (
            .in0(_gnd_net_),
            .in1(N__99596),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000_THRU_CRY_3_THRU_CO ),
            .carryout(\c0.n30000_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_5_LC_24_31_6 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_5_LC_24_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_5_LC_24_31_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_5_LC_24_31_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__99606),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000_THRU_CRY_4_THRU_CO ),
            .carryout(\c0.n30000_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_49_32_THRU_CRY_6_LC_24_31_7 .C_ON=1'b1;
    defparam \c0.add_49_32_THRU_CRY_6_LC_24_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_49_32_THRU_CRY_6_LC_24_31_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \c0.add_49_32_THRU_CRY_6_LC_24_31_7  (
            .in0(_gnd_net_),
            .in1(N__99600),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\c0.n30000_THRU_CRY_5_THRU_CO ),
            .carryout(\c0.n30000_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i31_LC_24_32_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_24_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_24_32_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_24_32_0  (
            .in0(N__92524),
            .in1(N__92872),
            .in2(_gnd_net_),
            .in3(N__92625),
            .lcout(\c0.FRAME_MATCHER_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97805),
            .ce(),
            .sr(N__92505));
    defparam \c0.select_369_Select_31_i3_2_lut_LC_24_32_1 .C_ON=1'b0;
    defparam \c0.select_369_Select_31_i3_2_lut_LC_24_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_31_i3_2_lut_LC_24_32_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_31_i3_2_lut_LC_24_32_1  (
            .in0(_gnd_net_),
            .in1(N__94835),
            .in2(_gnd_net_),
            .in3(N__92523),
            .lcout(\c0.n3_adj_4610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_28_i3_2_lut_LC_24_32_4 .C_ON=1'b0;
    defparam \c0.select_369_Select_28_i3_2_lut_LC_24_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_28_i3_2_lut_LC_24_32_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.select_369_Select_28_i3_2_lut_LC_24_32_4  (
            .in0(N__94836),
            .in1(N__92489),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n3_adj_4607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1251_LC_26_7_2 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1251_LC_26_7_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1251_LC_26_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1251_LC_26_7_2  (
            .in0(N__93379),
            .in1(N__92983),
            .in2(N__92952),
            .in3(N__93022),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1252_LC_26_7_3 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1252_LC_26_7_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1252_LC_26_7_3 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1252_LC_26_7_3  (
            .in0(N__93064),
            .in1(N__93340),
            .in2(N__93240),
            .in3(N__93103),
            .lcout(\quad_counter1.n1847 ),
            .ltout(\quad_counter1.n1847_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30711_1_lut_LC_26_7_4 .C_ON=1'b0;
    defparam \quad_counter1.i30711_1_lut_LC_26_7_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30711_1_lut_LC_26_7_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30711_1_lut_LC_26_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__93237),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_0_i3_2_lut_LC_26_7_6 .C_ON=1'b0;
    defparam \c0.select_369_Select_0_i3_2_lut_LC_26_7_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_0_i3_2_lut_LC_26_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.select_369_Select_0_i3_2_lut_LC_26_7_6  (
            .in0(_gnd_net_),
            .in1(N__93219),
            .in2(_gnd_net_),
            .in3(N__94834),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_2_lut_LC_26_8_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1281_2_lut_LC_26_8_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_2_lut_LC_26_8_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1281_2_lut_LC_26_8_0  (
            .in0(N__93105),
            .in1(N__93104),
            .in2(N__93301),
            .in3(N__93069),
            .lcout(\quad_counter1.n1919 ),
            .ltout(),
            .carryin(bfn_26_8_0_),
            .carryout(\quad_counter1.n30459 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_3_lut_LC_26_8_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1281_3_lut_LC_26_8_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_3_lut_LC_26_8_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1281_3_lut_LC_26_8_1  (
            .in0(N__93066),
            .in1(N__93065),
            .in2(N__93036),
            .in3(N__93027),
            .lcout(\quad_counter1.n1918 ),
            .ltout(),
            .carryin(\quad_counter1.n30459 ),
            .carryout(\quad_counter1.n30460 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_4_lut_LC_26_8_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1281_4_lut_LC_26_8_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_4_lut_LC_26_8_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1281_4_lut_LC_26_8_2  (
            .in0(N__93024),
            .in1(N__93023),
            .in2(N__93302),
            .in3(N__92988),
            .lcout(\quad_counter1.n1917 ),
            .ltout(),
            .carryin(\quad_counter1.n30460 ),
            .carryout(\quad_counter1.n30461 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_5_lut_LC_26_8_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1281_5_lut_LC_26_8_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_5_lut_LC_26_8_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1281_5_lut_LC_26_8_3  (
            .in0(N__92985),
            .in1(N__92984),
            .in2(N__93305),
            .in3(N__92955),
            .lcout(\quad_counter1.n1916 ),
            .ltout(),
            .carryin(\quad_counter1.n30461 ),
            .carryout(\quad_counter1.n30462 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_6_lut_LC_26_8_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1281_6_lut_LC_26_8_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_6_lut_LC_26_8_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1281_6_lut_LC_26_8_4  (
            .in0(N__92951),
            .in1(N__92950),
            .in2(N__93303),
            .in3(N__92919),
            .lcout(\quad_counter1.n1915 ),
            .ltout(),
            .carryin(\quad_counter1.n30462 ),
            .carryout(\quad_counter1.n30463 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_7_lut_LC_26_8_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1281_7_lut_LC_26_8_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_7_lut_LC_26_8_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1281_7_lut_LC_26_8_5  (
            .in0(N__93380),
            .in1(N__93381),
            .in2(N__93306),
            .in3(N__93345),
            .lcout(\quad_counter1.n1914 ),
            .ltout(),
            .carryin(\quad_counter1.n30463 ),
            .carryout(\quad_counter1.n30464 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1281_8_lut_LC_26_8_6 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1281_8_lut_LC_26_8_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1281_8_lut_LC_26_8_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1281_8_lut_LC_26_8_6  (
            .in0(N__93341),
            .in1(N__93342),
            .in2(N__93304),
            .in3(N__93264),
            .lcout(\quad_counter1.n1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_2_lut_LC_26_9_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_2_lut_LC_26_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_2_lut_LC_26_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_2_lut_LC_26_9_0  (
            .in0(_gnd_net_),
            .in1(N__95321),
            .in2(_gnd_net_),
            .in3(N__93261),
            .lcout(\quad_counter1.n1987 ),
            .ltout(),
            .carryin(bfn_26_9_0_),
            .carryout(\quad_counter1.n30465 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_3_lut_LC_26_9_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_3_lut_LC_26_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_3_lut_LC_26_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_3_lut_LC_26_9_1  (
            .in0(_gnd_net_),
            .in1(N__98777),
            .in2(N__95246),
            .in3(N__93258),
            .lcout(\quad_counter1.n1986 ),
            .ltout(),
            .carryin(\quad_counter1.n30465 ),
            .carryout(\quad_counter1.n30466 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_4_lut_LC_26_9_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_4_lut_LC_26_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_4_lut_LC_26_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_4_lut_LC_26_9_2  (
            .in0(_gnd_net_),
            .in1(N__95124),
            .in2(_gnd_net_),
            .in3(N__93255),
            .lcout(\quad_counter1.n1985 ),
            .ltout(),
            .carryin(\quad_counter1.n30466 ),
            .carryout(\quad_counter1.n30467 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_5_lut_LC_26_9_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_5_lut_LC_26_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_5_lut_LC_26_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_5_lut_LC_26_9_3  (
            .in0(_gnd_net_),
            .in1(N__95142),
            .in2(_gnd_net_),
            .in3(N__93252),
            .lcout(\quad_counter1.n1984 ),
            .ltout(),
            .carryin(\quad_counter1.n30467 ),
            .carryout(\quad_counter1.n30468 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_6_lut_LC_26_9_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_6_lut_LC_26_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_6_lut_LC_26_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_6_lut_LC_26_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__95094),
            .in3(N__93249),
            .lcout(\quad_counter1.n1983 ),
            .ltout(),
            .carryin(\quad_counter1.n30468 ),
            .carryout(\quad_counter1.n30469 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_7_lut_LC_26_9_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_7_lut_LC_26_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_7_lut_LC_26_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_7_lut_LC_26_9_5  (
            .in0(_gnd_net_),
            .in1(N__95065),
            .in2(_gnd_net_),
            .in3(N__93246),
            .lcout(\quad_counter1.n1982 ),
            .ltout(),
            .carryin(\quad_counter1.n30469 ),
            .carryout(\quad_counter1.n30470 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_8_lut_LC_26_9_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1348_8_lut_LC_26_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_8_lut_LC_26_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1348_8_lut_LC_26_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__100034),
            .in3(N__93243),
            .lcout(\quad_counter1.n1981 ),
            .ltout(),
            .carryin(\quad_counter1.n30470 ),
            .carryout(\quad_counter1.n30471 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1348_9_lut_LC_26_9_7 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1348_9_lut_LC_26_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1348_9_lut_LC_26_9_7 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \quad_counter1.mod_61_add_1348_9_lut_LC_26_9_7  (
            .in0(N__98778),
            .in1(N__95175),
            .in2(N__99996),
            .in3(N__93519),
            .lcout(\quad_counter1.n2012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23563_2_lut_LC_26_10_0 .C_ON=1'b0;
    defparam \quad_counter1.i23563_2_lut_LC_26_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23563_2_lut_LC_26_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23563_2_lut_LC_26_10_0  (
            .in0(_gnd_net_),
            .in1(N__93502),
            .in2(_gnd_net_),
            .in3(N__95527),
            .lcout(),
            .ltout(\quad_counter1.n28279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1258_LC_26_10_1 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1258_LC_26_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1258_LC_26_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1258_LC_26_10_1  (
            .in0(N__95473),
            .in1(N__95410),
            .in2(N__93516),
            .in3(N__95506),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_4_lut_LC_26_10_2 .C_ON=1'b0;
    defparam \quad_counter1.i2_4_lut_LC_26_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_4_lut_LC_26_10_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i2_4_lut_LC_26_10_2  (
            .in0(N__95431),
            .in1(N__95346),
            .in2(N__93513),
            .in3(N__95452),
            .lcout(),
            .ltout(\quad_counter1.n7_adj_4436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1259_LC_26_10_3 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1259_LC_26_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1259_LC_26_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1259_LC_26_10_3  (
            .in0(N__95389),
            .in1(N__95622),
            .in2(N__93510),
            .in3(N__95365),
            .lcout(\quad_counter1.n2243 ),
            .ltout(\quad_counter1.n2243_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30709_1_lut_LC_26_10_4 .C_ON=1'b0;
    defparam \quad_counter1.i30709_1_lut_LC_26_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30709_1_lut_LC_26_10_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30709_1_lut_LC_26_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__93507),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_2_lut_LC_26_11_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_2_lut_LC_26_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_2_lut_LC_26_11_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1549_2_lut_LC_26_11_0  (
            .in0(N__93504),
            .in1(N__93503),
            .in2(N__93697),
            .in3(N__93444),
            .lcout(\quad_counter1.n2319 ),
            .ltout(),
            .carryin(bfn_26_11_0_),
            .carryout(\quad_counter1.n30489 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_3_lut_LC_26_11_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_3_lut_LC_26_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_3_lut_LC_26_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1549_3_lut_LC_26_11_1  (
            .in0(N__95529),
            .in1(N__95528),
            .in2(N__93551),
            .in3(N__93411),
            .lcout(\quad_counter1.n2318 ),
            .ltout(),
            .carryin(\quad_counter1.n30489 ),
            .carryout(\quad_counter1.n30490 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_4_lut_LC_26_11_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_4_lut_LC_26_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_4_lut_LC_26_11_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1549_4_lut_LC_26_11_2  (
            .in0(N__95508),
            .in1(N__95507),
            .in2(N__93698),
            .in3(N__93384),
            .lcout(\quad_counter1.n2317 ),
            .ltout(),
            .carryin(\quad_counter1.n30490 ),
            .carryout(\quad_counter1.n30491 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_5_lut_LC_26_11_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_5_lut_LC_26_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_5_lut_LC_26_11_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1549_5_lut_LC_26_11_3  (
            .in0(N__95475),
            .in1(N__95474),
            .in2(N__93701),
            .in3(N__93759),
            .lcout(\quad_counter1.n2316 ),
            .ltout(),
            .carryin(\quad_counter1.n30491 ),
            .carryout(\quad_counter1.n30492 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_6_lut_LC_26_11_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_6_lut_LC_26_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_6_lut_LC_26_11_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1549_6_lut_LC_26_11_4  (
            .in0(N__95454),
            .in1(N__95453),
            .in2(N__93699),
            .in3(N__93732),
            .lcout(\quad_counter1.n2315 ),
            .ltout(),
            .carryin(\quad_counter1.n30492 ),
            .carryout(\quad_counter1.n30493 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_7_lut_LC_26_11_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_7_lut_LC_26_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_7_lut_LC_26_11_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1549_7_lut_LC_26_11_5  (
            .in0(N__95433),
            .in1(N__95432),
            .in2(N__93702),
            .in3(N__93705),
            .lcout(\quad_counter1.n2314 ),
            .ltout(),
            .carryin(\quad_counter1.n30493 ),
            .carryout(\quad_counter1.n30494 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_8_lut_LC_26_11_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_8_lut_LC_26_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_8_lut_LC_26_11_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1549_8_lut_LC_26_11_6  (
            .in0(N__95412),
            .in1(N__95411),
            .in2(N__93700),
            .in3(N__93627),
            .lcout(\quad_counter1.n2313 ),
            .ltout(),
            .carryin(\quad_counter1.n30494 ),
            .carryout(\quad_counter1.n30495 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_9_lut_LC_26_11_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_9_lut_LC_26_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_9_lut_LC_26_11_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1549_9_lut_LC_26_11_7  (
            .in0(N__95391),
            .in1(N__95390),
            .in2(N__93552),
            .in3(N__93624),
            .lcout(\quad_counter1.n2312 ),
            .ltout(),
            .carryin(\quad_counter1.n30495 ),
            .carryout(\quad_counter1.n30496 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_10_lut_LC_26_12_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_10_lut_LC_26_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_10_lut_LC_26_12_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1549_10_lut_LC_26_12_0  (
            .in0(N__95370),
            .in1(N__95366),
            .in2(N__93562),
            .in3(N__93594),
            .lcout(\quad_counter1.n2311 ),
            .ltout(),
            .carryin(bfn_26_12_0_),
            .carryout(\quad_counter1.n30497 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_11_lut_LC_26_12_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1549_11_lut_LC_26_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_11_lut_LC_26_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1549_11_lut_LC_26_12_1  (
            .in0(N__95345),
            .in1(N__95344),
            .in2(N__93564),
            .in3(N__93567),
            .lcout(\quad_counter1.n2310 ),
            .ltout(),
            .carryin(\quad_counter1.n30497 ),
            .carryout(\quad_counter1.n30498 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1549_12_lut_LC_26_12_2 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1549_12_lut_LC_26_12_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1549_12_lut_LC_26_12_2 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1549_12_lut_LC_26_12_2  (
            .in0(N__95620),
            .in1(N__95621),
            .in2(N__93563),
            .in3(N__93522),
            .lcout(\quad_counter1.n2309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_adj_1261_LC_26_12_7 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_adj_1261_LC_26_12_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_adj_1261_LC_26_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i2_2_lut_adj_1261_LC_26_12_7  (
            .in0(_gnd_net_),
            .in1(N__93944),
            .in2(_gnd_net_),
            .in3(N__93920),
            .lcout(\quad_counter1.n8_adj_4438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1922_LC_26_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1922_LC_26_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1922_LC_26_17_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1922_LC_26_17_0  (
            .in0(N__100102),
            .in1(N__101205),
            .in2(N__101343),
            .in3(N__100782),
            .lcout(),
            .ltout(\c0.n6_adj_4533_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__2__5299_LC_26_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__2__5299_LC_26_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__2__5299_LC_26_17_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__2__5299_LC_26_17_1  (
            .in0(N__100116),
            .in1(N__94095),
            .in2(N__93897),
            .in3(N__94035),
            .lcout(\c0.data_out_frame_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97715),
            .ce(N__96969),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_26_17_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_26_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_26_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_26_17_2  (
            .in0(N__96170),
            .in1(N__93894),
            .in2(_gnd_net_),
            .in3(N__95535),
            .lcout(\c0.n26_adj_4512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1731_LC_26_17_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1731_LC_26_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1731_LC_26_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1731_LC_26_17_3  (
            .in0(N__94928),
            .in1(N__96217),
            .in2(N__94021),
            .in3(N__94420),
            .lcout(\c0.n32271 ),
            .ltout(\c0.n32271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__1__5300_LC_26_17_4 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__1__5300_LC_26_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__1__5300_LC_26_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_frame_28__1__5300_LC_26_17_4  (
            .in0(_gnd_net_),
            .in1(N__96332),
            .in2(N__93870),
            .in3(N__101388),
            .lcout(\c0.data_out_frame_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97715),
            .ce(N__96969),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_26_17_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_26_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_26_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_26_17_5  (
            .in0(N__95589),
            .in1(N__93867),
            .in2(_gnd_net_),
            .in3(N__96169),
            .lcout(\c0.n26_adj_4506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__4__5297_LC_26_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__4__5297_LC_26_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__4__5297_LC_26_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__4__5297_LC_26_17_6  (
            .in0(N__96218),
            .in1(N__94015),
            .in2(N__98397),
            .in3(N__93830),
            .lcout(\c0.data_out_frame_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97715),
            .ce(N__96969),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1720_LC_26_18_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1720_LC_26_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1720_LC_26_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1720_LC_26_18_0  (
            .in0(N__94112),
            .in1(N__93831),
            .in2(N__93810),
            .in3(N__98034),
            .lcout(\c0.n32300 ),
            .ltout(\c0.n32300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1521_LC_26_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1521_LC_26_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1521_LC_26_18_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1521_LC_26_18_1  (
            .in0(N__94022),
            .in1(N__94094),
            .in2(N__94083),
            .in3(N__94034),
            .lcout(\c0.n32445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1347_LC_26_18_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1347_LC_26_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1347_LC_26_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1347_LC_26_18_2  (
            .in0(N__98168),
            .in1(N__94080),
            .in2(_gnd_net_),
            .in3(N__96810),
            .lcout(\c0.n32454 ),
            .ltout(\c0.n32454_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_26_18_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_26_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_26_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_26_18_3  (
            .in0(N__96328),
            .in1(N__96882),
            .in2(N__94044),
            .in3(N__101001),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1735_LC_26_18_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1735_LC_26_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1735_LC_26_18_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1735_LC_26_18_4  (
            .in0(N__94041),
            .in1(N__96417),
            .in2(N__93992),
            .in3(N__98111),
            .lcout(\c0.n35212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1775_LC_26_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1775_LC_26_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1775_LC_26_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1775_LC_26_18_5  (
            .in0(N__100099),
            .in1(N__98261),
            .in2(_gnd_net_),
            .in3(N__100999),
            .lcout(\c0.n31516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1497_LC_26_18_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1497_LC_26_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1497_LC_26_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1497_LC_26_18_6  (
            .in0(N__101000),
            .in1(N__96734),
            .in2(N__98274),
            .in3(N__100100),
            .lcout(\c0.n32331 ),
            .ltout(\c0.n32331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1379_LC_26_18_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1379_LC_26_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1379_LC_26_18_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \c0.i2_3_lut_adj_1379_LC_26_18_7  (
            .in0(N__94023),
            .in1(N__93988),
            .in2(N__93972),
            .in3(_gnd_net_),
            .lcout(n35623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1740_LC_26_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1740_LC_26_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1740_LC_26_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1740_LC_26_19_0  (
            .in0(N__94577),
            .in1(N__94535),
            .in2(_gnd_net_),
            .in3(N__98449),
            .lcout(\c0.n32403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_26_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_26_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_26_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_3_lut_3_lut_LC_26_19_1  (
            .in0(_gnd_net_),
            .in1(N__98351),
            .in2(_gnd_net_),
            .in3(N__94576),
            .lcout(\c0.n4_adj_4630 ),
            .ltout(\c0.n4_adj_4630_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__5__5288_LC_26_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__5__5288_LC_26_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__5__5288_LC_26_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__5__5288_LC_26_19_2  (
            .in0(N__95666),
            .in1(N__98119),
            .in2(N__94245),
            .in3(N__100425),
            .lcout(\c0.data_out_frame_29_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97750),
            .ce(N__96999),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1703_LC_26_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1703_LC_26_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1703_LC_26_19_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1703_LC_26_19_3  (
            .in0(N__96729),
            .in1(N__96350),
            .in2(_gnd_net_),
            .in3(N__101387),
            .lcout(\c0.n33557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1724_LC_26_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1724_LC_26_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1724_LC_26_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1724_LC_26_19_4  (
            .in0(N__94235),
            .in1(N__97876),
            .in2(N__100428),
            .in3(N__98118),
            .lcout(\c0.n31283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_26_19_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_26_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_26_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_26_19_5  (
            .in0(N__96183),
            .in1(N__94224),
            .in2(_gnd_net_),
            .in3(N__94215),
            .lcout(\c0.n26_adj_4620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1727_LC_26_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1727_LC_26_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1727_LC_26_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1727_LC_26_19_6  (
            .in0(N__98352),
            .in1(N__98450),
            .in2(N__100427),
            .in3(N__94536),
            .lcout(\c0.n32476 ),
            .ltout(\c0.n32476_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1356_LC_26_19_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1356_LC_26_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1356_LC_26_19_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_4_lut_adj_1356_LC_26_19_7  (
            .in0(N__96863),
            .in1(N__94113),
            .in2(N__94194),
            .in3(N__96837),
            .lcout(\c0.n33855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_1594_LC_26_20_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_1594_LC_26_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_1594_LC_26_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_adj_1594_LC_26_20_0  (
            .in0(N__94191),
            .in1(N__94863),
            .in2(N__94473),
            .in3(N__94158),
            .lcout(\c0.n44_adj_4639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1789_LC_26_20_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1789_LC_26_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1789_LC_26_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1789_LC_26_20_2  (
            .in0(N__94533),
            .in1(N__94924),
            .in2(N__100357),
            .in3(N__94575),
            .lcout(\c0.n33572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_2_lut_LC_26_20_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_2_lut_LC_26_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_2_lut_LC_26_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_3_lut_2_lut_LC_26_20_3  (
            .in0(_gnd_net_),
            .in1(N__96418),
            .in2(_gnd_net_),
            .in3(N__101380),
            .lcout(\c0.n31338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_17_i3_2_lut_LC_26_20_4 .C_ON=1'b0;
    defparam \c0.select_369_Select_17_i3_2_lut_LC_26_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_17_i3_2_lut_LC_26_20_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_17_i3_2_lut_LC_26_20_4  (
            .in0(N__94472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94796),
            .lcout(\c0.n3_adj_4596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1426_LC_26_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1426_LC_26_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1426_LC_26_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1426_LC_26_20_5  (
            .in0(_gnd_net_),
            .in1(N__98275),
            .in2(_gnd_net_),
            .in3(N__100078),
            .lcout(\c0.n31302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1373_LC_26_21_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1373_LC_26_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1373_LC_26_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1373_LC_26_21_0  (
            .in0(N__95009),
            .in1(N__96300),
            .in2(_gnd_net_),
            .in3(N__100415),
            .lcout(),
            .ltout(\c0.n17574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_LC_26_21_1 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_LC_26_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_LC_26_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_3_lut_4_lut_LC_26_21_1  (
            .in0(N__96419),
            .in1(N__98358),
            .in2(N__94437),
            .in3(N__98110),
            .lcout(\c0.n33936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1428_LC_26_21_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1428_LC_26_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1428_LC_26_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1428_LC_26_21_2  (
            .in0(N__94434),
            .in1(N__95576),
            .in2(N__94421),
            .in3(N__98369),
            .lcout(\c0.n33509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1349_LC_26_21_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1349_LC_26_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1349_LC_26_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1349_LC_26_21_3  (
            .in0(N__96420),
            .in1(N__94388),
            .in2(N__95037),
            .in3(N__94370),
            .lcout(\c0.n14_adj_4523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1410_LC_26_21_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1410_LC_26_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1410_LC_26_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1410_LC_26_21_4  (
            .in0(N__94325),
            .in1(N__95051),
            .in2(N__94578),
            .in3(N__100895),
            .lcout(\c0.n31463 ),
            .ltout(\c0.n31463_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1717_LC_26_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1717_LC_26_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1717_LC_26_21_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1717_LC_26_21_5  (
            .in0(N__100896),
            .in1(N__95008),
            .in2(N__94329),
            .in3(N__98447),
            .lcout(\c0.n17576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1487_LC_26_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1487_LC_26_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1487_LC_26_21_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i1_2_lut_adj_1487_LC_26_21_6  (
            .in0(N__94326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__100874),
            .lcout(\c0.n32361 ),
            .ltout(\c0.n32361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1489_LC_26_21_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1489_LC_26_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1489_LC_26_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1489_LC_26_21_7  (
            .in0(N__95052),
            .in1(N__95033),
            .in2(N__95013),
            .in3(N__94572),
            .lcout(\c0.n31857 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_4_lut_adj_2049_LC_26_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_4_lut_adj_2049_LC_26_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_4_lut_adj_2049_LC_26_22_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_4_lut_adj_2049_LC_26_22_1  (
            .in0(N__98344),
            .in1(N__94574),
            .in2(N__95010),
            .in3(N__96299),
            .lcout(\c0.n32457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1517_LC_26_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1517_LC_26_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1517_LC_26_22_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1517_LC_26_22_2  (
            .in0(N__96298),
            .in1(N__101347),
            .in2(N__100836),
            .in3(N__101188),
            .lcout(\c0.n32410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1419_LC_26_22_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1419_LC_26_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1419_LC_26_22_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i8_4_lut_adj_1419_LC_26_22_3  (
            .in0(N__98343),
            .in1(N__100832),
            .in2(N__94962),
            .in3(N__100380),
            .lcout(),
            .ltout(\c0.n20_adj_4549_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_adj_1422_LC_26_22_4 .C_ON=1'b0;
    defparam \c0.i11_3_lut_adj_1422_LC_26_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_adj_1422_LC_26_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_3_lut_adj_1422_LC_26_22_4  (
            .in0(_gnd_net_),
            .in1(N__94941),
            .in2(N__94932),
            .in3(N__98049),
            .lcout(),
            .ltout(\c0.n34466_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1423_LC_26_22_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1423_LC_26_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1423_LC_26_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_1423_LC_26_22_5  (
            .in0(N__94909),
            .in1(N__94889),
            .in2(N__94866),
            .in3(N__98132),
            .lcout(\c0.n33839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_369_Select_21_i3_2_lut_LC_26_22_6 .C_ON=1'b0;
    defparam \c0.select_369_Select_21_i3_2_lut_LC_26_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_369_Select_21_i3_2_lut_LC_26_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.select_369_Select_21_i3_2_lut_LC_26_22_6  (
            .in0(N__94862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__94825),
            .lcout(\c0.n3_adj_4600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1491_LC_26_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1491_LC_26_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1491_LC_26_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1491_LC_26_22_7  (
            .in0(_gnd_net_),
            .in1(N__94573),
            .in2(_gnd_net_),
            .in3(N__94514),
            .lcout(\c0.n15744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1713_LC_26_23_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1713_LC_26_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1713_LC_26_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1713_LC_26_23_3  (
            .in0(N__101112),
            .in1(N__101054),
            .in2(N__100255),
            .in3(N__96510),
            .lcout(\c0.n31878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1550_LC_26_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1550_LC_26_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1550_LC_26_23_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1550_LC_26_23_7  (
            .in0(N__98033),
            .in1(N__96297),
            .in2(N__101349),
            .in3(N__101196),
            .lcout(\c0.n31387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23790_4_lut_LC_27_9_0 .C_ON=1'b0;
    defparam \quad_counter1.i23790_4_lut_LC_27_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23790_4_lut_LC_27_9_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \quad_counter1.i23790_4_lut_LC_27_9_0  (
            .in0(N__95109),
            .in1(N__95174),
            .in2(N__95070),
            .in3(N__95089),
            .lcout(\quad_counter1.n1946 ),
            .ltout(\quad_counter1.n1946_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1355_3_lut_LC_27_9_1 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1355_3_lut_LC_27_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1355_3_lut_LC_27_9_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter1.mod_61_i1355_3_lut_LC_27_9_1  (
            .in0(_gnd_net_),
            .in1(N__95123),
            .in2(N__95163),
            .in3(N__95160),
            .lcout(\quad_counter1.n2017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1354_3_lut_LC_27_9_2 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1354_3_lut_LC_27_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1354_3_lut_LC_27_9_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \quad_counter1.mod_61_i1354_3_lut_LC_27_9_2  (
            .in0(_gnd_net_),
            .in1(N__99982),
            .in2(N__95154),
            .in3(N__95141),
            .lcout(\quad_counter1.n2016 ),
            .ltout(\quad_counter1.n2016_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_2_lut_LC_27_9_3 .C_ON=1'b0;
    defparam \quad_counter1.i3_2_lut_LC_27_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_2_lut_LC_27_9_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter1.i3_2_lut_LC_27_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__95145),
            .in3(N__99832),
            .lcout(\quad_counter1.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23569_2_lut_LC_27_9_4 .C_ON=1'b0;
    defparam \quad_counter1.i23569_2_lut_LC_27_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23569_2_lut_LC_27_9_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \quad_counter1.i23569_2_lut_LC_27_9_4  (
            .in0(_gnd_net_),
            .in1(N__95322),
            .in2(_gnd_net_),
            .in3(N__95239),
            .lcout(),
            .ltout(\quad_counter1.n28285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1253_LC_27_9_5 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1253_LC_27_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1253_LC_27_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1253_LC_27_9_5  (
            .in0(N__95140),
            .in1(N__100027),
            .in2(N__95127),
            .in3(N__95122),
            .lcout(\quad_counter1.n10_adj_4431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1353_3_lut_LC_27_9_6 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1353_3_lut_LC_27_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1353_3_lut_LC_27_9_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \quad_counter1.mod_61_i1353_3_lut_LC_27_9_6  (
            .in0(_gnd_net_),
            .in1(N__99981),
            .in2(N__95103),
            .in3(N__95090),
            .lcout(\quad_counter1.n2015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1352_3_lut_LC_27_9_7 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1352_3_lut_LC_27_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1352_3_lut_LC_27_9_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \quad_counter1.mod_61_i1352_3_lut_LC_27_9_7  (
            .in0(N__95076),
            .in1(N__95069),
            .in2(N__99994),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n2014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1357_3_lut_LC_27_10_0 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1357_3_lut_LC_27_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1357_3_lut_LC_27_10_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter1.mod_61_i1357_3_lut_LC_27_10_0  (
            .in0(_gnd_net_),
            .in1(N__95320),
            .in2(N__95283),
            .in3(N__99986),
            .lcout(\quad_counter1.n2019 ),
            .ltout(\quad_counter1.n2019_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i23567_2_lut_LC_27_10_1 .C_ON=1'b0;
    defparam \quad_counter1.i23567_2_lut_LC_27_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i23567_2_lut_LC_27_10_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \quad_counter1.i23567_2_lut_LC_27_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__95274),
            .in3(N__99929),
            .lcout(),
            .ltout(\quad_counter1.n28283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i4_4_lut_adj_1254_LC_27_10_2 .C_ON=1'b0;
    defparam \quad_counter1.i4_4_lut_adj_1254_LC_27_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i4_4_lut_adj_1254_LC_27_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i4_4_lut_adj_1254_LC_27_10_2  (
            .in0(N__99952),
            .in1(N__99869),
            .in2(N__95271),
            .in3(N__99778),
            .lcout(),
            .ltout(\quad_counter1.n10_adj_4432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i28696_4_lut_LC_27_10_3 .C_ON=1'b0;
    defparam \quad_counter1.i28696_4_lut_LC_27_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i28696_4_lut_LC_27_10_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \quad_counter1.i28696_4_lut_LC_27_10_3  (
            .in0(N__95268),
            .in1(N__99808),
            .in2(N__95262),
            .in3(N__98468),
            .lcout(\quad_counter1.n2045 ),
            .ltout(\quad_counter1.n2045_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1421_3_lut_LC_27_10_4 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1421_3_lut_LC_27_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1421_3_lut_LC_27_10_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter1.mod_61_i1421_3_lut_LC_27_10_4  (
            .in0(_gnd_net_),
            .in1(N__99638),
            .in2(N__95259),
            .in3(N__99624),
            .lcout(\quad_counter1.n2115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1424_3_lut_LC_27_10_5 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1424_3_lut_LC_27_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1424_3_lut_LC_27_10_5 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \quad_counter1.mod_61_i1424_3_lut_LC_27_10_5  (
            .in0(N__99654),
            .in1(N__99757),
            .in2(N__99672),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n2118 ),
            .ltout(\quad_counter1.n2118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i1_3_lut_adj_1256_LC_27_10_6 .C_ON=1'b0;
    defparam \quad_counter1.i1_3_lut_adj_1256_LC_27_10_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i1_3_lut_adj_1256_LC_27_10_6 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \quad_counter1.i1_3_lut_adj_1256_LC_27_10_6  (
            .in0(_gnd_net_),
            .in1(N__95221),
            .in2(N__95256),
            .in3(N__99886),
            .lcout(\quad_counter1.n7_adj_4434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1356_3_lut_LC_27_10_7 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1356_3_lut_LC_27_10_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1356_3_lut_LC_27_10_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \quad_counter1.mod_61_i1356_3_lut_LC_27_10_7  (
            .in0(N__95253),
            .in1(_gnd_net_),
            .in2(N__99995),
            .in3(N__95247),
            .lcout(\quad_counter1.n2018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_2_lut_LC_27_11_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_2_lut_LC_27_11_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_2_lut_LC_27_11_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1482_2_lut_LC_27_11_0  (
            .in0(N__95223),
            .in1(N__95222),
            .in2(N__100465),
            .in3(N__95511),
            .lcout(\quad_counter1.n2219 ),
            .ltout(),
            .carryin(bfn_27_11_0_),
            .carryout(\quad_counter1.n30480 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_3_lut_LC_27_11_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_3_lut_LC_27_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_3_lut_LC_27_11_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1482_3_lut_LC_27_11_1  (
            .in0(N__99888),
            .in1(N__99887),
            .in2(N__100503),
            .in3(N__95490),
            .lcout(\quad_counter1.n2218 ),
            .ltout(),
            .carryin(\quad_counter1.n30480 ),
            .carryout(\quad_counter1.n30481 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_4_lut_LC_27_11_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_4_lut_LC_27_11_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_4_lut_LC_27_11_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1482_4_lut_LC_27_11_2  (
            .in0(N__95487),
            .in1(N__95486),
            .in2(N__100466),
            .in3(N__95457),
            .lcout(\quad_counter1.n2217 ),
            .ltout(),
            .carryin(\quad_counter1.n30481 ),
            .carryout(\quad_counter1.n30482 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_5_lut_LC_27_11_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_5_lut_LC_27_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_5_lut_LC_27_11_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1482_5_lut_LC_27_11_3  (
            .in0(N__99711),
            .in1(N__99710),
            .in2(N__100469),
            .in3(N__95436),
            .lcout(\quad_counter1.n2216 ),
            .ltout(),
            .carryin(\quad_counter1.n30482 ),
            .carryout(\quad_counter1.n30483 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_6_lut_LC_27_11_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_6_lut_LC_27_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_6_lut_LC_27_11_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1482_6_lut_LC_27_11_4  (
            .in0(N__100619),
            .in1(N__100620),
            .in2(N__100467),
            .in3(N__95415),
            .lcout(\quad_counter1.n2215 ),
            .ltout(),
            .carryin(\quad_counter1.n30483 ),
            .carryout(\quad_counter1.n30484 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_7_lut_LC_27_11_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_7_lut_LC_27_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_7_lut_LC_27_11_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1482_7_lut_LC_27_11_5  (
            .in0(N__100589),
            .in1(N__100590),
            .in2(N__100470),
            .in3(N__95394),
            .lcout(\quad_counter1.n2214 ),
            .ltout(),
            .carryin(\quad_counter1.n30484 ),
            .carryout(\quad_counter1.n30485 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_8_lut_LC_27_11_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_8_lut_LC_27_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_8_lut_LC_27_11_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \quad_counter1.mod_61_add_1482_8_lut_LC_27_11_6  (
            .in0(N__99696),
            .in1(N__99695),
            .in2(N__100468),
            .in3(N__95373),
            .lcout(\quad_counter1.n2213 ),
            .ltout(),
            .carryin(\quad_counter1.n30485 ),
            .carryout(\quad_counter1.n30486 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_9_lut_LC_27_11_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_9_lut_LC_27_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_9_lut_LC_27_11_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1482_9_lut_LC_27_11_7  (
            .in0(N__100569),
            .in1(N__100568),
            .in2(N__100504),
            .in3(N__95349),
            .lcout(\quad_counter1.n2212 ),
            .ltout(),
            .carryin(\quad_counter1.n30486 ),
            .carryout(\quad_counter1.n30487 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_10_lut_LC_27_12_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1482_10_lut_LC_27_12_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_10_lut_LC_27_12_0 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1482_10_lut_LC_27_12_0  (
            .in0(N__100551),
            .in1(N__100550),
            .in2(N__100505),
            .in3(N__95325),
            .lcout(\quad_counter1.n2211 ),
            .ltout(),
            .carryin(bfn_27_12_0_),
            .carryout(\quad_counter1.n30488 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1482_11_lut_LC_27_12_1 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1482_11_lut_LC_27_12_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1482_11_lut_LC_27_12_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \quad_counter1.mod_61_add_1482_11_lut_LC_27_12_1  (
            .in0(N__100530),
            .in1(N__100529),
            .in2(N__100506),
            .in3(N__95625),
            .lcout(\quad_counter1.n2210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__3__5290_LC_27_16_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__3__5290_LC_27_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__3__5290_LC_27_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_frame_29__3__5290_LC_27_16_0  (
            .in0(N__96698),
            .in1(N__96819),
            .in2(_gnd_net_),
            .in3(N__96246),
            .lcout(\c0.data_out_frame_29_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97716),
            .ce(N__96948),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__1__5292_LC_27_17_0 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__1__5292_LC_27_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__1__5292_LC_27_17_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__1__5292_LC_27_17_0  (
            .in0(N__95544),
            .in1(N__96242),
            .in2(N__96699),
            .in3(N__96818),
            .lcout(\c0.data_out_frame_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97732),
            .ce(N__96988),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1346_LC_27_17_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1346_LC_27_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1346_LC_27_17_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i7_4_lut_adj_1346_LC_27_17_2  (
            .in0(N__96356),
            .in1(N__96239),
            .in2(N__96674),
            .in3(N__100268),
            .lcout(),
            .ltout(\c0.data_out_frame_29__2__N_1749_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__0__5293_LC_27_17_3 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__0__5293_LC_27_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__0__5293_LC_27_17_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.data_out_frame_29__0__5293_LC_27_17_3  (
            .in0(N__96241),
            .in1(_gnd_net_),
            .in2(N__95583),
            .in3(N__95543),
            .lcout(\c0.data_out_frame_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97732),
            .ce(N__96988),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_27_17_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_27_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_27_17_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_27_17_4  (
            .in0(N__95580),
            .in1(N__96372),
            .in2(N__100326),
            .in3(N__95642),
            .lcout(),
            .ltout(\c0.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_LC_27_17_5 .C_ON=1'b0;
    defparam \c0.i11_3_lut_LC_27_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_LC_27_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i11_3_lut_LC_27_17_5  (
            .in0(_gnd_net_),
            .in1(N__95565),
            .in2(N__95553),
            .in3(N__95550),
            .lcout(\c0.n31403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__2__5291_LC_27_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__2__5291_LC_27_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__2__5291_LC_27_17_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_29__2__5291_LC_27_17_6  (
            .in0(N__96357),
            .in1(N__96240),
            .in2(N__96675),
            .in3(N__100269),
            .lcout(\c0.data_out_frame_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97732),
            .ce(N__96988),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1716_LC_27_18_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1716_LC_27_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_1716_LC_27_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_1716_LC_27_18_0  (
            .in0(N__101046),
            .in1(N__96512),
            .in2(N__98457),
            .in3(N__96451),
            .lcout(),
            .ltout(\c0.n7_adj_4521_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_27_18_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_27_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_27_18_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_LC_27_18_1  (
            .in0(N__100319),
            .in1(N__96296),
            .in2(N__96249),
            .in3(N__98120),
            .lcout(\c0.data_out_frame_29__4__N_1639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1714_LC_27_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1714_LC_27_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1714_LC_27_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1714_LC_27_18_2  (
            .in0(N__100159),
            .in1(N__101045),
            .in2(_gnd_net_),
            .in3(N__96511),
            .lcout(\c0.n33588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1382_LC_27_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1382_LC_27_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1382_LC_27_18_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_1382_LC_27_18_3  (
            .in0(N__101100),
            .in1(N__100161),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n33656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1756_LC_27_18_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1756_LC_27_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1756_LC_27_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1756_LC_27_18_4  (
            .in0(N__100160),
            .in1(N__101099),
            .in2(N__100776),
            .in3(N__100670),
            .lcout(\c0.n32383 ),
            .ltout(\c0.n32383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__0__5301_LC_27_18_5 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__0__5301_LC_27_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__0__5301_LC_27_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame_28__0__5301_LC_27_18_5  (
            .in0(N__96222),
            .in1(N__98121),
            .in2(N__96198),
            .in3(N__96371),
            .lcout(\c0.data_out_frame_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97751),
            .ce(N__96995),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_27_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_27_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_27_18_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_27_18_6  (
            .in0(N__96195),
            .in1(N__96189),
            .in2(_gnd_net_),
            .in3(N__96181),
            .lcout(),
            .ltout(\c0.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i30392_4_lut_LC_27_18_7 .C_ON=1'b0;
    defparam \c0.i30392_4_lut_LC_27_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i30392_4_lut_LC_27_18_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.i30392_4_lut_LC_27_18_7  (
            .in0(N__95829),
            .in1(N__95814),
            .in2(N__95799),
            .in3(N__95796),
            .lcout(\c0.n35819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1498_LC_27_19_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1498_LC_27_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1498_LC_27_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1498_LC_27_19_0  (
            .in0(N__95667),
            .in1(N__97875),
            .in2(N__96531),
            .in3(N__100280),
            .lcout(data_out_frame_29__6__N_1518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_29__7__5286_LC_27_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame_29__7__5286_LC_27_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_29__7__5286_LC_27_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_frame_29__7__5286_LC_27_19_1  (
            .in0(_gnd_net_),
            .in1(N__96530),
            .in2(N__98280),
            .in3(N__96387),
            .lcout(\c0.data_out_frame_29_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97767),
            .ce(N__96998),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1493_LC_27_19_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1493_LC_27_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1493_LC_27_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i4_4_lut_adj_1493_LC_27_19_2  (
            .in0(N__96385),
            .in1(N__96809),
            .in2(N__96733),
            .in3(N__96426),
            .lcout(),
            .ltout(\c0.n10_adj_4573_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1494_LC_27_19_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1494_LC_27_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1494_LC_27_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1494_LC_27_19_3  (
            .in0(_gnd_net_),
            .in1(N__100101),
            .in2(N__96534),
            .in3(N__100990),
            .lcout(\c0.n31236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1715_LC_27_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1715_LC_27_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1715_LC_27_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1715_LC_27_19_4  (
            .in0(N__101055),
            .in1(N__97874),
            .in2(N__96516),
            .in3(N__96458),
            .lcout(\c0.n31372 ),
            .ltout(\c0.n31372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1702_LC_27_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1702_LC_27_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1702_LC_27_19_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1702_LC_27_19_5  (
            .in0(N__96416),
            .in1(N__96725),
            .in2(N__96390),
            .in3(N__101373),
            .lcout(\c0.n32437 ),
            .ltout(\c0.n32437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1730_LC_27_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1730_LC_27_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1730_LC_27_19_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1730_LC_27_19_6  (
            .in0(N__96386),
            .in1(_gnd_net_),
            .in2(N__96375),
            .in3(N__98276),
            .lcout(\c0.n31287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1542_LC_27_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1542_LC_27_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1542_LC_27_19_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1542_LC_27_19_7  (
            .in0(N__100254),
            .in1(N__98448),
            .in2(N__97880),
            .in3(N__98117),
            .lcout(\c0.n32273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1375_LC_27_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1375_LC_27_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1375_LC_27_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1375_LC_27_20_0  (
            .in0(N__96349),
            .in1(N__100958),
            .in2(N__100359),
            .in3(N__100878),
            .lcout(\c0.n4_adj_4525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1358_LC_27_20_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1358_LC_27_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1358_LC_27_20_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i6_4_lut_adj_1358_LC_27_20_1  (
            .in0(N__96333),
            .in1(N__98298),
            .in2(N__96312),
            .in3(N__100304),
            .lcout(),
            .ltout(\c0.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame_28__7__5294_LC_27_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame_28__7__5294_LC_27_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame_28__7__5294_LC_27_20_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame_28__7__5294_LC_27_20_2  (
            .in0(N__97908),
            .in1(N__97881),
            .in2(N__97827),
            .in3(N__96741),
            .lcout(\c0.data_out_frame_28_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__97782),
            .ce(N__96996),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_27_20_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_27_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_27_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_LC_27_20_3  (
            .in0(N__96881),
            .in1(N__96870),
            .in2(N__96864),
            .in3(N__96833),
            .lcout(\c0.n33644 ),
            .ltout(\c0.n33644_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_27_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_27_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_27_20_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_LC_27_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__96822),
            .in3(N__96811),
            .lcout(),
            .ltout(\c0.n31357_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1359_LC_27_20_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1359_LC_27_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1359_LC_27_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1359_LC_27_20_5  (
            .in0(N__100379),
            .in1(N__96776),
            .in2(N__96765),
            .in3(N__96762),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1384_LC_27_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1384_LC_27_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1384_LC_27_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1384_LC_27_21_1  (
            .in0(N__98446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__100253),
            .lcout(\c0.n32355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_27_21_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_27_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_27_21_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \c0.i2_2_lut_LC_27_21_3  (
            .in0(N__96735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__96688),
            .lcout(\c0.n10_adj_4520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1767_LC_27_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1767_LC_27_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1767_LC_27_21_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1767_LC_27_21_4  (
            .in0(N__101337),
            .in1(N__100824),
            .in2(_gnd_net_),
            .in3(N__101202),
            .lcout(\c0.n31468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1462_LC_27_21_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1462_LC_27_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1462_LC_27_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1462_LC_27_21_5  (
            .in0(N__96657),
            .in1(N__96634),
            .in2(N__96570),
            .in3(N__96558),
            .lcout(\c0.n35280 ),
            .ltout(\c0.n35280_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1945_LC_27_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1945_LC_27_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1945_LC_27_21_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1945_LC_27_21_6  (
            .in0(N__98187),
            .in1(N__98445),
            .in2(N__98412),
            .in3(N__100957),
            .lcout(\c0.n31461 ),
            .ltout(\c0.n31461_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1357_LC_27_21_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1357_LC_27_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1357_LC_27_21_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i3_4_lut_adj_1357_LC_27_21_7  (
            .in0(N__98390),
            .in1(N__100414),
            .in2(N__98373),
            .in3(N__98370),
            .lcout(\c0.n8_adj_4529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1390_LC_27_22_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1390_LC_27_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1390_LC_27_22_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_adj_1390_LC_27_22_0  (
            .in0(N__98342),
            .in1(N__98291),
            .in2(_gnd_net_),
            .in3(N__98273),
            .lcout(\c0.n33670 ),
            .ltout(\c0.n33670_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1397_LC_27_22_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1397_LC_27_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1397_LC_27_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1397_LC_27_22_1  (
            .in0(N__100256),
            .in1(N__98205),
            .in2(N__98190),
            .in3(N__100631),
            .lcout(),
            .ltout(\c0.n14_adj_4543_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1398_LC_27_22_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1398_LC_27_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1398_LC_27_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1398_LC_27_22_2  (
            .in0(N__97914),
            .in1(N__98183),
            .in2(N__98172),
            .in3(N__98169),
            .lcout(\c0.n32071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1420_LC_27_22_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1420_LC_27_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1420_LC_27_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1420_LC_27_22_5  (
            .in0(N__100632),
            .in1(N__98087),
            .in2(N__100082),
            .in3(N__98064),
            .lcout(\c0.n19_adj_4550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1396_LC_27_22_7 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1396_LC_27_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1396_LC_27_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_adj_1396_LC_27_22_7  (
            .in0(_gnd_net_),
            .in1(N__98042),
            .in2(_gnd_net_),
            .in3(N__97980),
            .lcout(\c0.n10_adj_4542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_28_8_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_28_8_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_28_8_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_28_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_2_lut_LC_28_9_0 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_2_lut_LC_28_9_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_2_lut_LC_28_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_2_lut_LC_28_9_0  (
            .in0(_gnd_net_),
            .in1(N__99922),
            .in2(_gnd_net_),
            .in3(N__99675),
            .lcout(\quad_counter1.n2087 ),
            .ltout(),
            .carryin(bfn_28_9_0_),
            .carryout(\quad_counter1.n30472 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_3_lut_LC_28_9_1 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_3_lut_LC_28_9_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_3_lut_LC_28_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_3_lut_LC_28_9_1  (
            .in0(_gnd_net_),
            .in1(N__98518),
            .in2(N__99671),
            .in3(N__99648),
            .lcout(\quad_counter1.n2086 ),
            .ltout(),
            .carryin(\quad_counter1.n30472 ),
            .carryout(\quad_counter1.n30473 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_4_lut_LC_28_9_2 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_4_lut_LC_28_9_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_4_lut_LC_28_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_4_lut_LC_28_9_2  (
            .in0(_gnd_net_),
            .in1(N__99779),
            .in2(_gnd_net_),
            .in3(N__99645),
            .lcout(\quad_counter1.n2085 ),
            .ltout(),
            .carryin(\quad_counter1.n30473 ),
            .carryout(\quad_counter1.n30474 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_5_lut_LC_28_9_3 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_5_lut_LC_28_9_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_5_lut_LC_28_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_5_lut_LC_28_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__99870),
            .in3(N__99642),
            .lcout(\quad_counter1.n2084 ),
            .ltout(),
            .carryin(\quad_counter1.n30474 ),
            .carryout(\quad_counter1.n30475 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_6_lut_LC_28_9_4 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_6_lut_LC_28_9_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_6_lut_LC_28_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_6_lut_LC_28_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__99639),
            .in3(N__99618),
            .lcout(\quad_counter1.n2083 ),
            .ltout(),
            .carryin(\quad_counter1.n30475 ),
            .carryout(\quad_counter1.n30476 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_7_lut_LC_28_9_5 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_7_lut_LC_28_9_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_7_lut_LC_28_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_7_lut_LC_28_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__99839),
            .in3(N__99615),
            .lcout(\quad_counter1.n2082 ),
            .ltout(),
            .carryin(\quad_counter1.n30476 ),
            .carryout(\quad_counter1.n30477 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_8_lut_LC_28_9_6 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_8_lut_LC_28_9_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_8_lut_LC_28_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_8_lut_LC_28_9_6  (
            .in0(_gnd_net_),
            .in1(N__99953),
            .in2(_gnd_net_),
            .in3(N__99612),
            .lcout(\quad_counter1.n2081 ),
            .ltout(),
            .carryin(\quad_counter1.n30477 ),
            .carryout(\quad_counter1.n30478 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_9_lut_LC_28_9_7 .C_ON=1'b1;
    defparam \quad_counter1.mod_61_add_1415_9_lut_LC_28_9_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_9_lut_LC_28_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter1.mod_61_add_1415_9_lut_LC_28_9_7  (
            .in0(_gnd_net_),
            .in1(N__99809),
            .in2(N__98748),
            .in3(N__99609),
            .lcout(\quad_counter1.n2080 ),
            .ltout(),
            .carryin(\quad_counter1.n30478 ),
            .carryout(\quad_counter1.n30479 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_add_1415_10_lut_LC_28_10_0 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_add_1415_10_lut_LC_28_10_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_add_1415_10_lut_LC_28_10_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \quad_counter1.mod_61_add_1415_10_lut_LC_28_10_0  (
            .in0(N__98589),
            .in1(N__98475),
            .in2(N__99761),
            .in3(N__100041),
            .lcout(\quad_counter1.n2111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1351_3_lut_LC_28_10_1 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1351_3_lut_LC_28_10_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1351_3_lut_LC_28_10_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter1.mod_61_i1351_3_lut_LC_28_10_1  (
            .in0(_gnd_net_),
            .in1(N__100038),
            .in2(N__100011),
            .in3(N__99990),
            .lcout(\quad_counter1.n2013 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1419_3_lut_LC_28_10_2 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1419_3_lut_LC_28_10_2 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1419_3_lut_LC_28_10_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter1.mod_61_i1419_3_lut_LC_28_10_2  (
            .in0(_gnd_net_),
            .in1(N__99954),
            .in2(N__99762),
            .in3(N__99936),
            .lcout(\quad_counter1.n2113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1425_3_lut_LC_28_10_3 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1425_3_lut_LC_28_10_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1425_3_lut_LC_28_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \quad_counter1.mod_61_i1425_3_lut_LC_28_10_3  (
            .in0(N__99930),
            .in1(N__99894),
            .in2(_gnd_net_),
            .in3(N__99746),
            .lcout(\quad_counter1.n2119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1422_3_lut_LC_28_10_4 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1422_3_lut_LC_28_10_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1422_3_lut_LC_28_10_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \quad_counter1.mod_61_i1422_3_lut_LC_28_10_4  (
            .in0(_gnd_net_),
            .in1(N__99868),
            .in2(N__99760),
            .in3(N__99846),
            .lcout(\quad_counter1.n2116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1420_3_lut_LC_28_10_5 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1420_3_lut_LC_28_10_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1420_3_lut_LC_28_10_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \quad_counter1.mod_61_i1420_3_lut_LC_28_10_5  (
            .in0(_gnd_net_),
            .in1(N__99747),
            .in2(N__99840),
            .in3(N__99816),
            .lcout(\quad_counter1.n2114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1418_3_lut_LC_28_11_1 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1418_3_lut_LC_28_11_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1418_3_lut_LC_28_11_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \quad_counter1.mod_61_i1418_3_lut_LC_28_11_1  (
            .in0(_gnd_net_),
            .in1(N__99810),
            .in2(N__99792),
            .in3(N__99759),
            .lcout(\quad_counter1.n2112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.mod_61_i1423_3_lut_LC_28_11_3 .C_ON=1'b0;
    defparam \quad_counter1.mod_61_i1423_3_lut_LC_28_11_3 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.mod_61_i1423_3_lut_LC_28_11_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \quad_counter1.mod_61_i1423_3_lut_LC_28_11_3  (
            .in0(N__99780),
            .in1(N__99758),
            .in2(_gnd_net_),
            .in3(N__99720),
            .lcout(\quad_counter1.n2117 ),
            .ltout(\quad_counter1.n2117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i2_2_lut_adj_1255_LC_28_11_4 .C_ON=1'b0;
    defparam \quad_counter1.i2_2_lut_adj_1255_LC_28_11_4 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i2_2_lut_adj_1255_LC_28_11_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \quad_counter1.i2_2_lut_adj_1255_LC_28_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__99699),
            .in3(N__99688),
            .lcout(),
            .ltout(\quad_counter1.n8_adj_4433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i5_4_lut_adj_1257_LC_28_11_5 .C_ON=1'b0;
    defparam \quad_counter1.i5_4_lut_adj_1257_LC_28_11_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i5_4_lut_adj_1257_LC_28_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \quad_counter1.i5_4_lut_adj_1257_LC_28_11_5  (
            .in0(N__100615),
            .in1(N__100599),
            .in2(N__100593),
            .in3(N__100585),
            .lcout(),
            .ltout(\quad_counter1.n34427_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i3_4_lut_LC_28_11_6 .C_ON=1'b0;
    defparam \quad_counter1.i3_4_lut_LC_28_11_6 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i3_4_lut_LC_28_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \quad_counter1.i3_4_lut_LC_28_11_6  (
            .in0(N__100567),
            .in1(N__100549),
            .in2(N__100533),
            .in3(N__100519),
            .lcout(\quad_counter1.n2144 ),
            .ltout(\quad_counter1.n2144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter1.i30710_1_lut_LC_28_11_7 .C_ON=1'b0;
    defparam \quad_counter1.i30710_1_lut_LC_28_11_7 .SEQ_MODE=4'b0000;
    defparam \quad_counter1.i30710_1_lut_LC_28_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \quad_counter1.i30710_1_lut_LC_28_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__100473),
            .in3(_gnd_net_),
            .lcout(\quad_counter1.n36137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1558_LC_28_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1558_LC_28_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1558_LC_28_18_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1558_LC_28_18_4  (
            .in0(N__100959),
            .in1(N__100879),
            .in2(N__100682),
            .in3(N__100426),
            .lcout(\c0.n33960 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1957_LC_28_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1957_LC_28_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1957_LC_28_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1957_LC_28_19_2  (
            .in0(N__100358),
            .in1(N__100940),
            .in2(_gnd_net_),
            .in3(N__100880),
            .lcout(\c0.n32412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_28_20_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_28_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_28_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_28_20_0  (
            .in0(N__100991),
            .in1(N__100308),
            .in2(N__100290),
            .in3(N__100281),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1380_LC_28_20_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1380_LC_28_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1380_LC_28_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1380_LC_28_20_2  (
            .in0(N__100246),
            .in1(N__100167),
            .in2(_gnd_net_),
            .in3(N__100986),
            .lcout(\c0.n33548 ),
            .ltout(\c0.n33548_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1381_LC_28_20_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1381_LC_28_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1381_LC_28_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1381_LC_28_20_3  (
            .in0(_gnd_net_),
            .in1(N__100070),
            .in2(N__101391),
            .in3(N__101111),
            .lcout(\c0.n33635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_3_lut_4_lut_LC_28_20_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_3_lut_4_lut_LC_28_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_3_lut_4_lut_LC_28_20_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.i2_3_lut_3_lut_4_lut_LC_28_20_5  (
            .in0(N__101348),
            .in1(N__101201),
            .in2(_gnd_net_),
            .in3(N__100685),
            .lcout(),
            .ltout(\c0.n33673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1723_LC_28_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1723_LC_28_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1723_LC_28_20_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1723_LC_28_20_6  (
            .in0(N__101110),
            .in1(N__100965),
            .in2(N__101058),
            .in3(N__101050),
            .lcout(\c0.n15782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_3_lut_LC_28_20_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_3_lut_LC_28_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_3_lut_LC_28_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_3_lut_LC_28_20_7  (
            .in0(N__100772),
            .in1(N__100826),
            .in2(_gnd_net_),
            .in3(N__100684),
            .lcout(\c0.n34929 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1409_LC_28_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1409_LC_28_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1409_LC_28_21_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \c0.i1_2_lut_adj_1409_LC_28_21_0  (
            .in0(_gnd_net_),
            .in1(N__100953),
            .in2(_gnd_net_),
            .in3(N__100866),
            .lcout(\c0.n32296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_4_lut_LC_28_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_4_lut_LC_28_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_4_lut_LC_28_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_4_lut_LC_28_21_5  (
            .in0(N__100867),
            .in1(N__100825),
            .in2(N__100781),
            .in3(N__100689),
            .lcout(\c0.n33899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
