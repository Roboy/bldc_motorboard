-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 12 2019 19:45:28

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : inout std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__50887\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50842\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50774\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50745\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50742\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50720\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50699\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50677\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50130\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49725\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49644\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49169\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49006\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41389\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.n17610_cascade_\ : std_logic;
signal \c0.n18214\ : std_logic;
signal \c0.n18217\ : std_logic;
signal \c0.n18094_cascade_\ : std_logic;
signal \c0.n18097_cascade_\ : std_logic;
signal \c0.n18262_cascade_\ : std_logic;
signal \c0.n22_adj_2365\ : std_logic;
signal \c0.n18265_cascade_\ : std_logic;
signal \c0.n10468_cascade_\ : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n15_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_5\ : std_logic;
signal \c0.n17306_cascade_\ : std_logic;
signal data_out_frame2_18_5 : std_logic;
signal \c0.n24_cascade_\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.n17174\ : std_logic;
signal \c0.n17174_cascade_\ : std_logic;
signal \c0.n10356_cascade_\ : std_logic;
signal \c0.n18139\ : std_logic;
signal \c0.n5_adj_2315_cascade_\ : std_logic;
signal data_out_frame2_13_7 : std_logic;
signal \c0.n18022\ : std_logic;
signal \c0.n5_adj_2353_cascade_\ : std_logic;
signal \c0.n6\ : std_logic;
signal \c0.n6_adj_2138\ : std_logic;
signal \c0.n17440\ : std_logic;
signal \c0.n18037_cascade_\ : std_logic;
signal \c0.n18274_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_4\ : std_logic;
signal \c0.n18277_cascade_\ : std_logic;
signal \c0.n22_adj_2367\ : std_logic;
signal \c0.n18034\ : std_logic;
signal \c0.n17225\ : std_logic;
signal \c0.n17135_cascade_\ : std_logic;
signal \c0.n21_cascade_\ : std_logic;
signal \c0.n20_adj_2223\ : std_logic;
signal \c0.n19_adj_2224\ : std_logic;
signal \c0.n14_adj_2308_cascade_\ : std_logic;
signal \c0.n17135\ : std_logic;
signal \c0.n17092_cascade_\ : std_logic;
signal \c0.n17_adj_2294_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_4\ : std_logic;
signal \c0.n12\ : std_logic;
signal data_out_frame2_14_0 : std_logic;
signal \c0.n17237_cascade_\ : std_logic;
signal \c0.n16_adj_2293\ : std_logic;
signal \c0.n18136\ : std_logic;
signal \c0.data_out_frame2_19_2\ : std_logic;
signal \c0.n10520_cascade_\ : std_logic;
signal \c0.n10349\ : std_logic;
signal \c0.n10462\ : std_logic;
signal \c0.n15_adj_2312\ : std_logic;
signal \c0.n17285\ : std_logic;
signal \c0.n10530\ : std_logic;
signal \c0.n10530_cascade_\ : std_logic;
signal \c0.n10371\ : std_logic;
signal data_out_frame2_7_0 : std_logic;
signal data_out_frame2_6_0 : std_logic;
signal \c0.n5_adj_2343\ : std_logic;
signal data_out_frame2_15_5 : std_logic;
signal \c0.n18100_cascade_\ : std_logic;
signal \c0.n18103\ : std_logic;
signal \c0.n18010_cascade_\ : std_logic;
signal \c0.n18013_cascade_\ : std_logic;
signal \c0.n22_adj_2375\ : std_logic;
signal \c0.n18025\ : std_logic;
signal \c0.n18238_cascade_\ : std_logic;
signal \c0.n18241\ : std_logic;
signal data_out_frame2_7_7 : std_logic;
signal \c0.n5_adj_2137\ : std_logic;
signal \c0.n18154\ : std_logic;
signal \c0.n18130_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_7\ : std_logic;
signal \c0.n18133_cascade_\ : std_logic;
signal \c0.n22_adj_2363\ : std_logic;
signal \c0.n18028\ : std_logic;
signal \c0.n18040_cascade_\ : std_logic;
signal \c0.n6_adj_2215\ : std_logic;
signal \c0.n17219\ : std_logic;
signal \c0.n17141\ : std_logic;
signal \c0.n17219_cascade_\ : std_logic;
signal \c0.n17_cascade_\ : std_logic;
signal \c0.n17228\ : std_logic;
signal \c0.n17246_cascade_\ : std_logic;
signal \c0.n17187\ : std_logic;
signal \c0.n33_cascade_\ : std_logic;
signal \c0.data_out_frame2_19_7\ : std_logic;
signal \c0.n30_adj_2218\ : std_logic;
signal \c0.n17300_cascade_\ : std_logic;
signal \c0.n34\ : std_logic;
signal \c0.n17237\ : std_logic;
signal \c0.n10440\ : std_logic;
signal \c0.n17569\ : std_logic;
signal data_out_frame2_17_5 : std_logic;
signal \c0.n17138\ : std_logic;
signal \c0.n6_adj_2228_cascade_\ : std_logic;
signal \c0.n17312\ : std_logic;
signal data_out_frame2_14_3 : std_logic;
signal \c0.n17267\ : std_logic;
signal data_out_frame2_13_2 : std_logic;
signal \c0.n17309\ : std_logic;
signal \c0.n17291\ : std_logic;
signal \c0.n17303\ : std_logic;
signal \c0.n25\ : std_logic;
signal \c0.n28_adj_2200_cascade_\ : std_logic;
signal \c0.n27_adj_2204\ : std_logic;
signal \c0.n10223_cascade_\ : std_logic;
signal \c0.n6_adj_2318\ : std_logic;
signal data_out_frame2_9_1 : std_logic;
signal \c0.n10346\ : std_logic;
signal \c0.n17231\ : std_logic;
signal \c0.n18076\ : std_logic;
signal data_out_frame2_9_5 : std_logic;
signal \c0.n18109\ : std_logic;
signal data_out_frame2_6_3 : std_logic;
signal \c0.n10334_cascade_\ : std_logic;
signal \c0.n10533\ : std_logic;
signal \c0.n10_adj_2297\ : std_logic;
signal \c0.n14_adj_2296_cascade_\ : std_logic;
signal tx2_enable : std_logic;
signal \c0.n3_adj_2232\ : std_logic;
signal \c0.n3_adj_2278\ : std_logic;
signal \c0.n3_adj_2266\ : std_logic;
signal \c0.data_out_frame2_19_6\ : std_logic;
signal \c0.n18178_cascade_\ : std_logic;
signal \c0.n6_adj_2161\ : std_logic;
signal \c0.n18181\ : std_logic;
signal data_out_frame2_16_6 : std_logic;
signal \c0.n18112\ : std_logic;
signal data_out_frame2_17_6 : std_logic;
signal \c0.data_out_frame2_20_6\ : std_logic;
signal \c0.n18115_cascade_\ : std_logic;
signal \c0.n22_adj_2364\ : std_logic;
signal data_out_frame2_18_6 : std_logic;
signal \c0.n18031\ : std_logic;
signal \c0.n10548\ : std_logic;
signal \c0.n10437\ : std_logic;
signal \c0.n17249_cascade_\ : std_logic;
signal \c0.n12_adj_2298\ : std_logic;
signal data_out_frame2_8_1 : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.n17678\ : std_logic;
signal \c0.n17279\ : std_logic;
signal \c0.data_out_frame2_20_1\ : std_logic;
signal data_out_frame2_13_0 : std_logic;
signal \c0.n10424\ : std_logic;
signal \c0.n14_adj_2346\ : std_logic;
signal \c0.n15_adj_2341_cascade_\ : std_logic;
signal data_out_frame2_14_5 : std_logic;
signal \c0.n16_adj_2320_cascade_\ : std_logic;
signal \c0.n17216\ : std_logic;
signal \c0.data_out_frame2_19_1\ : std_logic;
signal \c0.n18058\ : std_logic;
signal \c0.n6_adj_2175_cascade_\ : std_logic;
signal \c0.n17258\ : std_logic;
signal data_out_frame2_11_2 : std_logic;
signal \c0.n17171\ : std_logic;
signal \c0.n17132\ : std_logic;
signal \c0.n17184\ : std_logic;
signal \c0.n32\ : std_logic;
signal data_out_frame2_18_4 : std_logic;
signal data_out_frame2_5_5 : std_logic;
signal data_out_frame2_7_3 : std_logic;
signal data_out_frame2_17_4 : std_logic;
signal data_out_frame2_17_7 : std_logic;
signal \c0.n10356\ : std_logic;
signal \c0.n10572\ : std_logic;
signal \c0.n16_adj_2170\ : std_logic;
signal data_out_frame2_6_5 : std_logic;
signal data_out_frame2_6_7 : std_logic;
signal data_out_frame2_16_1 : std_logic;
signal \c0.n17153\ : std_logic;
signal \c0.n17168\ : std_logic;
signal \c0.n17153_cascade_\ : std_logic;
signal \c0.n26_adj_2203\ : std_logic;
signal data_out_frame2_5_7 : std_logic;
signal data_out_frame2_13_3 : std_logic;
signal data_out_frame2_7_6 : std_logic;
signal data_out_frame2_6_4 : std_logic;
signal \c0.n6_adj_2339\ : std_logic;
signal \c0.n10507\ : std_logic;
signal data_out_frame2_15_0 : std_logic;
signal \c0.n17273\ : std_logic;
signal data_out_frame2_9_2 : std_logic;
signal \c0.n18046\ : std_logic;
signal \c0.n17165\ : std_logic;
signal \c0.n10334\ : std_logic;
signal \c0.n10223\ : std_logic;
signal \c0.n10_adj_2190\ : std_logic;
signal \c0.n3_adj_2282\ : std_logic;
signal \c0.n3_adj_2227\ : std_logic;
signal \c0.n3_adj_2179\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_0\ : std_logic;
signal \bfn_4_27_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_1\ : std_logic;
signal \c0.n16079\ : std_logic;
signal \c0.n16080\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_3\ : std_logic;
signal \c0.FRAME_MATCHER_i_3\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_3\ : std_logic;
signal \c0.n16081\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_4\ : std_logic;
signal \c0.FRAME_MATCHER_i_4\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_4\ : std_logic;
signal \c0.n16082\ : std_logic;
signal \c0.n43\ : std_logic;
signal \c0.FRAME_MATCHER_i_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_5\ : std_logic;
signal \c0.n16083\ : std_logic;
signal \c0.n16084\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_7\ : std_logic;
signal \c0.n16085\ : std_logic;
signal \c0.n16086\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_8\ : std_logic;
signal \bfn_4_28_0_\ : std_logic;
signal \c0.n16087\ : std_logic;
signal \c0.n16088\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_11\ : std_logic;
signal \c0.n16089\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_12\ : std_logic;
signal \c0.n16090\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_13\ : std_logic;
signal \c0.n16091\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_14\ : std_logic;
signal \c0.n16092\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_15\ : std_logic;
signal \c0.n16093\ : std_logic;
signal \c0.n16094\ : std_logic;
signal \bfn_4_29_0_\ : std_logic;
signal \c0.n16095\ : std_logic;
signal \c0.n16096\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_19\ : std_logic;
signal \c0.n16097\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_20\ : std_logic;
signal \c0.n16098\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_21\ : std_logic;
signal \c0.n16099\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_22\ : std_logic;
signal \c0.n16100\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_23\ : std_logic;
signal \c0.n16101\ : std_logic;
signal \c0.n16102\ : std_logic;
signal \bfn_4_30_0_\ : std_logic;
signal \c0.n16103\ : std_logic;
signal \c0.n16104\ : std_logic;
signal \c0.n16105\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_28\ : std_logic;
signal \c0.n16106\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_29\ : std_logic;
signal \c0.FRAME_MATCHER_i_29\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_29\ : std_logic;
signal \c0.n16107\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_30\ : std_logic;
signal \c0.n16108\ : std_logic;
signal \c0.n16109\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_31\ : std_logic;
signal \n5244_cascade_\ : std_logic;
signal \n11018_cascade_\ : std_logic;
signal \c0.n18008\ : std_logic;
signal \n13692_cascade_\ : std_logic;
signal \bfn_4_32_0_\ : std_logic;
signal \c0.rx.n16125\ : std_logic;
signal \c0.rx.n16126\ : std_logic;
signal \c0.rx.n16127\ : std_logic;
signal \c0.rx.n16128\ : std_logic;
signal \c0.rx.n16129\ : std_logic;
signal \c0.rx.n16130\ : std_logic;
signal \c0.rx.n16131\ : std_logic;
signal data_out_frame2_18_1 : std_logic;
signal data_out_frame2_5_6 : std_logic;
signal \c0.n14_adj_2188_cascade_\ : std_logic;
signal \c0.n15_adj_2185\ : std_logic;
signal \c0.data_out_frame2_20_2\ : std_logic;
signal data_out_frame2_7_4 : std_logic;
signal \c0.n17240\ : std_logic;
signal \c0.n17240_cascade_\ : std_logic;
signal \c0.n14_adj_2206\ : std_logic;
signal \c0.n17439\ : std_logic;
signal \c0.n17249\ : std_logic;
signal \c0.data_out_frame2_19_5\ : std_logic;
signal \c0.n17116\ : std_logic;
signal \c0.n17234\ : std_logic;
signal \c0.n15_adj_2291\ : std_logic;
signal \c0.n17288\ : std_logic;
signal data_out_frame2_12_4 : std_logic;
signal \c0.n17288_cascade_\ : std_logic;
signal \c0.n14_adj_2292\ : std_logic;
signal \c0.n17294\ : std_logic;
signal \c0.n10428_cascade_\ : std_logic;
signal \c0.n12_adj_2178\ : std_logic;
signal \c0.n10504\ : std_logic;
signal data_out_frame2_17_1 : std_logic;
signal data_out_frame2_9_4 : std_logic;
signal \c0.n17568\ : std_logic;
signal \c0.n10554\ : std_logic;
signal \c0.n10263\ : std_logic;
signal \c0.n15_adj_2205\ : std_logic;
signal \c0.n5_adj_2337\ : std_logic;
signal data_out_frame2_10_2 : std_logic;
signal \c0.n10492\ : std_logic;
signal data_out_frame2_12_5 : std_logic;
signal \c0.n17255\ : std_logic;
signal data_out_frame2_16_4 : std_logic;
signal data_out_frame2_11_1 : std_logic;
signal \c0.n17156\ : std_logic;
signal \c0.n6_adj_2182_cascade_\ : std_logic;
signal \c0.n10229\ : std_logic;
signal \n10725_cascade_\ : std_logic;
signal data_out_frame2_12_7 : std_logic;
signal data_out_frame2_10_3 : std_logic;
signal \c0.n18106\ : std_logic;
signal data_out_frame2_16_2 : std_logic;
signal data_out_frame2_15_2 : std_logic;
signal data_out_frame2_18_2 : std_logic;
signal data_out_frame2_16_5 : std_logic;
signal data_out_frame2_15_4 : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal n15979 : std_logic;
signal n15980 : std_logic;
signal n15981 : std_logic;
signal n15982 : std_logic;
signal n15983 : std_logic;
signal n15984 : std_logic;
signal n15985 : std_logic;
signal n15986 : std_logic;
signal \bfn_5_24_0_\ : std_logic;
signal n15987 : std_logic;
signal n15988 : std_logic;
signal n15989 : std_logic;
signal n15990 : std_logic;
signal n15991 : std_logic;
signal n15992 : std_logic;
signal n15993 : std_logic;
signal n15994 : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal n15995 : std_logic;
signal n15996 : std_logic;
signal n15997 : std_logic;
signal n15998 : std_logic;
signal n15999 : std_logic;
signal n16000 : std_logic;
signal n16001 : std_logic;
signal n16002 : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal n16003 : std_logic;
signal n16004 : std_logic;
signal n16005 : std_logic;
signal n16006 : std_logic;
signal n16007 : std_logic;
signal n16008 : std_logic;
signal n16009 : std_logic;
signal \c0.n3\ : std_logic;
signal \c0.n26_adj_2373_cascade_\ : std_logic;
signal \c0.n3_adj_2280\ : std_logic;
signal \c0.FRAME_MATCHER_i_6\ : std_logic;
signal \c0.n41\ : std_logic;
signal \c0.n3_adj_2261\ : std_logic;
signal \c0.n3_adj_2270\ : std_logic;
signal \c0.n3_adj_2252\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_17\ : std_logic;
signal \c0.n3_adj_2257\ : std_logic;
signal \c0.FRAME_MATCHER_i_17\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_17\ : std_logic;
signal \c0.n3_adj_2248\ : std_logic;
signal \c0.n3_adj_2250\ : std_logic;
signal \c0.n3_adj_2244\ : std_logic;
signal \c0.FRAME_MATCHER_i_21\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_21\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_27\ : std_logic;
signal \c0.n3_adj_2276\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_8\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_9\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_31\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_25\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_26\ : std_logic;
signal \c0.rx.n10845\ : std_logic;
signal n1 : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.n10656\ : std_logic;
signal \n17708_cascade_\ : std_logic;
signal n5244 : std_logic;
signal n11018 : std_logic;
signal \c0.data_out_frame2_20_0\ : std_logic;
signal \c0.n18049\ : std_logic;
signal \c0.n18043\ : std_logic;
signal \c0.n17586\ : std_logic;
signal \c0.n18244_cascade_\ : std_logic;
signal \c0.n6_adj_2140\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.tx2.n18232_cascade_\ : std_logic;
signal \c0.n22_adj_2387\ : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal \c0.n18157\ : std_logic;
signal \c0.n17603\ : std_logic;
signal \c0.n18226_cascade_\ : std_logic;
signal \c0.n18229\ : std_logic;
signal data_out_frame2_10_0 : std_logic;
signal \c0.n18148_cascade_\ : std_logic;
signal \c0.n18151\ : std_logic;
signal data_out_frame2_5_0 : std_logic;
signal \c0.n5_adj_2217\ : std_logic;
signal \c0.n6_adj_2143\ : std_logic;
signal \c0.data_out_frame2_19_3\ : std_logic;
signal \c0.n18052_cascade_\ : std_logic;
signal \c0.data_out_frame2_20_3\ : std_logic;
signal \c0.n18055_cascade_\ : std_logic;
signal \c0.n9157\ : std_logic;
signal \c0.n18061\ : std_logic;
signal \c0.n18256_cascade_\ : std_logic;
signal \c0.n6_adj_2139\ : std_logic;
signal \c0.n22_adj_2371\ : std_logic;
signal \c0.n18259_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal data_out_frame2_10_1 : std_logic;
signal \c0.n17203\ : std_logic;
signal data_out_frame2_8_6 : std_logic;
signal data_out_frame2_9_6 : std_logic;
signal \c0.n18127\ : std_logic;
signal data_out_frame2_18_3 : std_logic;
signal data_out_frame2_17_0 : std_logic;
signal \c0.n18163\ : std_logic;
signal \c0.n18208\ : std_logic;
signal data_out_frame2_17_3 : std_logic;
signal data_out_frame2_14_2 : std_logic;
signal \c0.n10_adj_2207\ : std_logic;
signal data_out_frame2_11_4 : std_logic;
signal data_out_frame2_11_5 : std_logic;
signal \c0.n10359\ : std_logic;
signal data_out_frame2_5_4 : std_logic;
signal data_out_frame2_10_7 : std_logic;
signal \c0.tx2.n13748_cascade_\ : std_logic;
signal data_out_frame2_18_7 : std_logic;
signal data_out_frame2_17_2 : std_logic;
signal data_out_frame2_7_5 : std_logic;
signal \c0.tx2.n10\ : std_logic;
signal tx2_o : std_logic;
signal data_out_frame2_14_7 : std_logic;
signal \c0.tx2.n17322\ : std_logic;
signal \c0.tx2.n17018\ : std_logic;
signal \c0.tx2.r_Clock_Count_0\ : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal \c0.tx2.r_Clock_Count_1\ : std_logic;
signal \c0.tx2.n16132\ : std_logic;
signal \c0.tx2.r_Clock_Count_2\ : std_logic;
signal \c0.tx2.n16133\ : std_logic;
signal \c0.tx2.r_Clock_Count_3\ : std_logic;
signal \c0.tx2.n16134\ : std_logic;
signal \c0.tx2.r_Clock_Count_4\ : std_logic;
signal \c0.tx2.n16135\ : std_logic;
signal \c0.tx2.r_Clock_Count_5\ : std_logic;
signal \c0.tx2.n16136\ : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal \c0.tx2.n16137\ : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal \c0.tx2.n16138\ : std_logic;
signal \c0.tx2.n16139\ : std_logic;
signal \bfn_6_25_0_\ : std_logic;
signal \c0.tx2.r_Clock_Count_8\ : std_logic;
signal \c0.tx2.n10852\ : std_logic;
signal \c0.FRAME_MATCHER_i_8\ : std_logic;
signal \c0.n42\ : std_logic;
signal \c0.n41_adj_2376_cascade_\ : std_logic;
signal \c0.n39_adj_2377\ : std_logic;
signal \c0.n43_adj_2380\ : std_logic;
signal \c0.n48_adj_2379_cascade_\ : std_logic;
signal \c0.n44_adj_2378\ : std_logic;
signal \c0.n9995_cascade_\ : std_logic;
signal \c0.n9995\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_2\ : std_logic;
signal \c0.n3_adj_2286\ : std_logic;
signal \c0.n3_adj_2226\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_2\ : std_logic;
signal \c0.n40\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_24\ : std_logic;
signal \c0.n3_adj_2242\ : std_logic;
signal \c0.n3_adj_2240\ : std_logic;
signal \c0.n3_adj_2234\ : std_logic;
signal \c0.n3_adj_2230\ : std_logic;
signal \c0.n10009_cascade_\ : std_logic;
signal \c0.n3_adj_2181\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_18\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_27\ : std_logic;
signal \c0.FRAME_MATCHER_i_27\ : std_logic;
signal \c0.n3_adj_2236\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_9\ : std_logic;
signal \c0.FRAME_MATCHER_i_9\ : std_logic;
signal \c0.n3_adj_2274\ : std_logic;
signal \c0.rx.n17636\ : std_logic;
signal n17707 : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal \c0.rx.r_Clock_Count_0\ : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \c0.rx.n6\ : std_logic;
signal \c0.rx.n17022_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2094_0_cascade_\ : std_logic;
signal \c0.rx.n17380_cascade_\ : std_logic;
signal \c0.rx.n17635\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2094_0\ : std_logic;
signal \c0.rx.n6_adj_2130\ : std_logic;
signal \c0.n18247\ : std_logic;
signal \c0.n22_adj_2372\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal \c0.n17620\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \c0.tx2.n18082_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal \c0.tx2.n18085_cascade_\ : std_logic;
signal \c0.tx2.n18235\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_2062_cascade_\ : std_logic;
signal n3 : std_logic;
signal \c0.tx2.n13614_cascade_\ : std_logic;
signal \c0.n17587\ : std_logic;
signal \c0.n17107\ : std_logic;
signal data_out_frame2_15_6 : std_logic;
signal data_out_frame2_12_6 : std_logic;
signal \c0.n18118_cascade_\ : std_logic;
signal data_out_frame2_13_6 : std_logic;
signal \c0.n18121\ : std_logic;
signal \c0.tx2.n13614\ : std_logic;
signal n10976 : std_logic;
signal \n10976_cascade_\ : std_logic;
signal \r_Bit_Index_2_adj_2440\ : std_logic;
signal data_out_frame2_5_1 : std_logic;
signal \c0.n6_adj_2142\ : std_logic;
signal \c0.n18064\ : std_logic;
signal \c0.n18067\ : std_logic;
signal n8191 : std_logic;
signal data_out_frame2_6_1 : std_logic;
signal \c0.n5_adj_2289\ : std_logic;
signal data_out_frame2_11_7 : std_logic;
signal \c0.n10413_cascade_\ : std_logic;
signal \c0.n17282\ : std_logic;
signal data_out_frame2_10_6 : std_logic;
signal data_out_frame2_11_6 : std_logic;
signal \c0.n18124\ : std_logic;
signal \c0.data_out_frame2_19_0\ : std_logic;
signal data_out_frame2_18_0 : std_logic;
signal \c0.n18160\ : std_logic;
signal \c0.n10563\ : std_logic;
signal data_out_frame2_13_5 : std_logic;
signal \c0.n17095\ : std_logic;
signal \c0.n31\ : std_logic;
signal data_out_frame2_13_1 : std_logic;
signal data_out_frame2_12_1 : std_logic;
signal \c0.n18019\ : std_logic;
signal data_out_frame2_12_3 : std_logic;
signal data_out_frame2_5_3 : std_logic;
signal \c0.n18142\ : std_logic;
signal data_out_frame2_8_7 : std_logic;
signal data_out_frame2_9_7 : std_logic;
signal \c0.n18145\ : std_logic;
signal \c0.tx2.n9269\ : std_logic;
signal data_out_frame2_5_2 : std_logic;
signal data_out_frame2_10_4 : std_logic;
signal \c0.n10456\ : std_logic;
signal data_out_frame2_10_5 : std_logic;
signal data_out_frame2_11_3 : std_logic;
signal data_out_frame2_14_1 : std_logic;
signal data_out_frame2_15_1 : std_logic;
signal \c0.n18016\ : std_logic;
signal data_out_frame2_12_2 : std_logic;
signal data_out_frame2_7_2 : std_logic;
signal data_out_frame2_6_2 : std_logic;
signal \c0.n5_adj_2290\ : std_logic;
signal data_out_frame2_14_4 : std_logic;
signal data_out_frame2_11_0 : std_logic;
signal \c0.n17276\ : std_logic;
signal n17412 : std_logic;
signal data_out_frame2_9_3 : std_logic;
signal \c0.n6_adj_2197\ : std_logic;
signal data_out_frame2_15_7 : std_logic;
signal \c0.n17123\ : std_logic;
signal data_out_frame2_14_6 : std_logic;
signal \c0.n10434\ : std_logic;
signal data_out_frame2_16_3 : std_logic;
signal data_out_frame2_15_3 : std_logic;
signal \c0.n10482\ : std_logic;
signal data_out_frame2_8_4 : std_logic;
signal data_out_frame2_8_0 : std_logic;
signal \c0.n10513\ : std_logic;
signal data_out_frame2_16_0 : std_logic;
signal \c0.n17098\ : std_logic;
signal data_out_frame2_8_3 : std_logic;
signal \c0.n17_adj_2321\ : std_logic;
signal \c0.n30_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_26\ : std_logic;
signal \c0.FRAME_MATCHER_i_25\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_25\ : std_logic;
signal \c0.FRAME_MATCHER_i_24\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_24\ : std_logic;
signal \c0.FRAME_MATCHER_i_23\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_23\ : std_logic;
signal \c0.FRAME_MATCHER_i_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_20\ : std_logic;
signal \c0.FRAME_MATCHER_i_19\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_19\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_16\ : std_logic;
signal \c0.n3_adj_2254\ : std_logic;
signal \c0.FRAME_MATCHER_i_18\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_18\ : std_logic;
signal \c0.n3_adj_2288\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_1\ : std_logic;
signal \c0.n3_adj_2246\ : std_logic;
signal \c0.FRAME_MATCHER_i_22\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_22\ : std_logic;
signal \c0.FRAME_MATCHER_i_26\ : std_logic;
signal \c0.n3_adj_2238\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_10\ : std_logic;
signal \r_Bit_Index_1_adj_2441\ : std_logic;
signal \r_Bit_Index_0_adj_2442\ : std_logic;
signal n5266 : std_logic;
signal tx_enable : std_logic;
signal n10674 : std_logic;
signal \c0.n17574\ : std_logic;
signal \c0.rx.n10620\ : std_logic;
signal n17361 : std_logic;
signal \c0.rx.r_SM_Main_2_N_2088_2\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_2088_2_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_0\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_12\ : std_logic;
signal \c0.FRAME_MATCHER_i_12\ : std_logic;
signal \c0.n3_adj_2268\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \c0.n15972\ : std_logic;
signal \c0.n15973\ : std_logic;
signal \c0.n15974\ : std_logic;
signal \c0.n17606\ : std_logic;
signal \c0.n15975\ : std_logic;
signal \c0.n15976\ : std_logic;
signal \c0.n15977\ : std_logic;
signal \c0.n15978\ : std_logic;
signal \c0.n17714\ : std_logic;
signal \c0.n17589\ : std_logic;
signal data_out_frame2_7_1 : std_logic;
signal n10725 : std_logic;
signal data_out_frame2_12_0 : std_logic;
signal \r_SM_Main_2_N_2031_1\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \r_SM_Main_2_adj_2438\ : std_logic;
signal n4_adj_2484 : std_logic;
signal \r_SM_Main_1_adj_2439\ : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.n10133_cascade_\ : std_logic;
signal \c0.n6_adj_2356_cascade_\ : std_logic;
signal \c0.n10027_cascade_\ : std_logic;
signal data_in_0_7 : std_logic;
signal data_in_1_3 : std_logic;
signal \c0.n17331_cascade_\ : std_logic;
signal \c0.n17410\ : std_logic;
signal data_in_2_6 : std_logic;
signal \c0.n12_adj_2355\ : std_logic;
signal data_in_2_4 : std_logic;
signal \c0.n4_adj_2150\ : std_logic;
signal \c0.n10133\ : std_logic;
signal \c0.n17406\ : std_logic;
signal data_in_0_6 : std_logic;
signal \c0.FRAME_MATCHER_i_15\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_15\ : std_logic;
signal \c0.FRAME_MATCHER_i_13\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_13\ : std_logic;
signal \c0.FRAME_MATCHER_i_11\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_11\ : std_logic;
signal \c0.FRAME_MATCHER_i_7\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_7\ : std_logic;
signal \c0.n37\ : std_logic;
signal \c0.FRAME_MATCHER_i_28\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_28\ : std_logic;
signal \c0.FRAME_MATCHER_state_13\ : std_logic;
signal \c0.n8_adj_2332\ : std_logic;
signal \c0.FRAME_MATCHER_state_19\ : std_logic;
signal \c0.n8_adj_2328\ : std_logic;
signal \c0.FRAME_MATCHER_state_6\ : std_logic;
signal \c0.n8_adj_2334\ : std_logic;
signal \c0.FRAME_MATCHER_state_12\ : std_logic;
signal \c0.n16708\ : std_logic;
signal \c0.FRAME_MATCHER_state_14\ : std_logic;
signal \c0.n8_adj_2331\ : std_logic;
signal data_out_frame2_16_7 : std_logic;
signal \c0.n17194\ : std_logic;
signal \c0.n10459\ : std_logic;
signal data_in_0_5 : std_logic;
signal data_in_0_4 : std_logic;
signal data_in_0_2 : std_logic;
signal data_in_1_5 : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1278_16\ : std_logic;
signal \c0.FRAME_MATCHER_state_4\ : std_logic;
signal \c0.n16716\ : std_logic;
signal data_in_1_2 : std_logic;
signal \c0.n17388\ : std_logic;
signal \c0.n3_adj_2272\ : std_logic;
signal \c0.FRAME_MATCHER_i_10\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_10\ : std_logic;
signal \c0.n3_adj_2264\ : std_logic;
signal \c0.FRAME_MATCHER_i_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_14\ : std_logic;
signal \c0.FRAME_MATCHER_i_16\ : std_logic;
signal \c0.n10009\ : std_logic;
signal \c0.n3_adj_2259\ : std_logic;
signal n26_adj_2423 : std_logic;
signal \bfn_9_29_0_\ : std_logic;
signal n25_adj_2424 : std_logic;
signal n16041 : std_logic;
signal n24 : std_logic;
signal n16042 : std_logic;
signal n23_adj_2425 : std_logic;
signal n16043 : std_logic;
signal n22_adj_2426 : std_logic;
signal n16044 : std_logic;
signal n21 : std_logic;
signal n16045 : std_logic;
signal n20 : std_logic;
signal n16046 : std_logic;
signal n19 : std_logic;
signal n16047 : std_logic;
signal n16048 : std_logic;
signal n18 : std_logic;
signal \bfn_9_30_0_\ : std_logic;
signal n17 : std_logic;
signal n16049 : std_logic;
signal n16 : std_logic;
signal n16050 : std_logic;
signal n15 : std_logic;
signal n16051 : std_logic;
signal n14 : std_logic;
signal n16052 : std_logic;
signal n13 : std_logic;
signal n16053 : std_logic;
signal n12 : std_logic;
signal n16054 : std_logic;
signal n11 : std_logic;
signal n16055 : std_logic;
signal n16056 : std_logic;
signal n10_adj_2420 : std_logic;
signal \bfn_9_31_0_\ : std_logic;
signal n9_adj_2421 : std_logic;
signal n16057 : std_logic;
signal n8_adj_2412 : std_logic;
signal n16058 : std_logic;
signal n7 : std_logic;
signal n16059 : std_logic;
signal n6_adj_2429 : std_logic;
signal n16060 : std_logic;
signal n16061 : std_logic;
signal n16062 : std_logic;
signal n16063 : std_logic;
signal n16064 : std_logic;
signal \bfn_9_32_0_\ : std_logic;
signal n16065 : std_logic;
signal \c0.n17711\ : std_logic;
signal \c0.n17659\ : std_logic;
signal \c0.n11867_cascade_\ : std_logic;
signal \c0.n4_adj_2187\ : std_logic;
signal \c0.n4_adj_2152\ : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal \c0.n17761\ : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.n4_adj_2155\ : std_logic;
signal \c0.data_in_frame_3_6\ : std_logic;
signal \c0.n15_adj_2310_cascade_\ : std_logic;
signal \c0.data_in_frame_3_3\ : std_logic;
signal \n17075_cascade_\ : std_logic;
signal data_in_2_5 : std_logic;
signal data_in_2_0 : std_logic;
signal \c0.n17400_cascade_\ : std_logic;
signal \c0.n8_adj_2359_cascade_\ : std_logic;
signal \c0.n13450\ : std_logic;
signal \c0.data_in_frame_3_4\ : std_logic;
signal data_in_0_1 : std_logic;
signal \c0.n7_adj_2384_cascade_\ : std_logic;
signal \c0.n6_adj_2336\ : std_logic;
signal \c0.n10136\ : std_logic;
signal data_in_1_4 : std_logic;
signal data_in_2_3 : std_logic;
signal \c0.n16_adj_2361_cascade_\ : std_logic;
signal \c0.n17_adj_2362\ : std_logic;
signal \n63_cascade_\ : std_logic;
signal data_in_2_7 : std_logic;
signal \c0.n10141\ : std_logic;
signal \c0.n10027\ : std_logic;
signal \c0.n17_adj_2370\ : std_logic;
signal \c0.n16_adj_2366_cascade_\ : std_logic;
signal data_in_1_7 : std_logic;
signal \n9378_cascade_\ : std_logic;
signal \c0.n47_adj_2347_cascade_\ : std_logic;
signal \c0.n13146_cascade_\ : std_logic;
signal data_in_3_4 : std_logic;
signal data_in_1_6 : std_logic;
signal data_in_3_5 : std_logic;
signal \c0.n17402\ : std_logic;
signal \c0.FRAME_MATCHER_state_20\ : std_logic;
signal \c0.n8_adj_2327\ : std_logic;
signal \c0.FRAME_MATCHER_i_31\ : std_logic;
signal \c0.n10161\ : std_logic;
signal \n2061_cascade_\ : std_logic;
signal \c0.n47_adj_2347\ : std_logic;
signal \c0.n9334_cascade_\ : std_logic;
signal \c0.n4\ : std_logic;
signal \c0.n15821_cascade_\ : std_logic;
signal \c0.n8_adj_2335\ : std_logic;
signal rand_data_0 : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal rand_data_1 : std_logic;
signal n16010 : std_logic;
signal rand_data_2 : std_logic;
signal n16011 : std_logic;
signal rand_data_3 : std_logic;
signal n16012 : std_logic;
signal rand_data_4 : std_logic;
signal n16013 : std_logic;
signal rand_data_5 : std_logic;
signal n16014 : std_logic;
signal rand_data_6 : std_logic;
signal n16015 : std_logic;
signal rand_data_7 : std_logic;
signal n16016 : std_logic;
signal n16017 : std_logic;
signal rand_data_8 : std_logic;
signal \bfn_10_26_0_\ : std_logic;
signal rand_data_9 : std_logic;
signal rand_setpoint_9 : std_logic;
signal n16018 : std_logic;
signal rand_data_10 : std_logic;
signal n16019 : std_logic;
signal rand_data_11 : std_logic;
signal n16020 : std_logic;
signal rand_data_12 : std_logic;
signal n16021 : std_logic;
signal rand_data_13 : std_logic;
signal n16022 : std_logic;
signal rand_data_14 : std_logic;
signal n16023 : std_logic;
signal rand_data_15 : std_logic;
signal n16024 : std_logic;
signal n16025 : std_logic;
signal rand_data_16 : std_logic;
signal \bfn_10_27_0_\ : std_logic;
signal rand_data_17 : std_logic;
signal rand_setpoint_17 : std_logic;
signal n16026 : std_logic;
signal rand_data_18 : std_logic;
signal n16027 : std_logic;
signal rand_data_19 : std_logic;
signal n16028 : std_logic;
signal rand_data_20 : std_logic;
signal n16029 : std_logic;
signal rand_data_21 : std_logic;
signal n16030 : std_logic;
signal rand_data_22 : std_logic;
signal n16031 : std_logic;
signal rand_data_23 : std_logic;
signal n16032 : std_logic;
signal n16033 : std_logic;
signal rand_data_24 : std_logic;
signal rand_setpoint_24 : std_logic;
signal \bfn_10_28_0_\ : std_logic;
signal rand_data_25 : std_logic;
signal n16034 : std_logic;
signal rand_data_26 : std_logic;
signal n16035 : std_logic;
signal rand_data_27 : std_logic;
signal n16036 : std_logic;
signal rand_data_28 : std_logic;
signal n16037 : std_logic;
signal rand_data_29 : std_logic;
signal n16038 : std_logic;
signal rand_data_30 : std_logic;
signal n16039 : std_logic;
signal rand_data_31 : std_logic;
signal n16040 : std_logic;
signal rand_setpoint_31 : std_logic;
signal rand_setpoint_26 : std_logic;
signal rand_setpoint_29 : std_logic;
signal rand_setpoint_27 : std_logic;
signal rand_setpoint_28 : std_logic;
signal rand_setpoint_11 : std_logic;
signal \c0.n17585\ : std_logic;
signal rand_setpoint_10 : std_logic;
signal \c0.n17583_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.n17022\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \c0.rx.n17058\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.n17080\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.n17710\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.n4_adj_2154\ : std_logic;
signal \c0.n4_adj_2345\ : std_logic;
signal \c0.n2122_cascade_\ : std_logic;
signal \c0.data_in_frame_2_5\ : std_logic;
signal \c0.data_in_frame_5_6\ : std_logic;
signal \c0.n2124_cascade_\ : std_logic;
signal \c0.data_in_frame_5_3\ : std_logic;
signal \c0.n16475\ : std_logic;
signal \c0.data_in_frame_5_5\ : std_logic;
signal \c0.n17373\ : std_logic;
signal \c0.n19_adj_2303\ : std_logic;
signal \c0.n17076_cascade_\ : std_logic;
signal n17075 : std_logic;
signal data_in_frame_6_4 : std_logic;
signal \c0.n10215\ : std_logic;
signal \c0.data_in_frame_0_4\ : std_logic;
signal \c0.n10215_cascade_\ : std_logic;
signal \c0.n17206_cascade_\ : std_logic;
signal \c0.n20_adj_2195\ : std_logic;
signal \c0.n39\ : std_logic;
signal \c0.n2137\ : std_logic;
signal \c0.n23_cascade_\ : std_logic;
signal \c0.n26_adj_2210\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n30_adj_2213_cascade_\ : std_logic;
signal \c0.n17_adj_2214\ : std_logic;
signal \n31_adj_2415_cascade_\ : std_logic;
signal data_in_frame_6_3 : std_logic;
signal data_in_3_7 : std_logic;
signal \c0.n6_adj_2358\ : std_logic;
signal \c0.FRAME_MATCHER_i_1\ : std_logic;
signal \c0.n15164\ : std_logic;
signal \c0.n17072_cascade_\ : std_logic;
signal \c0.data_in_frame_2_4\ : std_logic;
signal \FRAME_MATCHER_i_31__N_1273_cascade_\ : std_logic;
signal \n17086_cascade_\ : std_logic;
signal n63_adj_2428 : std_logic;
signal n63 : std_logic;
signal \c0.FRAME_MATCHER_state_8\ : std_logic;
signal \c0.n16666\ : std_logic;
signal \c0.FRAME_MATCHER_state_9\ : std_logic;
signal \c0.n16674\ : std_logic;
signal \c0.n1034\ : std_logic;
signal \n10140_cascade_\ : std_logic;
signal \c0.n8_adj_2385_cascade_\ : std_logic;
signal \c0.n16670\ : std_logic;
signal \c0.n17367_cascade_\ : std_logic;
signal \n9_cascade_\ : std_logic;
signal \c0.n10139\ : std_logic;
signal \c0.n11833\ : std_logic;
signal \c0.FRAME_MATCHER_state_3\ : std_logic;
signal \c0.FRAME_MATCHER_state_5\ : std_logic;
signal n9 : std_logic;
signal \n21_adj_2487_cascade_\ : std_logic;
signal n63_adj_2418 : std_logic;
signal n6_adj_2410 : std_logic;
signal n2061 : std_logic;
signal \c0.n51_adj_2173\ : std_logic;
signal \c0.n10166\ : std_logic;
signal \c0.FRAME_MATCHER_i_30\ : std_logic;
signal \c0.FRAME_MATCHER_i_31_N_1310_30\ : std_logic;
signal \c0.n16696\ : std_logic;
signal rand_setpoint_2 : std_logic;
signal rand_setpoint_3 : std_logic;
signal \c0.FRAME_MATCHER_state_7\ : std_logic;
signal \c0.n16141\ : std_logic;
signal rand_setpoint_23 : std_logic;
signal \c0.n17639_cascade_\ : std_logic;
signal rand_setpoint_20 : std_logic;
signal rand_setpoint_22 : std_logic;
signal \c0.n17647\ : std_logic;
signal rand_setpoint_19 : std_logic;
signal \c0.n17631_cascade_\ : std_logic;
signal rand_setpoint_18 : std_logic;
signal \c0.n17627_cascade_\ : std_logic;
signal rand_setpoint_21 : std_logic;
signal \c0.n17643\ : std_logic;
signal \c0.n18268_cascade_\ : std_logic;
signal \c0.tx.n55_cascade_\ : std_logic;
signal \c0.n5_adj_2136\ : std_logic;
signal rand_setpoint_12 : std_logic;
signal \c0.n5\ : std_logic;
signal \c0.n18172_cascade_\ : std_logic;
signal \c0.n17764\ : std_logic;
signal \c0.n17676\ : std_logic;
signal rand_setpoint_14 : std_logic;
signal \c0.n17703\ : std_logic;
signal \c0.data_out_1_4\ : std_logic;
signal \c0.n17675\ : std_logic;
signal \c0.n17697\ : std_logic;
signal n18271 : std_logic;
signal \n10_adj_2408_cascade_\ : std_logic;
signal \c0.data_out_2_3\ : std_logic;
signal data_out_0_5 : std_logic;
signal data_out_2_2 : std_logic;
signal \n2699_cascade_\ : std_logic;
signal data_out_3_4 : std_logic;
signal n2699 : std_logic;
signal data_out_3_2 : std_logic;
signal \c0.data_in_frame_2_6\ : std_logic;
signal \c0.n17713\ : std_logic;
signal \c0.n4_adj_2325\ : std_logic;
signal \c0.tx2_transmit_N_1996\ : std_logic;
signal \c0.byte_transmit_counter2_7\ : std_logic;
signal \c0.byte_transmit_counter2_6\ : std_logic;
signal \c0.n13284\ : std_logic;
signal \c0.n13628\ : std_logic;
signal \c0.n13628_cascade_\ : std_logic;
signal tx2_active : std_logic;
signal \c0.data_in_frame_3_2\ : std_logic;
signal data_in_frame_6_2 : std_logic;
signal \c0.n17475_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_5\ : std_logic;
signal \c0.n16352\ : std_logic;
signal \c0.n24_adj_2340\ : std_logic;
signal data_in_frame_6_5 : std_logic;
signal \c0.n2122\ : std_logic;
signal \c0.n17469_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_7\ : std_logic;
signal data_in_frame_6_1 : std_logic;
signal \c0.data_in_frame_5_1\ : std_logic;
signal \c0.n17114_cascade_\ : std_logic;
signal \c0.data_in_frame_5_7\ : std_logic;
signal \c0.data_in_frame_1_4\ : std_logic;
signal \c0.n17101_cascade_\ : std_logic;
signal \c0.n10_adj_2299_cascade_\ : std_logic;
signal \c0.n17206\ : std_logic;
signal \c0.n10407\ : std_logic;
signal data_in_frame_6_0 : std_logic;
signal \c0.n10407_cascade_\ : std_logic;
signal \c0.data_in_frame_1_5\ : std_logic;
signal \c0.n17215\ : std_logic;
signal \c0.n2128\ : std_logic;
signal data_in_frame_6_7 : std_logic;
signal \c0.data_in_frame_5_0\ : std_logic;
signal \c0.n2128_cascade_\ : std_logic;
signal \c0.n19_adj_2324\ : std_logic;
signal data_in_3_0 : std_logic;
signal \c0.data_in_frame_0_3\ : std_logic;
signal \c0.data_in_frame_0_2\ : std_logic;
signal \c0.n2120\ : std_logic;
signal \c0.n22_adj_2201_cascade_\ : std_logic;
signal \c0.n27_adj_2202\ : std_logic;
signal \c0.data_in_frame_0_5\ : std_logic;
signal \c0.data_in_frame_0_6\ : std_logic;
signal \c0.data_in_frame_2_0\ : std_logic;
signal data_in_3_6 : std_logic;
signal data_in_1_0 : std_logic;
signal data_in_0_0 : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_2_1 : std_logic;
signal data_in_1_1 : std_logic;
signal \c0.data_in_frame_3_5\ : std_logic;
signal \c0.data_in_frame_2_3\ : std_logic;
signal rx_data_3 : std_logic;
signal data_in_3_3 : std_logic;
signal \c0.FRAME_MATCHER_state_28\ : std_logic;
signal \c0.n50\ : std_logic;
signal \c0.n47_cascade_\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.n51\ : std_logic;
signal \c0.n56_cascade_\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.n10018_cascade_\ : std_logic;
signal n5 : std_logic;
signal n1_adj_2486 : std_logic;
signal n9378 : std_logic;
signal \FRAME_MATCHER_state_1\ : std_logic;
signal \c0.n16261\ : std_logic;
signal \c0.r_SM_Main_2_N_2034_0_adj_2167\ : std_logic;
signal \c0.n10018\ : std_logic;
signal n10088 : std_logic;
signal n17086 : std_logic;
signal n17063 : std_logic;
signal n17089 : std_logic;
signal n17090 : std_logic;
signal n3_adj_2485 : std_logic;
signal n6 : std_logic;
signal n17349 : std_logic;
signal \n3_adj_2485_cascade_\ : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_23 : std_logic;
signal blink_counter_22 : std_logic;
signal blink_counter_21 : std_logic;
signal n10140 : std_logic;
signal n8 : std_logic;
signal \n4_adj_2417_cascade_\ : std_logic;
signal \FRAME_MATCHER_state_31_N_1406_2\ : std_logic;
signal \FRAME_MATCHER_state_2\ : std_logic;
signal blink_counter_25 : std_logic;
signal n17428 : std_logic;
signal n17427 : std_logic;
signal \LED_c\ : std_logic;
signal n3779 : std_logic;
signal \FRAME_MATCHER_i_31__N_1273\ : std_logic;
signal n6_adj_2488 : std_logic;
signal data_out_3_0 : std_logic;
signal n18175 : std_logic;
signal \n10_adj_2409_cascade_\ : std_logic;
signal \c0.n8_adj_2183_cascade_\ : std_logic;
signal \c0.n17671\ : std_logic;
signal rand_setpoint_4 : std_logic;
signal \data_out_10__7__N_110_cascade_\ : std_logic;
signal rand_setpoint_6 : std_logic;
signal \c0.data_out_1_2\ : std_logic;
signal \c0.n17696\ : std_logic;
signal \n18073_cascade_\ : std_logic;
signal \c0.tx.n10688_cascade_\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal rand_setpoint_1 : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal n18070 : std_logic;
signal \c0.tx.n10688\ : std_logic;
signal \n4_adj_2419_cascade_\ : std_logic;
signal \n5_adj_2407_cascade_\ : std_logic;
signal \n10_adj_2444_cascade_\ : std_logic;
signal n8_adj_2447 : std_logic;
signal n4_adj_2419 : std_logic;
signal \bfn_12_31_0_\ : std_logic;
signal \c0.n27\ : std_logic;
signal \c0.n16066\ : std_logic;
signal \c0.n16067\ : std_logic;
signal \c0.n25_adj_2386\ : std_logic;
signal \c0.n16068\ : std_logic;
signal \c0.n16069\ : std_logic;
signal \c0.n16070\ : std_logic;
signal \c0.n22_adj_2313\ : std_logic;
signal \c0.n16071\ : std_logic;
signal \c0.n21_adj_2262\ : std_logic;
signal \c0.n16072\ : std_logic;
signal \c0.n16073\ : std_logic;
signal \bfn_12_32_0_\ : std_logic;
signal \c0.n16074\ : std_logic;
signal \c0.n16075\ : std_logic;
signal \c0.n16076\ : std_logic;
signal \c0.n16077\ : std_logic;
signal \c0.n16078\ : std_logic;
signal \c0.n10594\ : std_logic;
signal \c0.n16353\ : std_logic;
signal \c0.n26_adj_2368\ : std_logic;
signal \c0.n16474\ : std_logic;
signal \c0.n18_adj_2360\ : std_logic;
signal rx_data_0 : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal n10010 : std_logic;
signal rx_data_5 : std_logic;
signal \c0.n24_adj_2317\ : std_logic;
signal \c0.n22_adj_2319\ : std_logic;
signal \c0.n21_adj_2323\ : std_logic;
signal \c0.FRAME_MATCHER_i_0\ : std_logic;
signal \c0.FRAME_MATCHER_i_2\ : std_logic;
signal \c0.n15171_cascade_\ : std_logic;
signal \c0.data_in_frame_1_6\ : std_logic;
signal \c0.n2124\ : std_logic;
signal data_in_frame_6_6 : std_logic;
signal \c0.n17214\ : std_logic;
signal \c0.n28_adj_2374\ : std_logic;
signal \c0.n27_adj_2381_cascade_\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n12491_cascade_\ : std_logic;
signal \c0.data_in_frame_0_1\ : std_logic;
signal \c0.n10259\ : std_logic;
signal \c0.data_in_frame_2_7\ : std_logic;
signal rx_data_2 : std_logic;
signal \c0.n15179\ : std_logic;
signal \c0.n17686\ : std_logic;
signal \c0.data_out_frame2_0_4\ : std_logic;
signal \c0.n17688\ : std_logic;
signal \c0.data_out_frame2_0_3\ : std_logic;
signal \c0.data_in_frame_3_7\ : std_logic;
signal \c0.n2126\ : std_logic;
signal \c0.data_in_frame_3_0\ : std_logic;
signal \c0.n2138\ : std_logic;
signal \c0.data_in_frame_2_1\ : std_logic;
signal \c0.data_in_frame_2_2\ : std_logic;
signal \c0.n18_adj_2316_cascade_\ : std_logic;
signal \c0.data_in_frame_0_7\ : std_logic;
signal \c0.n23_adj_2322\ : std_logic;
signal \c0.FRAME_MATCHER_state_23\ : std_logic;
signal \c0.n13381\ : std_logic;
signal \c0.FRAME_MATCHER_state_11\ : std_logic;
signal \c0.n8_adj_2333\ : std_logic;
signal data_out_frame2_8_2 : std_logic;
signal \c0.n16\ : std_logic;
signal n4_adj_2427 : std_logic;
signal n4_adj_2416 : std_logic;
signal \r_Bit_Index_1_adj_2436\ : std_logic;
signal \r_Bit_Index_2_adj_2435\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \c0.rx.n10158\ : std_logic;
signal \c0.FRAME_MATCHER_state_16\ : std_logic;
signal \c0.n48\ : std_logic;
signal \c0.FRAME_MATCHER_state_30\ : std_logic;
signal \c0.n16698\ : std_logic;
signal \c0.FRAME_MATCHER_state_27\ : std_logic;
signal \c0.n16718\ : std_logic;
signal rand_setpoint_0 : std_logic;
signal n2 : std_logic;
signal data_out_2_0 : std_logic;
signal rand_setpoint_7 : std_logic;
signal data_out_0_0 : std_logic;
signal rand_setpoint_16 : std_logic;
signal rand_setpoint_15 : std_logic;
signal n10_adj_2450 : std_logic;
signal \n10_adj_2411_cascade_\ : std_logic;
signal n5_adj_2407 : std_logic;
signal \c0.n5_adj_2141\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal \n18196_cascade_\ : std_logic;
signal n18199 : std_logic;
signal \c0.tx.n31\ : std_logic;
signal n17759 : std_logic;
signal n17664 : std_logic;
signal \c0.n18166\ : std_logic;
signal \c0.n2_adj_2145\ : std_logic;
signal \c0.n17701\ : std_logic;
signal n18169 : std_logic;
signal \c0.n453\ : std_logic;
signal n4_adj_2414 : std_logic;
signal \c0.n19\ : std_logic;
signal \n9524_cascade_\ : std_logic;
signal \c0.n16267_cascade_\ : std_logic;
signal \c0.n445\ : std_logic;
signal \c0.n23_adj_2314\ : std_logic;
signal \c0.n28\ : std_logic;
signal n17765 : std_logic;
signal \n17392_cascade_\ : std_logic;
signal n17416 : std_logic;
signal \c0.n20_adj_2255\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.n24_adj_2389_cascade_\ : std_logic;
signal n17327 : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.n26_adj_2391\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.n9453_cascade_\ : std_logic;
signal \c0.n24_adj_2342\ : std_logic;
signal \c0.delay_counter_12\ : std_logic;
signal \c0.n16_adj_2212\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.n26\ : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.n22_adj_2390\ : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal \c0.n18_adj_2220\ : std_logic;
signal \c0.delay_counter_13\ : std_logic;
signal \c0.n15_adj_2211\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \c0.delay_counter_11\ : std_logic;
signal \c0.n9453\ : std_logic;
signal \c0.n16267\ : std_logic;
signal \c0.n17_adj_2219\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.n18_adj_2388\ : std_logic;
signal \c0.n17712\ : std_logic;
signal \c0.n11867\ : std_logic;
signal \c0.byte_transmit_counter2_5\ : std_logic;
signal \c0.n4_adj_2147\ : std_logic;
signal n13116 : std_logic;
signal rx_data_6 : std_logic;
signal rx_data_1 : std_logic;
signal \c0.n17072\ : std_logic;
signal \c0.data_in_frame_3_1\ : std_logic;
signal \c0.n17472_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_6\ : std_logic;
signal rx_data_ready : std_logic;
signal data_in_3_2 : std_logic;
signal data_in_2_2 : std_logic;
signal \c0.data_in_frame_1_3\ : std_logic;
signal \c0.data_in_frame_5_4\ : std_logic;
signal \c0.data_in_frame_1_2\ : std_logic;
signal \c0.n21_adj_2357\ : std_logic;
signal \c0.data_out_frame2_0_0\ : std_logic;
signal \c0.n17490\ : std_logic;
signal \c0.n15171\ : std_logic;
signal rx_data_7 : std_logic;
signal \c0.n17076\ : std_logic;
signal \c0.n26_adj_2174\ : std_logic;
signal \c0.n17487_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_1\ : std_logic;
signal \FRAME_MATCHER_state_0\ : std_logic;
signal \c0.n12491\ : std_logic;
signal \c0.n17690_cascade_\ : std_logic;
signal \c0.data_out_frame2_0_2\ : std_logic;
signal \c0.data_in_frame_5_2\ : std_logic;
signal \c0.data_in_frame_1_0\ : std_logic;
signal \c0.data_in_frame_1_1\ : std_logic;
signal \c0.n17102\ : std_logic;
signal \c0.n5815\ : std_logic;
signal \c0.n4494\ : std_logic;
signal \c0.n5817\ : std_logic;
signal n31_adj_2415 : std_logic;
signal \c0.n18202\ : std_logic;
signal \c0.FRAME_MATCHER_state_29\ : std_logic;
signal \c0.n16658\ : std_logic;
signal \c0.FRAME_MATCHER_state_10\ : std_logic;
signal \c0.n16710\ : std_logic;
signal data_out_frame2_13_4 : std_logic;
signal data_out_frame2_9_0 : std_logic;
signal \c0.n17315\ : std_logic;
signal \c0.data_in_frame_0_0\ : std_logic;
signal \c0.data_in_frame_1_7\ : std_logic;
signal \c0.n17213\ : std_logic;
signal data_out_frame2_8_5 : std_logic;
signal data_out_frame2_6_6 : std_logic;
signal \c0.n10472\ : std_logic;
signal \c0.n15821\ : std_logic;
signal \c0.FRAME_MATCHER_state_18\ : std_logic;
signal \c0.n8_adj_2329\ : std_logic;
signal \c0.n8_adj_2385\ : std_logic;
signal \c0.n46\ : std_logic;
signal \FRAME_MATCHER_i_31__N_1272\ : std_logic;
signal n488 : std_logic;
signal \c0.n13146\ : std_logic;
signal n4408 : std_logic;
signal \c0.n276_cascade_\ : std_logic;
signal \c0.n4_adj_2135\ : std_logic;
signal \c0.n4_adj_2135_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_31\ : std_logic;
signal \c0.n16700\ : std_logic;
signal \c0.n9334\ : std_logic;
signal n44 : std_logic;
signal \c0.n17069\ : std_logic;
signal \c0.FRAME_MATCHER_state_17\ : std_logic;
signal \c0.n16704\ : std_logic;
signal \c0.n3_adj_2193\ : std_logic;
signal n10_adj_2431 : std_logic;
signal \c0.n6_adj_2221\ : std_logic;
signal \c0.n17147\ : std_logic;
signal rand_setpoint_8 : std_logic;
signal \c0.n17653\ : std_logic;
signal data_out_8_1 : std_logic;
signal \c0.n1_adj_2160\ : std_logic;
signal \c0.n18184_cascade_\ : std_logic;
signal \n18187_cascade_\ : std_logic;
signal \c0.data_out_6_6\ : std_logic;
signal \c0.n5_adj_2159\ : std_logic;
signal rand_setpoint_30 : std_logic;
signal \c0.n17698\ : std_logic;
signal \c0.n17612\ : std_logic;
signal \c0.n17626\ : std_logic;
signal n25 : std_logic;
signal n28 : std_logic;
signal \n5_adj_2448_cascade_\ : std_logic;
signal \n31_cascade_\ : std_logic;
signal n22 : std_logic;
signal n9524 : std_logic;
signal n450 : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal \c0.tx.r_Bit_Index_0\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \c0.tx.n17673_cascade_\ : std_logic;
signal \c0.n10326\ : std_logic;
signal \c0.n17126\ : std_logic;
signal \c0.n17126_cascade_\ : std_logic;
signal \c0.n17651\ : std_logic;
signal n10705 : std_logic;
signal n10_adj_2444 : std_logic;
signal \bfn_14_30_0_\ : std_logic;
signal \c0.n16110\ : std_logic;
signal \c0.n16111\ : std_logic;
signal \c0.n16112\ : std_logic;
signal \c0.n16113\ : std_logic;
signal byte_transmit_counter_5 : std_logic;
signal \c0.n16114\ : std_logic;
signal byte_transmit_counter_6 : std_logic;
signal \c0.n16115\ : std_logic;
signal byte_transmit_counter_7 : std_logic;
signal \c0.n16116\ : std_logic;
signal \c0.n68_cascade_\ : std_logic;
signal \tx_transmit_N_1947_7\ : std_logic;
signal \c0.n4650\ : std_logic;
signal \tx_transmit_N_1947_3\ : std_logic;
signal \c0.n59\ : std_logic;
signal \c0.n65\ : std_logic;
signal \tx_transmit_N_1947_4\ : std_logic;
signal \tx_transmit_N_1947_5\ : std_logic;
signal \tx_transmit_N_1947_6\ : std_logic;
signal \c0.n17404\ : std_logic;
signal \tx_transmit_N_1947_1\ : std_logic;
signal \tx_transmit_N_1947_0\ : std_logic;
signal \c0.n13662\ : std_logic;
signal \c0.n13662_cascade_\ : std_logic;
signal \tx_transmit_N_1947_2\ : std_logic;
signal \c0.n13726\ : std_logic;
signal \c0.n10815\ : std_logic;
signal data_out_0_3 : std_logic;
signal n10_adj_2483 : std_logic;
signal \c0.data_out_3_6\ : std_logic;
signal \c0.FRAME_MATCHER_state_25\ : std_logic;
signal \c0.n16690\ : std_logic;
signal \c0.FRAME_MATCHER_state_26\ : std_logic;
signal \c0.n16702\ : std_logic;
signal \c0.FRAME_MATCHER_state_15\ : std_logic;
signal \c0.n8_adj_2330\ : std_logic;
signal \c0.FRAME_MATCHER_state_21\ : std_logic;
signal \c0.n16686\ : std_logic;
signal \c0.FRAME_MATCHER_state_24\ : std_logic;
signal \c0.n16688\ : std_logic;
signal \c0.n15_adj_2177\ : std_logic;
signal \c0.n17270\ : std_logic;
signal \c0.data_out_7_2\ : std_logic;
signal \c0.n10316\ : std_logic;
signal \c0.n17201\ : std_logic;
signal \c0.n10316_cascade_\ : std_logic;
signal \c0.n17177\ : std_logic;
signal data_out_8_6 : std_logic;
signal \c0.data_out_6__1__N_537\ : std_logic;
signal \c0.data_out_7_7\ : std_logic;
signal rand_setpoint_5 : std_logic;
signal n2594 : std_logic;
signal rand_setpoint_13 : std_logic;
signal \c0.data_out_7_5\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \c0.data_out_1_1\ : std_logic;
signal data_out_0_1 : std_logic;
signal n1_adj_2449 : std_logic;
signal \c0.n12630\ : std_logic;
signal \c0.data_out_7_0\ : std_logic;
signal \c0.n10395\ : std_logic;
signal \c0.n10_adj_2189_cascade_\ : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal \c0.n8_adj_2157\ : std_logic;
signal n10_adj_2422 : std_logic;
signal \c0.tx.n77_cascade_\ : std_logic;
signal \c0.tx.n12\ : std_logic;
signal tx_o : std_logic;
signal \c0.tx.n10\ : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal n10_adj_2443 : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \c0.tx.n12_adj_2134\ : std_logic;
signal \c0.n8_cascade_\ : std_logic;
signal n9257 : std_logic;
signal \c0.n65_adj_2192\ : std_logic;
signal \c0.tx.r_SM_Main_0\ : std_logic;
signal \c0.tx.n83\ : std_logic;
signal \n5142_cascade_\ : std_logic;
signal \c0.tx.n6759\ : std_logic;
signal \c0.tx.n13702\ : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \c0.data_out_5_5\ : std_logic;
signal \c0.n5_adj_2163\ : std_logic;
signal \c0.n17581_cascade_\ : std_logic;
signal n10_adj_2432 : std_logic;
signal \c0.tx.r_SM_Main_1\ : std_logic;
signal \c0.tx.n10613\ : std_logic;
signal \c0.n17622\ : std_logic;
signal \c0.n18088\ : std_logic;
signal \c0.n2_adj_2164_cascade_\ : std_logic;
signal n18091 : std_logic;
signal data_out_3_5 : std_logic;
signal \c0.data_out_0_6\ : std_logic;
signal n4 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n9999 : std_logic;
signal rx_data_4 : std_logic;
signal data_out_1_6 : std_logic;
signal \c0.n9369\ : std_logic;
signal \c0.n276\ : std_logic;
signal \FRAME_MATCHER_i_31__N_1275\ : std_logic;
signal \c0.FRAME_MATCHER_state_22\ : std_logic;
signal \c0.n16714\ : std_logic;
signal data_out_1_7 : std_logic;
signal \c0.n8_adj_2352\ : std_logic;
signal \c0.n10179\ : std_logic;
signal \c0.n10188\ : std_logic;
signal \c0.n17209_cascade_\ : std_logic;
signal \c0.data_out_10_2\ : std_logic;
signal \c0.n6_adj_2216\ : std_logic;
signal \c0.data_out_9_6\ : std_logic;
signal \c0.n17200\ : std_logic;
signal \c0.data_out_8_0\ : std_logic;
signal n8_adj_2445 : std_logic;
signal n6_adj_2446 : std_logic;
signal n23 : std_logic;
signal n32 : std_logic;
signal \n29_cascade_\ : std_logic;
signal n26 : std_logic;
signal \c0.data_out_5_2\ : std_logic;
signal \c0.n10196\ : std_logic;
signal \c0.n10196_cascade_\ : std_logic;
signal \c0.data_out_10_3\ : std_logic;
signal \c0.data_out_6_4\ : std_logic;
signal data_out_8_5 : std_logic;
signal \c0.n10392\ : std_logic;
signal \bfn_16_28_0_\ : std_logic;
signal \c0.tx.n16117\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal n10954 : std_logic;
signal \c0.tx.n16118\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal n10957 : std_logic;
signal \c0.tx.n16119\ : std_logic;
signal \c0.tx.n16120\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal n10963 : std_logic;
signal \c0.tx.n16121\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal n10966 : std_logic;
signal \c0.tx.n16122\ : std_logic;
signal \c0.tx.n16123\ : std_logic;
signal \c0.tx.n16124\ : std_logic;
signal \c0.tx.r_Clock_Count_8\ : std_logic;
signal \c0.tx.r_SM_Main_2\ : std_logic;
signal \bfn_16_29_0_\ : std_logic;
signal n10972 : std_logic;
signal data_out_8_7 : std_logic;
signal n10951 : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal n10969 : std_logic;
signal \c0.tx.r_Clock_Count_7\ : std_logic;
signal data_out_3_7 : std_logic;
signal data_out_2_7 : std_logic;
signal \c0.data_out_7__3__N_441\ : std_logic;
signal \c0.n1\ : std_logic;
signal \c0.n17747_cascade_\ : std_logic;
signal \c0.n2_adj_2156\ : std_logic;
signal \c0.n18220_cascade_\ : std_logic;
signal \c0.n17607\ : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal n10_adj_2413 : std_logic;
signal \n18223_cascade_\ : std_logic;
signal byte_transmit_counter_2 : std_logic;
signal n10 : std_logic;
signal n10960 : std_logic;
signal \c0.tx.r_Clock_Count_4\ : std_logic;
signal n10994 : std_logic;
signal n5142 : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal \c0.n10595\ : std_logic;
signal \c0.data_out_6_0\ : std_logic;
signal \c0.n17129\ : std_logic;
signal \c0.n10447_cascade_\ : std_logic;
signal \c0.data_out_6_1\ : std_logic;
signal \c0.n10183\ : std_logic;
signal \c0.data_out_6_3\ : std_logic;
signal \c0.n17222\ : std_logic;
signal \c0.data_out_9_7\ : std_logic;
signal \c0.n17243\ : std_logic;
signal \c0.n17264\ : std_logic;
signal \c0.n10_adj_2191_cascade_\ : std_logic;
signal byte_transmit_counter_0 : std_logic;
signal \c0.data_out_10_4\ : std_logic;
signal \c0.n8_adj_2198_cascade_\ : std_logic;
signal byte_transmit_counter_1 : std_logic;
signal n10_adj_2430 : std_logic;
signal \c0.n17209\ : std_logic;
signal \c0.n17297\ : std_logic;
signal \c0.n17297_cascade_\ : std_logic;
signal \c0.data_out_7__2__N_447\ : std_logic;
signal \c0.n14_adj_2176\ : std_logic;
signal \c0.data_out_7_6\ : std_logic;
signal \c0.n12_adj_2180\ : std_logic;
signal data_out_10_0 : std_logic;
signal \c0.data_out_7_3\ : std_logic;
signal \c0.data_out_5_3\ : std_logic;
signal \c0.n17180\ : std_logic;
signal \c0.data_out_9_4\ : std_logic;
signal \c0.n17162_cascade_\ : std_logic;
signal \c0.data_out_6_2\ : std_logic;
signal \c0.n17197\ : std_logic;
signal \c0.n10_adj_2196_cascade_\ : std_logic;
signal \c0.n17261\ : std_logic;
signal \c0.data_out_6_7\ : std_logic;
signal \c0.n26_adj_2165\ : std_logic;
signal \c0.data_out_6_5\ : std_logic;
signal data_out_8_3 : std_logic;
signal \c0.n10_adj_2166_cascade_\ : std_logic;
signal \c0.n10170\ : std_logic;
signal \c0.n17252\ : std_logic;
signal data_out_10_1 : std_logic;
signal data_out_8_2 : std_logic;
signal \c0.data_out_10_5\ : std_logic;
signal \c0.data_out_7_1\ : std_logic;
signal \c0.data_out_9_0\ : std_logic;
signal \c0.n6_adj_2169\ : std_logic;
signal \c0.n17162\ : std_logic;
signal \c0.n17150_cascade_\ : std_logic;
signal \c0.data_out_9_1\ : std_logic;
signal \c0.data_out_9_5\ : std_logic;
signal \c0.n17110\ : std_logic;
signal data_out_8_4 : std_logic;
signal \c0.data_out_10_7\ : std_logic;
signal \UART_TRANSMITTER_state_2\ : std_logic;
signal \UART_TRANSMITTER_state_0\ : std_logic;
signal rand_setpoint_25 : std_logic;
signal data_out_5_1 : std_logic;
signal \c0.r_SM_Main_2_N_2034_0\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal n444 : std_logic;
signal n10596 : std_logic;
signal \UART_TRANSMITTER_state_1\ : std_logic;
signal data_out_2_5 : std_logic;
signal \data_out_10__7__N_110\ : std_logic;
signal \data_out_9__2__N_367\ : std_logic;
signal \CLK_c\ : std_logic;
signal data_out_9_2 : std_logic;
signal \c0.data_out_5_4\ : std_logic;
signal \c0.data_out_10_6\ : std_logic;
signal \c0.data_out_9_3\ : std_logic;
signal \c0.n10204_cascade_\ : std_logic;
signal \c0.data_out_7_4\ : std_logic;
signal \c0.n10_adj_2172\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50887\,
            DIN => \N__50886\,
            DOUT => \N__50885\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50887\,
            PADOUT => \N__50886\,
            PADIN => \N__50885\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35976\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50878\,
            DIN => \N__50877\,
            DOUT => \N__50876\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50878\,
            PADOUT => \N__50877\,
            PADIN => \N__50876\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50869\,
            DIN => \N__50868\,
            DOUT => \N__50867\,
            PACKAGEPIN => PIN_2
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50869\,
            PADOUT => \N__50868\,
            PADIN => \N__50867\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__49762\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50860\,
            DIN => \N__50859\,
            DOUT => \N__50858\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50860\,
            PADOUT => \N__50859\,
            PADIN => \N__50858\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22131\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__17694\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50851\,
            DIN => \N__50850\,
            DOUT => \N__50849\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50851\,
            PADOUT => \N__50850\,
            PADIN => \N__50849\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__43887\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__25689\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50842\,
            DIN => \N__50841\,
            DOUT => \N__50840\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50842\,
            PADOUT => \N__50841\,
            PADIN => \N__50840\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__12827\ : InMux
    port map (
            O => \N__50823\,
            I => \N__50820\
        );

    \I__12826\ : LocalMux
    port map (
            O => \N__50820\,
            I => \N__50813\
        );

    \I__12825\ : InMux
    port map (
            O => \N__50819\,
            I => \N__50808\
        );

    \I__12824\ : InMux
    port map (
            O => \N__50818\,
            I => \N__50808\
        );

    \I__12823\ : InMux
    port map (
            O => \N__50817\,
            I => \N__50805\
        );

    \I__12822\ : InMux
    port map (
            O => \N__50816\,
            I => \N__50802\
        );

    \I__12821\ : Span4Mux_v
    port map (
            O => \N__50813\,
            I => \N__50799\
        );

    \I__12820\ : LocalMux
    port map (
            O => \N__50808\,
            I => \N__50796\
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__50805\,
            I => \N__50793\
        );

    \I__12818\ : LocalMux
    port map (
            O => \N__50802\,
            I => \N__50790\
        );

    \I__12817\ : Odrv4
    port map (
            O => \N__50799\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__12816\ : Odrv4
    port map (
            O => \N__50796\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__12815\ : Odrv4
    port map (
            O => \N__50793\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__12814\ : Odrv4
    port map (
            O => \N__50790\,
            I => \c0.r_SM_Main_2_N_2034_0\
        );

    \I__12813\ : CascadeMux
    port map (
            O => \N__50781\,
            I => \N__50777\
        );

    \I__12812\ : InMux
    port map (
            O => \N__50780\,
            I => \N__50774\
        );

    \I__12811\ : InMux
    port map (
            O => \N__50777\,
            I => \N__50770\
        );

    \I__12810\ : LocalMux
    port map (
            O => \N__50774\,
            I => \N__50767\
        );

    \I__12809\ : InMux
    port map (
            O => \N__50773\,
            I => \N__50764\
        );

    \I__12808\ : LocalMux
    port map (
            O => \N__50770\,
            I => \N__50755\
        );

    \I__12807\ : Span4Mux_v
    port map (
            O => \N__50767\,
            I => \N__50755\
        );

    \I__12806\ : LocalMux
    port map (
            O => \N__50764\,
            I => \N__50755\
        );

    \I__12805\ : InMux
    port map (
            O => \N__50763\,
            I => \N__50750\
        );

    \I__12804\ : InMux
    port map (
            O => \N__50762\,
            I => \N__50750\
        );

    \I__12803\ : Odrv4
    port map (
            O => \N__50755\,
            I => \c0.tx_active\
        );

    \I__12802\ : LocalMux
    port map (
            O => \N__50750\,
            I => \c0.tx_active\
        );

    \I__12801\ : CascadeMux
    port map (
            O => \N__50745\,
            I => \N__50737\
        );

    \I__12800\ : CascadeMux
    port map (
            O => \N__50744\,
            I => \N__50734\
        );

    \I__12799\ : CascadeMux
    port map (
            O => \N__50743\,
            I => \N__50730\
        );

    \I__12798\ : CascadeMux
    port map (
            O => \N__50742\,
            I => \N__50727\
        );

    \I__12797\ : CascadeMux
    port map (
            O => \N__50741\,
            I => \N__50724\
        );

    \I__12796\ : InMux
    port map (
            O => \N__50740\,
            I => \N__50710\
        );

    \I__12795\ : InMux
    port map (
            O => \N__50737\,
            I => \N__50710\
        );

    \I__12794\ : InMux
    port map (
            O => \N__50734\,
            I => \N__50710\
        );

    \I__12793\ : InMux
    port map (
            O => \N__50733\,
            I => \N__50707\
        );

    \I__12792\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50700\
        );

    \I__12791\ : InMux
    port map (
            O => \N__50727\,
            I => \N__50700\
        );

    \I__12790\ : InMux
    port map (
            O => \N__50724\,
            I => \N__50700\
        );

    \I__12789\ : CascadeMux
    port map (
            O => \N__50723\,
            I => \N__50695\
        );

    \I__12788\ : CascadeMux
    port map (
            O => \N__50722\,
            I => \N__50692\
        );

    \I__12787\ : CascadeMux
    port map (
            O => \N__50721\,
            I => \N__50689\
        );

    \I__12786\ : CascadeMux
    port map (
            O => \N__50720\,
            I => \N__50685\
        );

    \I__12785\ : InMux
    port map (
            O => \N__50719\,
            I => \N__50681\
        );

    \I__12784\ : InMux
    port map (
            O => \N__50718\,
            I => \N__50678\
        );

    \I__12783\ : CascadeMux
    port map (
            O => \N__50717\,
            I => \N__50673\
        );

    \I__12782\ : LocalMux
    port map (
            O => \N__50710\,
            I => \N__50670\
        );

    \I__12781\ : LocalMux
    port map (
            O => \N__50707\,
            I => \N__50667\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__50700\,
            I => \N__50664\
        );

    \I__12779\ : InMux
    port map (
            O => \N__50699\,
            I => \N__50657\
        );

    \I__12778\ : InMux
    port map (
            O => \N__50698\,
            I => \N__50657\
        );

    \I__12777\ : InMux
    port map (
            O => \N__50695\,
            I => \N__50657\
        );

    \I__12776\ : InMux
    port map (
            O => \N__50692\,
            I => \N__50654\
        );

    \I__12775\ : InMux
    port map (
            O => \N__50689\,
            I => \N__50649\
        );

    \I__12774\ : InMux
    port map (
            O => \N__50688\,
            I => \N__50649\
        );

    \I__12773\ : InMux
    port map (
            O => \N__50685\,
            I => \N__50646\
        );

    \I__12772\ : InMux
    port map (
            O => \N__50684\,
            I => \N__50643\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__50681\,
            I => \N__50638\
        );

    \I__12770\ : LocalMux
    port map (
            O => \N__50678\,
            I => \N__50638\
        );

    \I__12769\ : InMux
    port map (
            O => \N__50677\,
            I => \N__50631\
        );

    \I__12768\ : InMux
    port map (
            O => \N__50676\,
            I => \N__50631\
        );

    \I__12767\ : InMux
    port map (
            O => \N__50673\,
            I => \N__50631\
        );

    \I__12766\ : Span4Mux_s2_v
    port map (
            O => \N__50670\,
            I => \N__50622\
        );

    \I__12765\ : Span4Mux_v
    port map (
            O => \N__50667\,
            I => \N__50622\
        );

    \I__12764\ : Span4Mux_h
    port map (
            O => \N__50664\,
            I => \N__50622\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__50657\,
            I => \N__50622\
        );

    \I__12762\ : LocalMux
    port map (
            O => \N__50654\,
            I => \N__50617\
        );

    \I__12761\ : LocalMux
    port map (
            O => \N__50649\,
            I => \N__50617\
        );

    \I__12760\ : LocalMux
    port map (
            O => \N__50646\,
            I => \N__50612\
        );

    \I__12759\ : LocalMux
    port map (
            O => \N__50643\,
            I => \N__50612\
        );

    \I__12758\ : Span4Mux_v
    port map (
            O => \N__50638\,
            I => \N__50607\
        );

    \I__12757\ : LocalMux
    port map (
            O => \N__50631\,
            I => \N__50607\
        );

    \I__12756\ : Span4Mux_h
    port map (
            O => \N__50622\,
            I => \N__50604\
        );

    \I__12755\ : Span12Mux_h
    port map (
            O => \N__50617\,
            I => \N__50601\
        );

    \I__12754\ : Span4Mux_h
    port map (
            O => \N__50612\,
            I => \N__50596\
        );

    \I__12753\ : Span4Mux_h
    port map (
            O => \N__50607\,
            I => \N__50596\
        );

    \I__12752\ : Odrv4
    port map (
            O => \N__50604\,
            I => n444
        );

    \I__12751\ : Odrv12
    port map (
            O => \N__50601\,
            I => n444
        );

    \I__12750\ : Odrv4
    port map (
            O => \N__50596\,
            I => n444
        );

    \I__12749\ : CEMux
    port map (
            O => \N__50589\,
            I => \N__50584\
        );

    \I__12748\ : CEMux
    port map (
            O => \N__50588\,
            I => \N__50580\
        );

    \I__12747\ : CascadeMux
    port map (
            O => \N__50587\,
            I => \N__50577\
        );

    \I__12746\ : LocalMux
    port map (
            O => \N__50584\,
            I => \N__50571\
        );

    \I__12745\ : CascadeMux
    port map (
            O => \N__50583\,
            I => \N__50568\
        );

    \I__12744\ : LocalMux
    port map (
            O => \N__50580\,
            I => \N__50563\
        );

    \I__12743\ : InMux
    port map (
            O => \N__50577\,
            I => \N__50560\
        );

    \I__12742\ : CascadeMux
    port map (
            O => \N__50576\,
            I => \N__50557\
        );

    \I__12741\ : CEMux
    port map (
            O => \N__50575\,
            I => \N__50549\
        );

    \I__12740\ : CascadeMux
    port map (
            O => \N__50574\,
            I => \N__50543\
        );

    \I__12739\ : Span4Mux_s3_h
    port map (
            O => \N__50571\,
            I => \N__50538\
        );

    \I__12738\ : InMux
    port map (
            O => \N__50568\,
            I => \N__50534\
        );

    \I__12737\ : CEMux
    port map (
            O => \N__50567\,
            I => \N__50530\
        );

    \I__12736\ : CEMux
    port map (
            O => \N__50566\,
            I => \N__50526\
        );

    \I__12735\ : Span4Mux_v
    port map (
            O => \N__50563\,
            I => \N__50521\
        );

    \I__12734\ : LocalMux
    port map (
            O => \N__50560\,
            I => \N__50521\
        );

    \I__12733\ : InMux
    port map (
            O => \N__50557\,
            I => \N__50518\
        );

    \I__12732\ : InMux
    port map (
            O => \N__50556\,
            I => \N__50511\
        );

    \I__12731\ : InMux
    port map (
            O => \N__50555\,
            I => \N__50511\
        );

    \I__12730\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50511\
        );

    \I__12729\ : InMux
    port map (
            O => \N__50553\,
            I => \N__50506\
        );

    \I__12728\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50506\
        );

    \I__12727\ : LocalMux
    port map (
            O => \N__50549\,
            I => \N__50502\
        );

    \I__12726\ : CEMux
    port map (
            O => \N__50548\,
            I => \N__50499\
        );

    \I__12725\ : CascadeMux
    port map (
            O => \N__50547\,
            I => \N__50496\
        );

    \I__12724\ : CascadeMux
    port map (
            O => \N__50546\,
            I => \N__50493\
        );

    \I__12723\ : InMux
    port map (
            O => \N__50543\,
            I => \N__50484\
        );

    \I__12722\ : InMux
    port map (
            O => \N__50542\,
            I => \N__50484\
        );

    \I__12721\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50484\
        );

    \I__12720\ : Span4Mux_h
    port map (
            O => \N__50538\,
            I => \N__50481\
        );

    \I__12719\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50478\
        );

    \I__12718\ : LocalMux
    port map (
            O => \N__50534\,
            I => \N__50475\
        );

    \I__12717\ : InMux
    port map (
            O => \N__50533\,
            I => \N__50472\
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__50530\,
            I => \N__50467\
        );

    \I__12715\ : CascadeMux
    port map (
            O => \N__50529\,
            I => \N__50464\
        );

    \I__12714\ : LocalMux
    port map (
            O => \N__50526\,
            I => \N__50457\
        );

    \I__12713\ : Span4Mux_h
    port map (
            O => \N__50521\,
            I => \N__50457\
        );

    \I__12712\ : LocalMux
    port map (
            O => \N__50518\,
            I => \N__50457\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__50511\,
            I => \N__50452\
        );

    \I__12710\ : LocalMux
    port map (
            O => \N__50506\,
            I => \N__50452\
        );

    \I__12709\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50449\
        );

    \I__12708\ : Span4Mux_v
    port map (
            O => \N__50502\,
            I => \N__50446\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__50499\,
            I => \N__50443\
        );

    \I__12706\ : InMux
    port map (
            O => \N__50496\,
            I => \N__50436\
        );

    \I__12705\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50436\
        );

    \I__12704\ : InMux
    port map (
            O => \N__50492\,
            I => \N__50436\
        );

    \I__12703\ : CEMux
    port map (
            O => \N__50491\,
            I => \N__50433\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__50484\,
            I => \N__50430\
        );

    \I__12701\ : Span4Mux_h
    port map (
            O => \N__50481\,
            I => \N__50427\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__50478\,
            I => \N__50424\
        );

    \I__12699\ : Span4Mux_v
    port map (
            O => \N__50475\,
            I => \N__50419\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__50472\,
            I => \N__50419\
        );

    \I__12697\ : CascadeMux
    port map (
            O => \N__50471\,
            I => \N__50415\
        );

    \I__12696\ : CascadeMux
    port map (
            O => \N__50470\,
            I => \N__50412\
        );

    \I__12695\ : Span4Mux_v
    port map (
            O => \N__50467\,
            I => \N__50408\
        );

    \I__12694\ : InMux
    port map (
            O => \N__50464\,
            I => \N__50405\
        );

    \I__12693\ : Span4Mux_v
    port map (
            O => \N__50457\,
            I => \N__50398\
        );

    \I__12692\ : Span4Mux_s1_v
    port map (
            O => \N__50452\,
            I => \N__50398\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__50449\,
            I => \N__50398\
        );

    \I__12690\ : Span4Mux_h
    port map (
            O => \N__50446\,
            I => \N__50391\
        );

    \I__12689\ : Span4Mux_v
    port map (
            O => \N__50443\,
            I => \N__50391\
        );

    \I__12688\ : LocalMux
    port map (
            O => \N__50436\,
            I => \N__50391\
        );

    \I__12687\ : LocalMux
    port map (
            O => \N__50433\,
            I => \N__50387\
        );

    \I__12686\ : Span12Mux_v
    port map (
            O => \N__50430\,
            I => \N__50384\
        );

    \I__12685\ : Span4Mux_h
    port map (
            O => \N__50427\,
            I => \N__50377\
        );

    \I__12684\ : Span4Mux_v
    port map (
            O => \N__50424\,
            I => \N__50377\
        );

    \I__12683\ : Span4Mux_v
    port map (
            O => \N__50419\,
            I => \N__50377\
        );

    \I__12682\ : InMux
    port map (
            O => \N__50418\,
            I => \N__50372\
        );

    \I__12681\ : InMux
    port map (
            O => \N__50415\,
            I => \N__50372\
        );

    \I__12680\ : InMux
    port map (
            O => \N__50412\,
            I => \N__50369\
        );

    \I__12679\ : InMux
    port map (
            O => \N__50411\,
            I => \N__50366\
        );

    \I__12678\ : Span4Mux_v
    port map (
            O => \N__50408\,
            I => \N__50357\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__50405\,
            I => \N__50357\
        );

    \I__12676\ : Span4Mux_h
    port map (
            O => \N__50398\,
            I => \N__50357\
        );

    \I__12675\ : Span4Mux_s1_v
    port map (
            O => \N__50391\,
            I => \N__50357\
        );

    \I__12674\ : InMux
    port map (
            O => \N__50390\,
            I => \N__50354\
        );

    \I__12673\ : Odrv4
    port map (
            O => \N__50387\,
            I => n10596
        );

    \I__12672\ : Odrv12
    port map (
            O => \N__50384\,
            I => n10596
        );

    \I__12671\ : Odrv4
    port map (
            O => \N__50377\,
            I => n10596
        );

    \I__12670\ : LocalMux
    port map (
            O => \N__50372\,
            I => n10596
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__50369\,
            I => n10596
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__50366\,
            I => n10596
        );

    \I__12667\ : Odrv4
    port map (
            O => \N__50357\,
            I => n10596
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__50354\,
            I => n10596
        );

    \I__12665\ : InMux
    port map (
            O => \N__50337\,
            I => \N__50334\
        );

    \I__12664\ : LocalMux
    port map (
            O => \N__50334\,
            I => \N__50330\
        );

    \I__12663\ : CascadeMux
    port map (
            O => \N__50333\,
            I => \N__50325\
        );

    \I__12662\ : Span4Mux_h
    port map (
            O => \N__50330\,
            I => \N__50311\
        );

    \I__12661\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50306\
        );

    \I__12660\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50306\
        );

    \I__12659\ : InMux
    port map (
            O => \N__50325\,
            I => \N__50301\
        );

    \I__12658\ : InMux
    port map (
            O => \N__50324\,
            I => \N__50301\
        );

    \I__12657\ : InMux
    port map (
            O => \N__50323\,
            I => \N__50296\
        );

    \I__12656\ : InMux
    port map (
            O => \N__50322\,
            I => \N__50296\
        );

    \I__12655\ : CascadeMux
    port map (
            O => \N__50321\,
            I => \N__50293\
        );

    \I__12654\ : InMux
    port map (
            O => \N__50320\,
            I => \N__50287\
        );

    \I__12653\ : InMux
    port map (
            O => \N__50319\,
            I => \N__50284\
        );

    \I__12652\ : InMux
    port map (
            O => \N__50318\,
            I => \N__50281\
        );

    \I__12651\ : InMux
    port map (
            O => \N__50317\,
            I => \N__50278\
        );

    \I__12650\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50272\
        );

    \I__12649\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50267\
        );

    \I__12648\ : CascadeMux
    port map (
            O => \N__50314\,
            I => \N__50263\
        );

    \I__12647\ : Span4Mux_h
    port map (
            O => \N__50311\,
            I => \N__50254\
        );

    \I__12646\ : LocalMux
    port map (
            O => \N__50306\,
            I => \N__50254\
        );

    \I__12645\ : LocalMux
    port map (
            O => \N__50301\,
            I => \N__50249\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__50296\,
            I => \N__50249\
        );

    \I__12643\ : InMux
    port map (
            O => \N__50293\,
            I => \N__50245\
        );

    \I__12642\ : InMux
    port map (
            O => \N__50292\,
            I => \N__50241\
        );

    \I__12641\ : InMux
    port map (
            O => \N__50291\,
            I => \N__50238\
        );

    \I__12640\ : InMux
    port map (
            O => \N__50290\,
            I => \N__50233\
        );

    \I__12639\ : LocalMux
    port map (
            O => \N__50287\,
            I => \N__50230\
        );

    \I__12638\ : LocalMux
    port map (
            O => \N__50284\,
            I => \N__50227\
        );

    \I__12637\ : LocalMux
    port map (
            O => \N__50281\,
            I => \N__50222\
        );

    \I__12636\ : LocalMux
    port map (
            O => \N__50278\,
            I => \N__50222\
        );

    \I__12635\ : InMux
    port map (
            O => \N__50277\,
            I => \N__50215\
        );

    \I__12634\ : InMux
    port map (
            O => \N__50276\,
            I => \N__50215\
        );

    \I__12633\ : InMux
    port map (
            O => \N__50275\,
            I => \N__50215\
        );

    \I__12632\ : LocalMux
    port map (
            O => \N__50272\,
            I => \N__50212\
        );

    \I__12631\ : InMux
    port map (
            O => \N__50271\,
            I => \N__50207\
        );

    \I__12630\ : InMux
    port map (
            O => \N__50270\,
            I => \N__50207\
        );

    \I__12629\ : LocalMux
    port map (
            O => \N__50267\,
            I => \N__50201\
        );

    \I__12628\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50198\
        );

    \I__12627\ : InMux
    port map (
            O => \N__50263\,
            I => \N__50195\
        );

    \I__12626\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50192\
        );

    \I__12625\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50187\
        );

    \I__12624\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50187\
        );

    \I__12623\ : InMux
    port map (
            O => \N__50259\,
            I => \N__50184\
        );

    \I__12622\ : Span4Mux_h
    port map (
            O => \N__50254\,
            I => \N__50179\
        );

    \I__12621\ : Span4Mux_h
    port map (
            O => \N__50249\,
            I => \N__50179\
        );

    \I__12620\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50176\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__50245\,
            I => \N__50173\
        );

    \I__12618\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50170\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__50241\,
            I => \N__50165\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__50238\,
            I => \N__50165\
        );

    \I__12615\ : InMux
    port map (
            O => \N__50237\,
            I => \N__50162\
        );

    \I__12614\ : InMux
    port map (
            O => \N__50236\,
            I => \N__50159\
        );

    \I__12613\ : LocalMux
    port map (
            O => \N__50233\,
            I => \N__50147\
        );

    \I__12612\ : Span4Mux_h
    port map (
            O => \N__50230\,
            I => \N__50138\
        );

    \I__12611\ : Span4Mux_s1_v
    port map (
            O => \N__50227\,
            I => \N__50138\
        );

    \I__12610\ : Span4Mux_h
    port map (
            O => \N__50222\,
            I => \N__50138\
        );

    \I__12609\ : LocalMux
    port map (
            O => \N__50215\,
            I => \N__50138\
        );

    \I__12608\ : Span4Mux_s3_v
    port map (
            O => \N__50212\,
            I => \N__50130\
        );

    \I__12607\ : LocalMux
    port map (
            O => \N__50207\,
            I => \N__50130\
        );

    \I__12606\ : InMux
    port map (
            O => \N__50206\,
            I => \N__50125\
        );

    \I__12605\ : InMux
    port map (
            O => \N__50205\,
            I => \N__50125\
        );

    \I__12604\ : InMux
    port map (
            O => \N__50204\,
            I => \N__50122\
        );

    \I__12603\ : Span4Mux_v
    port map (
            O => \N__50201\,
            I => \N__50119\
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__50198\,
            I => \N__50116\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__50195\,
            I => \N__50111\
        );

    \I__12600\ : LocalMux
    port map (
            O => \N__50192\,
            I => \N__50111\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__50187\,
            I => \N__50108\
        );

    \I__12598\ : LocalMux
    port map (
            O => \N__50184\,
            I => \N__50105\
        );

    \I__12597\ : IoSpan4Mux
    port map (
            O => \N__50179\,
            I => \N__50100\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__50176\,
            I => \N__50100\
        );

    \I__12595\ : Span4Mux_v
    port map (
            O => \N__50173\,
            I => \N__50097\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__50170\,
            I => \N__50088\
        );

    \I__12593\ : Span12Mux_v
    port map (
            O => \N__50165\,
            I => \N__50088\
        );

    \I__12592\ : LocalMux
    port map (
            O => \N__50162\,
            I => \N__50088\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__50159\,
            I => \N__50088\
        );

    \I__12590\ : InMux
    port map (
            O => \N__50158\,
            I => \N__50081\
        );

    \I__12589\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50081\
        );

    \I__12588\ : InMux
    port map (
            O => \N__50156\,
            I => \N__50081\
        );

    \I__12587\ : InMux
    port map (
            O => \N__50155\,
            I => \N__50076\
        );

    \I__12586\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50076\
        );

    \I__12585\ : InMux
    port map (
            O => \N__50153\,
            I => \N__50073\
        );

    \I__12584\ : InMux
    port map (
            O => \N__50152\,
            I => \N__50066\
        );

    \I__12583\ : InMux
    port map (
            O => \N__50151\,
            I => \N__50066\
        );

    \I__12582\ : InMux
    port map (
            O => \N__50150\,
            I => \N__50066\
        );

    \I__12581\ : Span4Mux_v
    port map (
            O => \N__50147\,
            I => \N__50061\
        );

    \I__12580\ : Span4Mux_v
    port map (
            O => \N__50138\,
            I => \N__50061\
        );

    \I__12579\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50054\
        );

    \I__12578\ : InMux
    port map (
            O => \N__50136\,
            I => \N__50054\
        );

    \I__12577\ : InMux
    port map (
            O => \N__50135\,
            I => \N__50054\
        );

    \I__12576\ : Span4Mux_h
    port map (
            O => \N__50130\,
            I => \N__50047\
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__50125\,
            I => \N__50047\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__50122\,
            I => \N__50047\
        );

    \I__12573\ : Span4Mux_h
    port map (
            O => \N__50119\,
            I => \N__50044\
        );

    \I__12572\ : Span4Mux_h
    port map (
            O => \N__50116\,
            I => \N__50033\
        );

    \I__12571\ : Span4Mux_h
    port map (
            O => \N__50111\,
            I => \N__50033\
        );

    \I__12570\ : Span4Mux_h
    port map (
            O => \N__50108\,
            I => \N__50033\
        );

    \I__12569\ : Span4Mux_h
    port map (
            O => \N__50105\,
            I => \N__50033\
        );

    \I__12568\ : Span4Mux_s2_v
    port map (
            O => \N__50100\,
            I => \N__50033\
        );

    \I__12567\ : Sp12to4
    port map (
            O => \N__50097\,
            I => \N__50028\
        );

    \I__12566\ : Span12Mux_s5_v
    port map (
            O => \N__50088\,
            I => \N__50028\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__50081\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12564\ : LocalMux
    port map (
            O => \N__50076\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12563\ : LocalMux
    port map (
            O => \N__50073\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__50066\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12561\ : Odrv4
    port map (
            O => \N__50061\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12560\ : LocalMux
    port map (
            O => \N__50054\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12559\ : Odrv4
    port map (
            O => \N__50047\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12558\ : Odrv4
    port map (
            O => \N__50044\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12557\ : Odrv4
    port map (
            O => \N__50033\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12556\ : Odrv12
    port map (
            O => \N__50028\,
            I => \UART_TRANSMITTER_state_1\
        );

    \I__12555\ : InMux
    port map (
            O => \N__50007\,
            I => \N__50004\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__50004\,
            I => \N__50000\
        );

    \I__12553\ : InMux
    port map (
            O => \N__50003\,
            I => \N__49997\
        );

    \I__12552\ : Span4Mux_s1_v
    port map (
            O => \N__50000\,
            I => \N__49994\
        );

    \I__12551\ : LocalMux
    port map (
            O => \N__49997\,
            I => data_out_2_5
        );

    \I__12550\ : Odrv4
    port map (
            O => \N__49994\,
            I => data_out_2_5
        );

    \I__12549\ : CEMux
    port map (
            O => \N__49989\,
            I => \N__49985\
        );

    \I__12548\ : CEMux
    port map (
            O => \N__49988\,
            I => \N__49981\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__49985\,
            I => \N__49974\
        );

    \I__12546\ : CEMux
    port map (
            O => \N__49984\,
            I => \N__49971\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__49981\,
            I => \N__49967\
        );

    \I__12544\ : CEMux
    port map (
            O => \N__49980\,
            I => \N__49964\
        );

    \I__12543\ : CEMux
    port map (
            O => \N__49979\,
            I => \N__49959\
        );

    \I__12542\ : InMux
    port map (
            O => \N__49978\,
            I => \N__49956\
        );

    \I__12541\ : InMux
    port map (
            O => \N__49977\,
            I => \N__49953\
        );

    \I__12540\ : Span4Mux_v
    port map (
            O => \N__49974\,
            I => \N__49950\
        );

    \I__12539\ : LocalMux
    port map (
            O => \N__49971\,
            I => \N__49947\
        );

    \I__12538\ : CEMux
    port map (
            O => \N__49970\,
            I => \N__49944\
        );

    \I__12537\ : Span4Mux_v
    port map (
            O => \N__49967\,
            I => \N__49939\
        );

    \I__12536\ : LocalMux
    port map (
            O => \N__49964\,
            I => \N__49939\
        );

    \I__12535\ : CascadeMux
    port map (
            O => \N__49963\,
            I => \N__49936\
        );

    \I__12534\ : CascadeMux
    port map (
            O => \N__49962\,
            I => \N__49931\
        );

    \I__12533\ : LocalMux
    port map (
            O => \N__49959\,
            I => \N__49924\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__49956\,
            I => \N__49924\
        );

    \I__12531\ : LocalMux
    port map (
            O => \N__49953\,
            I => \N__49921\
        );

    \I__12530\ : Span4Mux_h
    port map (
            O => \N__49950\,
            I => \N__49916\
        );

    \I__12529\ : Span4Mux_h
    port map (
            O => \N__49947\,
            I => \N__49916\
        );

    \I__12528\ : LocalMux
    port map (
            O => \N__49944\,
            I => \N__49913\
        );

    \I__12527\ : Span4Mux_h
    port map (
            O => \N__49939\,
            I => \N__49910\
        );

    \I__12526\ : InMux
    port map (
            O => \N__49936\,
            I => \N__49907\
        );

    \I__12525\ : InMux
    port map (
            O => \N__49935\,
            I => \N__49902\
        );

    \I__12524\ : InMux
    port map (
            O => \N__49934\,
            I => \N__49902\
        );

    \I__12523\ : InMux
    port map (
            O => \N__49931\,
            I => \N__49897\
        );

    \I__12522\ : InMux
    port map (
            O => \N__49930\,
            I => \N__49897\
        );

    \I__12521\ : InMux
    port map (
            O => \N__49929\,
            I => \N__49894\
        );

    \I__12520\ : Span4Mux_h
    port map (
            O => \N__49924\,
            I => \N__49889\
        );

    \I__12519\ : Span4Mux_v
    port map (
            O => \N__49921\,
            I => \N__49889\
        );

    \I__12518\ : Span4Mux_h
    port map (
            O => \N__49916\,
            I => \N__49886\
        );

    \I__12517\ : Span4Mux_h
    port map (
            O => \N__49913\,
            I => \N__49881\
        );

    \I__12516\ : Span4Mux_h
    port map (
            O => \N__49910\,
            I => \N__49881\
        );

    \I__12515\ : LocalMux
    port map (
            O => \N__49907\,
            I => \data_out_10__7__N_110\
        );

    \I__12514\ : LocalMux
    port map (
            O => \N__49902\,
            I => \data_out_10__7__N_110\
        );

    \I__12513\ : LocalMux
    port map (
            O => \N__49897\,
            I => \data_out_10__7__N_110\
        );

    \I__12512\ : LocalMux
    port map (
            O => \N__49894\,
            I => \data_out_10__7__N_110\
        );

    \I__12511\ : Odrv4
    port map (
            O => \N__49889\,
            I => \data_out_10__7__N_110\
        );

    \I__12510\ : Odrv4
    port map (
            O => \N__49886\,
            I => \data_out_10__7__N_110\
        );

    \I__12509\ : Odrv4
    port map (
            O => \N__49881\,
            I => \data_out_10__7__N_110\
        );

    \I__12508\ : InMux
    port map (
            O => \N__49866\,
            I => \N__49862\
        );

    \I__12507\ : InMux
    port map (
            O => \N__49865\,
            I => \N__49859\
        );

    \I__12506\ : LocalMux
    port map (
            O => \N__49862\,
            I => \N__49854\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__49859\,
            I => \N__49854\
        );

    \I__12504\ : Odrv4
    port map (
            O => \N__49854\,
            I => \data_out_9__2__N_367\
        );

    \I__12503\ : ClkMux
    port map (
            O => \N__49851\,
            I => \N__49176\
        );

    \I__12502\ : ClkMux
    port map (
            O => \N__49850\,
            I => \N__49176\
        );

    \I__12501\ : ClkMux
    port map (
            O => \N__49849\,
            I => \N__49176\
        );

    \I__12500\ : ClkMux
    port map (
            O => \N__49848\,
            I => \N__49176\
        );

    \I__12499\ : ClkMux
    port map (
            O => \N__49847\,
            I => \N__49176\
        );

    \I__12498\ : ClkMux
    port map (
            O => \N__49846\,
            I => \N__49176\
        );

    \I__12497\ : ClkMux
    port map (
            O => \N__49845\,
            I => \N__49176\
        );

    \I__12496\ : ClkMux
    port map (
            O => \N__49844\,
            I => \N__49176\
        );

    \I__12495\ : ClkMux
    port map (
            O => \N__49843\,
            I => \N__49176\
        );

    \I__12494\ : ClkMux
    port map (
            O => \N__49842\,
            I => \N__49176\
        );

    \I__12493\ : ClkMux
    port map (
            O => \N__49841\,
            I => \N__49176\
        );

    \I__12492\ : ClkMux
    port map (
            O => \N__49840\,
            I => \N__49176\
        );

    \I__12491\ : ClkMux
    port map (
            O => \N__49839\,
            I => \N__49176\
        );

    \I__12490\ : ClkMux
    port map (
            O => \N__49838\,
            I => \N__49176\
        );

    \I__12489\ : ClkMux
    port map (
            O => \N__49837\,
            I => \N__49176\
        );

    \I__12488\ : ClkMux
    port map (
            O => \N__49836\,
            I => \N__49176\
        );

    \I__12487\ : ClkMux
    port map (
            O => \N__49835\,
            I => \N__49176\
        );

    \I__12486\ : ClkMux
    port map (
            O => \N__49834\,
            I => \N__49176\
        );

    \I__12485\ : ClkMux
    port map (
            O => \N__49833\,
            I => \N__49176\
        );

    \I__12484\ : ClkMux
    port map (
            O => \N__49832\,
            I => \N__49176\
        );

    \I__12483\ : ClkMux
    port map (
            O => \N__49831\,
            I => \N__49176\
        );

    \I__12482\ : ClkMux
    port map (
            O => \N__49830\,
            I => \N__49176\
        );

    \I__12481\ : ClkMux
    port map (
            O => \N__49829\,
            I => \N__49176\
        );

    \I__12480\ : ClkMux
    port map (
            O => \N__49828\,
            I => \N__49176\
        );

    \I__12479\ : ClkMux
    port map (
            O => \N__49827\,
            I => \N__49176\
        );

    \I__12478\ : ClkMux
    port map (
            O => \N__49826\,
            I => \N__49176\
        );

    \I__12477\ : ClkMux
    port map (
            O => \N__49825\,
            I => \N__49176\
        );

    \I__12476\ : ClkMux
    port map (
            O => \N__49824\,
            I => \N__49176\
        );

    \I__12475\ : ClkMux
    port map (
            O => \N__49823\,
            I => \N__49176\
        );

    \I__12474\ : ClkMux
    port map (
            O => \N__49822\,
            I => \N__49176\
        );

    \I__12473\ : ClkMux
    port map (
            O => \N__49821\,
            I => \N__49176\
        );

    \I__12472\ : ClkMux
    port map (
            O => \N__49820\,
            I => \N__49176\
        );

    \I__12471\ : ClkMux
    port map (
            O => \N__49819\,
            I => \N__49176\
        );

    \I__12470\ : ClkMux
    port map (
            O => \N__49818\,
            I => \N__49176\
        );

    \I__12469\ : ClkMux
    port map (
            O => \N__49817\,
            I => \N__49176\
        );

    \I__12468\ : ClkMux
    port map (
            O => \N__49816\,
            I => \N__49176\
        );

    \I__12467\ : ClkMux
    port map (
            O => \N__49815\,
            I => \N__49176\
        );

    \I__12466\ : ClkMux
    port map (
            O => \N__49814\,
            I => \N__49176\
        );

    \I__12465\ : ClkMux
    port map (
            O => \N__49813\,
            I => \N__49176\
        );

    \I__12464\ : ClkMux
    port map (
            O => \N__49812\,
            I => \N__49176\
        );

    \I__12463\ : ClkMux
    port map (
            O => \N__49811\,
            I => \N__49176\
        );

    \I__12462\ : ClkMux
    port map (
            O => \N__49810\,
            I => \N__49176\
        );

    \I__12461\ : ClkMux
    port map (
            O => \N__49809\,
            I => \N__49176\
        );

    \I__12460\ : ClkMux
    port map (
            O => \N__49808\,
            I => \N__49176\
        );

    \I__12459\ : ClkMux
    port map (
            O => \N__49807\,
            I => \N__49176\
        );

    \I__12458\ : ClkMux
    port map (
            O => \N__49806\,
            I => \N__49176\
        );

    \I__12457\ : ClkMux
    port map (
            O => \N__49805\,
            I => \N__49176\
        );

    \I__12456\ : ClkMux
    port map (
            O => \N__49804\,
            I => \N__49176\
        );

    \I__12455\ : ClkMux
    port map (
            O => \N__49803\,
            I => \N__49176\
        );

    \I__12454\ : ClkMux
    port map (
            O => \N__49802\,
            I => \N__49176\
        );

    \I__12453\ : ClkMux
    port map (
            O => \N__49801\,
            I => \N__49176\
        );

    \I__12452\ : ClkMux
    port map (
            O => \N__49800\,
            I => \N__49176\
        );

    \I__12451\ : ClkMux
    port map (
            O => \N__49799\,
            I => \N__49176\
        );

    \I__12450\ : ClkMux
    port map (
            O => \N__49798\,
            I => \N__49176\
        );

    \I__12449\ : ClkMux
    port map (
            O => \N__49797\,
            I => \N__49176\
        );

    \I__12448\ : ClkMux
    port map (
            O => \N__49796\,
            I => \N__49176\
        );

    \I__12447\ : ClkMux
    port map (
            O => \N__49795\,
            I => \N__49176\
        );

    \I__12446\ : ClkMux
    port map (
            O => \N__49794\,
            I => \N__49176\
        );

    \I__12445\ : ClkMux
    port map (
            O => \N__49793\,
            I => \N__49176\
        );

    \I__12444\ : ClkMux
    port map (
            O => \N__49792\,
            I => \N__49176\
        );

    \I__12443\ : ClkMux
    port map (
            O => \N__49791\,
            I => \N__49176\
        );

    \I__12442\ : ClkMux
    port map (
            O => \N__49790\,
            I => \N__49176\
        );

    \I__12441\ : ClkMux
    port map (
            O => \N__49789\,
            I => \N__49176\
        );

    \I__12440\ : ClkMux
    port map (
            O => \N__49788\,
            I => \N__49176\
        );

    \I__12439\ : ClkMux
    port map (
            O => \N__49787\,
            I => \N__49176\
        );

    \I__12438\ : ClkMux
    port map (
            O => \N__49786\,
            I => \N__49176\
        );

    \I__12437\ : ClkMux
    port map (
            O => \N__49785\,
            I => \N__49176\
        );

    \I__12436\ : ClkMux
    port map (
            O => \N__49784\,
            I => \N__49176\
        );

    \I__12435\ : ClkMux
    port map (
            O => \N__49783\,
            I => \N__49176\
        );

    \I__12434\ : ClkMux
    port map (
            O => \N__49782\,
            I => \N__49176\
        );

    \I__12433\ : ClkMux
    port map (
            O => \N__49781\,
            I => \N__49176\
        );

    \I__12432\ : ClkMux
    port map (
            O => \N__49780\,
            I => \N__49176\
        );

    \I__12431\ : ClkMux
    port map (
            O => \N__49779\,
            I => \N__49176\
        );

    \I__12430\ : ClkMux
    port map (
            O => \N__49778\,
            I => \N__49176\
        );

    \I__12429\ : ClkMux
    port map (
            O => \N__49777\,
            I => \N__49176\
        );

    \I__12428\ : ClkMux
    port map (
            O => \N__49776\,
            I => \N__49176\
        );

    \I__12427\ : ClkMux
    port map (
            O => \N__49775\,
            I => \N__49176\
        );

    \I__12426\ : ClkMux
    port map (
            O => \N__49774\,
            I => \N__49176\
        );

    \I__12425\ : ClkMux
    port map (
            O => \N__49773\,
            I => \N__49176\
        );

    \I__12424\ : ClkMux
    port map (
            O => \N__49772\,
            I => \N__49176\
        );

    \I__12423\ : ClkMux
    port map (
            O => \N__49771\,
            I => \N__49176\
        );

    \I__12422\ : ClkMux
    port map (
            O => \N__49770\,
            I => \N__49176\
        );

    \I__12421\ : ClkMux
    port map (
            O => \N__49769\,
            I => \N__49176\
        );

    \I__12420\ : ClkMux
    port map (
            O => \N__49768\,
            I => \N__49176\
        );

    \I__12419\ : ClkMux
    port map (
            O => \N__49767\,
            I => \N__49176\
        );

    \I__12418\ : ClkMux
    port map (
            O => \N__49766\,
            I => \N__49176\
        );

    \I__12417\ : ClkMux
    port map (
            O => \N__49765\,
            I => \N__49176\
        );

    \I__12416\ : ClkMux
    port map (
            O => \N__49764\,
            I => \N__49176\
        );

    \I__12415\ : ClkMux
    port map (
            O => \N__49763\,
            I => \N__49176\
        );

    \I__12414\ : ClkMux
    port map (
            O => \N__49762\,
            I => \N__49176\
        );

    \I__12413\ : ClkMux
    port map (
            O => \N__49761\,
            I => \N__49176\
        );

    \I__12412\ : ClkMux
    port map (
            O => \N__49760\,
            I => \N__49176\
        );

    \I__12411\ : ClkMux
    port map (
            O => \N__49759\,
            I => \N__49176\
        );

    \I__12410\ : ClkMux
    port map (
            O => \N__49758\,
            I => \N__49176\
        );

    \I__12409\ : ClkMux
    port map (
            O => \N__49757\,
            I => \N__49176\
        );

    \I__12408\ : ClkMux
    port map (
            O => \N__49756\,
            I => \N__49176\
        );

    \I__12407\ : ClkMux
    port map (
            O => \N__49755\,
            I => \N__49176\
        );

    \I__12406\ : ClkMux
    port map (
            O => \N__49754\,
            I => \N__49176\
        );

    \I__12405\ : ClkMux
    port map (
            O => \N__49753\,
            I => \N__49176\
        );

    \I__12404\ : ClkMux
    port map (
            O => \N__49752\,
            I => \N__49176\
        );

    \I__12403\ : ClkMux
    port map (
            O => \N__49751\,
            I => \N__49176\
        );

    \I__12402\ : ClkMux
    port map (
            O => \N__49750\,
            I => \N__49176\
        );

    \I__12401\ : ClkMux
    port map (
            O => \N__49749\,
            I => \N__49176\
        );

    \I__12400\ : ClkMux
    port map (
            O => \N__49748\,
            I => \N__49176\
        );

    \I__12399\ : ClkMux
    port map (
            O => \N__49747\,
            I => \N__49176\
        );

    \I__12398\ : ClkMux
    port map (
            O => \N__49746\,
            I => \N__49176\
        );

    \I__12397\ : ClkMux
    port map (
            O => \N__49745\,
            I => \N__49176\
        );

    \I__12396\ : ClkMux
    port map (
            O => \N__49744\,
            I => \N__49176\
        );

    \I__12395\ : ClkMux
    port map (
            O => \N__49743\,
            I => \N__49176\
        );

    \I__12394\ : ClkMux
    port map (
            O => \N__49742\,
            I => \N__49176\
        );

    \I__12393\ : ClkMux
    port map (
            O => \N__49741\,
            I => \N__49176\
        );

    \I__12392\ : ClkMux
    port map (
            O => \N__49740\,
            I => \N__49176\
        );

    \I__12391\ : ClkMux
    port map (
            O => \N__49739\,
            I => \N__49176\
        );

    \I__12390\ : ClkMux
    port map (
            O => \N__49738\,
            I => \N__49176\
        );

    \I__12389\ : ClkMux
    port map (
            O => \N__49737\,
            I => \N__49176\
        );

    \I__12388\ : ClkMux
    port map (
            O => \N__49736\,
            I => \N__49176\
        );

    \I__12387\ : ClkMux
    port map (
            O => \N__49735\,
            I => \N__49176\
        );

    \I__12386\ : ClkMux
    port map (
            O => \N__49734\,
            I => \N__49176\
        );

    \I__12385\ : ClkMux
    port map (
            O => \N__49733\,
            I => \N__49176\
        );

    \I__12384\ : ClkMux
    port map (
            O => \N__49732\,
            I => \N__49176\
        );

    \I__12383\ : ClkMux
    port map (
            O => \N__49731\,
            I => \N__49176\
        );

    \I__12382\ : ClkMux
    port map (
            O => \N__49730\,
            I => \N__49176\
        );

    \I__12381\ : ClkMux
    port map (
            O => \N__49729\,
            I => \N__49176\
        );

    \I__12380\ : ClkMux
    port map (
            O => \N__49728\,
            I => \N__49176\
        );

    \I__12379\ : ClkMux
    port map (
            O => \N__49727\,
            I => \N__49176\
        );

    \I__12378\ : ClkMux
    port map (
            O => \N__49726\,
            I => \N__49176\
        );

    \I__12377\ : ClkMux
    port map (
            O => \N__49725\,
            I => \N__49176\
        );

    \I__12376\ : ClkMux
    port map (
            O => \N__49724\,
            I => \N__49176\
        );

    \I__12375\ : ClkMux
    port map (
            O => \N__49723\,
            I => \N__49176\
        );

    \I__12374\ : ClkMux
    port map (
            O => \N__49722\,
            I => \N__49176\
        );

    \I__12373\ : ClkMux
    port map (
            O => \N__49721\,
            I => \N__49176\
        );

    \I__12372\ : ClkMux
    port map (
            O => \N__49720\,
            I => \N__49176\
        );

    \I__12371\ : ClkMux
    port map (
            O => \N__49719\,
            I => \N__49176\
        );

    \I__12370\ : ClkMux
    port map (
            O => \N__49718\,
            I => \N__49176\
        );

    \I__12369\ : ClkMux
    port map (
            O => \N__49717\,
            I => \N__49176\
        );

    \I__12368\ : ClkMux
    port map (
            O => \N__49716\,
            I => \N__49176\
        );

    \I__12367\ : ClkMux
    port map (
            O => \N__49715\,
            I => \N__49176\
        );

    \I__12366\ : ClkMux
    port map (
            O => \N__49714\,
            I => \N__49176\
        );

    \I__12365\ : ClkMux
    port map (
            O => \N__49713\,
            I => \N__49176\
        );

    \I__12364\ : ClkMux
    port map (
            O => \N__49712\,
            I => \N__49176\
        );

    \I__12363\ : ClkMux
    port map (
            O => \N__49711\,
            I => \N__49176\
        );

    \I__12362\ : ClkMux
    port map (
            O => \N__49710\,
            I => \N__49176\
        );

    \I__12361\ : ClkMux
    port map (
            O => \N__49709\,
            I => \N__49176\
        );

    \I__12360\ : ClkMux
    port map (
            O => \N__49708\,
            I => \N__49176\
        );

    \I__12359\ : ClkMux
    port map (
            O => \N__49707\,
            I => \N__49176\
        );

    \I__12358\ : ClkMux
    port map (
            O => \N__49706\,
            I => \N__49176\
        );

    \I__12357\ : ClkMux
    port map (
            O => \N__49705\,
            I => \N__49176\
        );

    \I__12356\ : ClkMux
    port map (
            O => \N__49704\,
            I => \N__49176\
        );

    \I__12355\ : ClkMux
    port map (
            O => \N__49703\,
            I => \N__49176\
        );

    \I__12354\ : ClkMux
    port map (
            O => \N__49702\,
            I => \N__49176\
        );

    \I__12353\ : ClkMux
    port map (
            O => \N__49701\,
            I => \N__49176\
        );

    \I__12352\ : ClkMux
    port map (
            O => \N__49700\,
            I => \N__49176\
        );

    \I__12351\ : ClkMux
    port map (
            O => \N__49699\,
            I => \N__49176\
        );

    \I__12350\ : ClkMux
    port map (
            O => \N__49698\,
            I => \N__49176\
        );

    \I__12349\ : ClkMux
    port map (
            O => \N__49697\,
            I => \N__49176\
        );

    \I__12348\ : ClkMux
    port map (
            O => \N__49696\,
            I => \N__49176\
        );

    \I__12347\ : ClkMux
    port map (
            O => \N__49695\,
            I => \N__49176\
        );

    \I__12346\ : ClkMux
    port map (
            O => \N__49694\,
            I => \N__49176\
        );

    \I__12345\ : ClkMux
    port map (
            O => \N__49693\,
            I => \N__49176\
        );

    \I__12344\ : ClkMux
    port map (
            O => \N__49692\,
            I => \N__49176\
        );

    \I__12343\ : ClkMux
    port map (
            O => \N__49691\,
            I => \N__49176\
        );

    \I__12342\ : ClkMux
    port map (
            O => \N__49690\,
            I => \N__49176\
        );

    \I__12341\ : ClkMux
    port map (
            O => \N__49689\,
            I => \N__49176\
        );

    \I__12340\ : ClkMux
    port map (
            O => \N__49688\,
            I => \N__49176\
        );

    \I__12339\ : ClkMux
    port map (
            O => \N__49687\,
            I => \N__49176\
        );

    \I__12338\ : ClkMux
    port map (
            O => \N__49686\,
            I => \N__49176\
        );

    \I__12337\ : ClkMux
    port map (
            O => \N__49685\,
            I => \N__49176\
        );

    \I__12336\ : ClkMux
    port map (
            O => \N__49684\,
            I => \N__49176\
        );

    \I__12335\ : ClkMux
    port map (
            O => \N__49683\,
            I => \N__49176\
        );

    \I__12334\ : ClkMux
    port map (
            O => \N__49682\,
            I => \N__49176\
        );

    \I__12333\ : ClkMux
    port map (
            O => \N__49681\,
            I => \N__49176\
        );

    \I__12332\ : ClkMux
    port map (
            O => \N__49680\,
            I => \N__49176\
        );

    \I__12331\ : ClkMux
    port map (
            O => \N__49679\,
            I => \N__49176\
        );

    \I__12330\ : ClkMux
    port map (
            O => \N__49678\,
            I => \N__49176\
        );

    \I__12329\ : ClkMux
    port map (
            O => \N__49677\,
            I => \N__49176\
        );

    \I__12328\ : ClkMux
    port map (
            O => \N__49676\,
            I => \N__49176\
        );

    \I__12327\ : ClkMux
    port map (
            O => \N__49675\,
            I => \N__49176\
        );

    \I__12326\ : ClkMux
    port map (
            O => \N__49674\,
            I => \N__49176\
        );

    \I__12325\ : ClkMux
    port map (
            O => \N__49673\,
            I => \N__49176\
        );

    \I__12324\ : ClkMux
    port map (
            O => \N__49672\,
            I => \N__49176\
        );

    \I__12323\ : ClkMux
    port map (
            O => \N__49671\,
            I => \N__49176\
        );

    \I__12322\ : ClkMux
    port map (
            O => \N__49670\,
            I => \N__49176\
        );

    \I__12321\ : ClkMux
    port map (
            O => \N__49669\,
            I => \N__49176\
        );

    \I__12320\ : ClkMux
    port map (
            O => \N__49668\,
            I => \N__49176\
        );

    \I__12319\ : ClkMux
    port map (
            O => \N__49667\,
            I => \N__49176\
        );

    \I__12318\ : ClkMux
    port map (
            O => \N__49666\,
            I => \N__49176\
        );

    \I__12317\ : ClkMux
    port map (
            O => \N__49665\,
            I => \N__49176\
        );

    \I__12316\ : ClkMux
    port map (
            O => \N__49664\,
            I => \N__49176\
        );

    \I__12315\ : ClkMux
    port map (
            O => \N__49663\,
            I => \N__49176\
        );

    \I__12314\ : ClkMux
    port map (
            O => \N__49662\,
            I => \N__49176\
        );

    \I__12313\ : ClkMux
    port map (
            O => \N__49661\,
            I => \N__49176\
        );

    \I__12312\ : ClkMux
    port map (
            O => \N__49660\,
            I => \N__49176\
        );

    \I__12311\ : ClkMux
    port map (
            O => \N__49659\,
            I => \N__49176\
        );

    \I__12310\ : ClkMux
    port map (
            O => \N__49658\,
            I => \N__49176\
        );

    \I__12309\ : ClkMux
    port map (
            O => \N__49657\,
            I => \N__49176\
        );

    \I__12308\ : ClkMux
    port map (
            O => \N__49656\,
            I => \N__49176\
        );

    \I__12307\ : ClkMux
    port map (
            O => \N__49655\,
            I => \N__49176\
        );

    \I__12306\ : ClkMux
    port map (
            O => \N__49654\,
            I => \N__49176\
        );

    \I__12305\ : ClkMux
    port map (
            O => \N__49653\,
            I => \N__49176\
        );

    \I__12304\ : ClkMux
    port map (
            O => \N__49652\,
            I => \N__49176\
        );

    \I__12303\ : ClkMux
    port map (
            O => \N__49651\,
            I => \N__49176\
        );

    \I__12302\ : ClkMux
    port map (
            O => \N__49650\,
            I => \N__49176\
        );

    \I__12301\ : ClkMux
    port map (
            O => \N__49649\,
            I => \N__49176\
        );

    \I__12300\ : ClkMux
    port map (
            O => \N__49648\,
            I => \N__49176\
        );

    \I__12299\ : ClkMux
    port map (
            O => \N__49647\,
            I => \N__49176\
        );

    \I__12298\ : ClkMux
    port map (
            O => \N__49646\,
            I => \N__49176\
        );

    \I__12297\ : ClkMux
    port map (
            O => \N__49645\,
            I => \N__49176\
        );

    \I__12296\ : ClkMux
    port map (
            O => \N__49644\,
            I => \N__49176\
        );

    \I__12295\ : ClkMux
    port map (
            O => \N__49643\,
            I => \N__49176\
        );

    \I__12294\ : ClkMux
    port map (
            O => \N__49642\,
            I => \N__49176\
        );

    \I__12293\ : ClkMux
    port map (
            O => \N__49641\,
            I => \N__49176\
        );

    \I__12292\ : ClkMux
    port map (
            O => \N__49640\,
            I => \N__49176\
        );

    \I__12291\ : ClkMux
    port map (
            O => \N__49639\,
            I => \N__49176\
        );

    \I__12290\ : ClkMux
    port map (
            O => \N__49638\,
            I => \N__49176\
        );

    \I__12289\ : ClkMux
    port map (
            O => \N__49637\,
            I => \N__49176\
        );

    \I__12288\ : ClkMux
    port map (
            O => \N__49636\,
            I => \N__49176\
        );

    \I__12287\ : ClkMux
    port map (
            O => \N__49635\,
            I => \N__49176\
        );

    \I__12286\ : ClkMux
    port map (
            O => \N__49634\,
            I => \N__49176\
        );

    \I__12285\ : ClkMux
    port map (
            O => \N__49633\,
            I => \N__49176\
        );

    \I__12284\ : ClkMux
    port map (
            O => \N__49632\,
            I => \N__49176\
        );

    \I__12283\ : ClkMux
    port map (
            O => \N__49631\,
            I => \N__49176\
        );

    \I__12282\ : ClkMux
    port map (
            O => \N__49630\,
            I => \N__49176\
        );

    \I__12281\ : ClkMux
    port map (
            O => \N__49629\,
            I => \N__49176\
        );

    \I__12280\ : ClkMux
    port map (
            O => \N__49628\,
            I => \N__49176\
        );

    \I__12279\ : ClkMux
    port map (
            O => \N__49627\,
            I => \N__49176\
        );

    \I__12278\ : GlobalMux
    port map (
            O => \N__49176\,
            I => \N__49173\
        );

    \I__12277\ : gio2CtrlBuf
    port map (
            O => \N__49173\,
            I => \CLK_c\
        );

    \I__12276\ : InMux
    port map (
            O => \N__49170\,
            I => \N__49165\
        );

    \I__12275\ : InMux
    port map (
            O => \N__49169\,
            I => \N__49162\
        );

    \I__12274\ : InMux
    port map (
            O => \N__49168\,
            I => \N__49158\
        );

    \I__12273\ : LocalMux
    port map (
            O => \N__49165\,
            I => \N__49155\
        );

    \I__12272\ : LocalMux
    port map (
            O => \N__49162\,
            I => \N__49152\
        );

    \I__12271\ : CascadeMux
    port map (
            O => \N__49161\,
            I => \N__49148\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__49158\,
            I => \N__49144\
        );

    \I__12269\ : Span4Mux_v
    port map (
            O => \N__49155\,
            I => \N__49141\
        );

    \I__12268\ : Span4Mux_v
    port map (
            O => \N__49152\,
            I => \N__49138\
        );

    \I__12267\ : InMux
    port map (
            O => \N__49151\,
            I => \N__49135\
        );

    \I__12266\ : InMux
    port map (
            O => \N__49148\,
            I => \N__49132\
        );

    \I__12265\ : InMux
    port map (
            O => \N__49147\,
            I => \N__49129\
        );

    \I__12264\ : Span4Mux_v
    port map (
            O => \N__49144\,
            I => \N__49122\
        );

    \I__12263\ : Span4Mux_h
    port map (
            O => \N__49141\,
            I => \N__49122\
        );

    \I__12262\ : Span4Mux_h
    port map (
            O => \N__49138\,
            I => \N__49122\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__49135\,
            I => data_out_9_2
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__49132\,
            I => data_out_9_2
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__49129\,
            I => data_out_9_2
        );

    \I__12258\ : Odrv4
    port map (
            O => \N__49122\,
            I => data_out_9_2
        );

    \I__12257\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49106\
        );

    \I__12256\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49103\
        );

    \I__12255\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49100\
        );

    \I__12254\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49094\
        );

    \I__12253\ : InMux
    port map (
            O => \N__49109\,
            I => \N__49094\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__49106\,
            I => \N__49091\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__49103\,
            I => \N__49088\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__49100\,
            I => \N__49085\
        );

    \I__12249\ : InMux
    port map (
            O => \N__49099\,
            I => \N__49081\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__49094\,
            I => \N__49078\
        );

    \I__12247\ : Span4Mux_v
    port map (
            O => \N__49091\,
            I => \N__49075\
        );

    \I__12246\ : Span4Mux_v
    port map (
            O => \N__49088\,
            I => \N__49072\
        );

    \I__12245\ : Span4Mux_v
    port map (
            O => \N__49085\,
            I => \N__49069\
        );

    \I__12244\ : InMux
    port map (
            O => \N__49084\,
            I => \N__49066\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__49081\,
            I => \N__49060\
        );

    \I__12242\ : Span4Mux_h
    port map (
            O => \N__49078\,
            I => \N__49060\
        );

    \I__12241\ : Sp12to4
    port map (
            O => \N__49075\,
            I => \N__49051\
        );

    \I__12240\ : Sp12to4
    port map (
            O => \N__49072\,
            I => \N__49051\
        );

    \I__12239\ : Sp12to4
    port map (
            O => \N__49069\,
            I => \N__49051\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__49066\,
            I => \N__49051\
        );

    \I__12237\ : InMux
    port map (
            O => \N__49065\,
            I => \N__49048\
        );

    \I__12236\ : Odrv4
    port map (
            O => \N__49060\,
            I => \c0.data_out_5_4\
        );

    \I__12235\ : Odrv12
    port map (
            O => \N__49051\,
            I => \c0.data_out_5_4\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__49048\,
            I => \c0.data_out_5_4\
        );

    \I__12233\ : InMux
    port map (
            O => \N__49041\,
            I => \N__49037\
        );

    \I__12232\ : CascadeMux
    port map (
            O => \N__49040\,
            I => \N__49034\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__49037\,
            I => \N__49030\
        );

    \I__12230\ : InMux
    port map (
            O => \N__49034\,
            I => \N__49025\
        );

    \I__12229\ : InMux
    port map (
            O => \N__49033\,
            I => \N__49025\
        );

    \I__12228\ : Span4Mux_v
    port map (
            O => \N__49030\,
            I => \N__49022\
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__49025\,
            I => \N__49019\
        );

    \I__12226\ : Odrv4
    port map (
            O => \N__49022\,
            I => \c0.data_out_10_6\
        );

    \I__12225\ : Odrv4
    port map (
            O => \N__49019\,
            I => \c0.data_out_10_6\
        );

    \I__12224\ : InMux
    port map (
            O => \N__49014\,
            I => \N__49010\
        );

    \I__12223\ : InMux
    port map (
            O => \N__49013\,
            I => \N__49007\
        );

    \I__12222\ : LocalMux
    port map (
            O => \N__49010\,
            I => \N__49000\
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__49007\,
            I => \N__49000\
        );

    \I__12220\ : InMux
    port map (
            O => \N__49006\,
            I => \N__48997\
        );

    \I__12219\ : InMux
    port map (
            O => \N__49005\,
            I => \N__48994\
        );

    \I__12218\ : Span4Mux_v
    port map (
            O => \N__49000\,
            I => \N__48991\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__48997\,
            I => \N__48988\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__48994\,
            I => \c0.data_out_9_3\
        );

    \I__12215\ : Odrv4
    port map (
            O => \N__48991\,
            I => \c0.data_out_9_3\
        );

    \I__12214\ : Odrv4
    port map (
            O => \N__48988\,
            I => \c0.data_out_9_3\
        );

    \I__12213\ : CascadeMux
    port map (
            O => \N__48981\,
            I => \c0.n10204_cascade_\
        );

    \I__12212\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48975\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__48975\,
            I => \N__48972\
        );

    \I__12210\ : Span4Mux_v
    port map (
            O => \N__48972\,
            I => \N__48968\
        );

    \I__12209\ : InMux
    port map (
            O => \N__48971\,
            I => \N__48965\
        );

    \I__12208\ : Sp12to4
    port map (
            O => \N__48968\,
            I => \N__48958\
        );

    \I__12207\ : LocalMux
    port map (
            O => \N__48965\,
            I => \N__48958\
        );

    \I__12206\ : InMux
    port map (
            O => \N__48964\,
            I => \N__48953\
        );

    \I__12205\ : InMux
    port map (
            O => \N__48963\,
            I => \N__48953\
        );

    \I__12204\ : Odrv12
    port map (
            O => \N__48958\,
            I => \c0.data_out_7_4\
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__48953\,
            I => \c0.data_out_7_4\
        );

    \I__12202\ : CascadeMux
    port map (
            O => \N__48948\,
            I => \N__48945\
        );

    \I__12201\ : InMux
    port map (
            O => \N__48945\,
            I => \N__48942\
        );

    \I__12200\ : LocalMux
    port map (
            O => \N__48942\,
            I => \N__48939\
        );

    \I__12199\ : Span4Mux_v
    port map (
            O => \N__48939\,
            I => \N__48936\
        );

    \I__12198\ : Odrv4
    port map (
            O => \N__48936\,
            I => \c0.n10_adj_2172\
        );

    \I__12197\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48930\
        );

    \I__12196\ : LocalMux
    port map (
            O => \N__48930\,
            I => \N__48927\
        );

    \I__12195\ : Span4Mux_h
    port map (
            O => \N__48927\,
            I => \N__48922\
        );

    \I__12194\ : InMux
    port map (
            O => \N__48926\,
            I => \N__48919\
        );

    \I__12193\ : InMux
    port map (
            O => \N__48925\,
            I => \N__48916\
        );

    \I__12192\ : Span4Mux_h
    port map (
            O => \N__48922\,
            I => \N__48913\
        );

    \I__12191\ : LocalMux
    port map (
            O => \N__48919\,
            I => \N__48908\
        );

    \I__12190\ : LocalMux
    port map (
            O => \N__48916\,
            I => \N__48908\
        );

    \I__12189\ : Odrv4
    port map (
            O => \N__48913\,
            I => \c0.data_out_6_7\
        );

    \I__12188\ : Odrv12
    port map (
            O => \N__48908\,
            I => \c0.data_out_6_7\
        );

    \I__12187\ : InMux
    port map (
            O => \N__48903\,
            I => \N__48900\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__48900\,
            I => \N__48897\
        );

    \I__12185\ : Span4Mux_h
    port map (
            O => \N__48897\,
            I => \N__48893\
        );

    \I__12184\ : InMux
    port map (
            O => \N__48896\,
            I => \N__48890\
        );

    \I__12183\ : Odrv4
    port map (
            O => \N__48893\,
            I => \c0.n26_adj_2165\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__48890\,
            I => \c0.n26_adj_2165\
        );

    \I__12181\ : InMux
    port map (
            O => \N__48885\,
            I => \N__48880\
        );

    \I__12180\ : InMux
    port map (
            O => \N__48884\,
            I => \N__48877\
        );

    \I__12179\ : InMux
    port map (
            O => \N__48883\,
            I => \N__48874\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__48880\,
            I => \N__48871\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48868\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__48874\,
            I => \N__48865\
        );

    \I__12175\ : Span4Mux_v
    port map (
            O => \N__48871\,
            I => \N__48861\
        );

    \I__12174\ : Span4Mux_h
    port map (
            O => \N__48868\,
            I => \N__48858\
        );

    \I__12173\ : Span4Mux_h
    port map (
            O => \N__48865\,
            I => \N__48855\
        );

    \I__12172\ : InMux
    port map (
            O => \N__48864\,
            I => \N__48852\
        );

    \I__12171\ : Span4Mux_h
    port map (
            O => \N__48861\,
            I => \N__48849\
        );

    \I__12170\ : Span4Mux_h
    port map (
            O => \N__48858\,
            I => \N__48844\
        );

    \I__12169\ : Span4Mux_v
    port map (
            O => \N__48855\,
            I => \N__48844\
        );

    \I__12168\ : LocalMux
    port map (
            O => \N__48852\,
            I => \N__48841\
        );

    \I__12167\ : Odrv4
    port map (
            O => \N__48849\,
            I => \c0.data_out_6_5\
        );

    \I__12166\ : Odrv4
    port map (
            O => \N__48844\,
            I => \c0.data_out_6_5\
        );

    \I__12165\ : Odrv4
    port map (
            O => \N__48841\,
            I => \c0.data_out_6_5\
        );

    \I__12164\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48831\
        );

    \I__12163\ : LocalMux
    port map (
            O => \N__48831\,
            I => \N__48828\
        );

    \I__12162\ : Span4Mux_v
    port map (
            O => \N__48828\,
            I => \N__48822\
        );

    \I__12161\ : InMux
    port map (
            O => \N__48827\,
            I => \N__48819\
        );

    \I__12160\ : InMux
    port map (
            O => \N__48826\,
            I => \N__48816\
        );

    \I__12159\ : InMux
    port map (
            O => \N__48825\,
            I => \N__48812\
        );

    \I__12158\ : Sp12to4
    port map (
            O => \N__48822\,
            I => \N__48805\
        );

    \I__12157\ : LocalMux
    port map (
            O => \N__48819\,
            I => \N__48805\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__48816\,
            I => \N__48805\
        );

    \I__12155\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48802\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__48812\,
            I => data_out_8_3
        );

    \I__12153\ : Odrv12
    port map (
            O => \N__48805\,
            I => data_out_8_3
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__48802\,
            I => data_out_8_3
        );

    \I__12151\ : CascadeMux
    port map (
            O => \N__48795\,
            I => \c0.n10_adj_2166_cascade_\
        );

    \I__12150\ : CascadeMux
    port map (
            O => \N__48792\,
            I => \N__48788\
        );

    \I__12149\ : InMux
    port map (
            O => \N__48791\,
            I => \N__48785\
        );

    \I__12148\ : InMux
    port map (
            O => \N__48788\,
            I => \N__48782\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__48785\,
            I => \N__48779\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__48782\,
            I => \c0.n10170\
        );

    \I__12145\ : Odrv4
    port map (
            O => \N__48779\,
            I => \c0.n10170\
        );

    \I__12144\ : InMux
    port map (
            O => \N__48774\,
            I => \N__48771\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__48771\,
            I => \N__48767\
        );

    \I__12142\ : InMux
    port map (
            O => \N__48770\,
            I => \N__48764\
        );

    \I__12141\ : Odrv12
    port map (
            O => \N__48767\,
            I => \c0.n17252\
        );

    \I__12140\ : LocalMux
    port map (
            O => \N__48764\,
            I => \c0.n17252\
        );

    \I__12139\ : CascadeMux
    port map (
            O => \N__48759\,
            I => \N__48756\
        );

    \I__12138\ : InMux
    port map (
            O => \N__48756\,
            I => \N__48753\
        );

    \I__12137\ : LocalMux
    port map (
            O => \N__48753\,
            I => \N__48750\
        );

    \I__12136\ : Span4Mux_v
    port map (
            O => \N__48750\,
            I => \N__48747\
        );

    \I__12135\ : Span4Mux_h
    port map (
            O => \N__48747\,
            I => \N__48742\
        );

    \I__12134\ : InMux
    port map (
            O => \N__48746\,
            I => \N__48737\
        );

    \I__12133\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48737\
        );

    \I__12132\ : Odrv4
    port map (
            O => \N__48742\,
            I => data_out_10_1
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__48737\,
            I => data_out_10_1
        );

    \I__12130\ : InMux
    port map (
            O => \N__48732\,
            I => \N__48729\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__48729\,
            I => \N__48725\
        );

    \I__12128\ : InMux
    port map (
            O => \N__48728\,
            I => \N__48722\
        );

    \I__12127\ : Span4Mux_h
    port map (
            O => \N__48725\,
            I => \N__48719\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__48722\,
            I => \N__48714\
        );

    \I__12125\ : Span4Mux_h
    port map (
            O => \N__48719\,
            I => \N__48710\
        );

    \I__12124\ : InMux
    port map (
            O => \N__48718\,
            I => \N__48707\
        );

    \I__12123\ : InMux
    port map (
            O => \N__48717\,
            I => \N__48704\
        );

    \I__12122\ : Span4Mux_h
    port map (
            O => \N__48714\,
            I => \N__48701\
        );

    \I__12121\ : InMux
    port map (
            O => \N__48713\,
            I => \N__48698\
        );

    \I__12120\ : Odrv4
    port map (
            O => \N__48710\,
            I => data_out_8_2
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__48707\,
            I => data_out_8_2
        );

    \I__12118\ : LocalMux
    port map (
            O => \N__48704\,
            I => data_out_8_2
        );

    \I__12117\ : Odrv4
    port map (
            O => \N__48701\,
            I => data_out_8_2
        );

    \I__12116\ : LocalMux
    port map (
            O => \N__48698\,
            I => data_out_8_2
        );

    \I__12115\ : CascadeMux
    port map (
            O => \N__48687\,
            I => \N__48684\
        );

    \I__12114\ : InMux
    port map (
            O => \N__48684\,
            I => \N__48680\
        );

    \I__12113\ : InMux
    port map (
            O => \N__48683\,
            I => \N__48677\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__48680\,
            I => \N__48674\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__48677\,
            I => \N__48668\
        );

    \I__12110\ : Span4Mux_s3_v
    port map (
            O => \N__48674\,
            I => \N__48668\
        );

    \I__12109\ : InMux
    port map (
            O => \N__48673\,
            I => \N__48665\
        );

    \I__12108\ : Odrv4
    port map (
            O => \N__48668\,
            I => \c0.data_out_10_5\
        );

    \I__12107\ : LocalMux
    port map (
            O => \N__48665\,
            I => \c0.data_out_10_5\
        );

    \I__12106\ : InMux
    port map (
            O => \N__48660\,
            I => \N__48656\
        );

    \I__12105\ : InMux
    port map (
            O => \N__48659\,
            I => \N__48653\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__48656\,
            I => \N__48647\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__48653\,
            I => \N__48647\
        );

    \I__12102\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48644\
        );

    \I__12101\ : Span4Mux_v
    port map (
            O => \N__48647\,
            I => \N__48641\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__48644\,
            I => \N__48638\
        );

    \I__12099\ : Span4Mux_h
    port map (
            O => \N__48641\,
            I => \N__48635\
        );

    \I__12098\ : Span4Mux_h
    port map (
            O => \N__48638\,
            I => \N__48632\
        );

    \I__12097\ : Span4Mux_h
    port map (
            O => \N__48635\,
            I => \N__48629\
        );

    \I__12096\ : Span4Mux_h
    port map (
            O => \N__48632\,
            I => \N__48626\
        );

    \I__12095\ : Odrv4
    port map (
            O => \N__48629\,
            I => \c0.data_out_7_1\
        );

    \I__12094\ : Odrv4
    port map (
            O => \N__48626\,
            I => \c0.data_out_7_1\
        );

    \I__12093\ : InMux
    port map (
            O => \N__48621\,
            I => \N__48617\
        );

    \I__12092\ : CascadeMux
    port map (
            O => \N__48620\,
            I => \N__48611\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__48617\,
            I => \N__48608\
        );

    \I__12090\ : InMux
    port map (
            O => \N__48616\,
            I => \N__48603\
        );

    \I__12089\ : InMux
    port map (
            O => \N__48615\,
            I => \N__48603\
        );

    \I__12088\ : InMux
    port map (
            O => \N__48614\,
            I => \N__48598\
        );

    \I__12087\ : InMux
    port map (
            O => \N__48611\,
            I => \N__48598\
        );

    \I__12086\ : Odrv4
    port map (
            O => \N__48608\,
            I => \c0.data_out_9_0\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__48603\,
            I => \c0.data_out_9_0\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__48598\,
            I => \c0.data_out_9_0\
        );

    \I__12083\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48588\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__48588\,
            I => \N__48585\
        );

    \I__12081\ : Odrv4
    port map (
            O => \N__48585\,
            I => \c0.n6_adj_2169\
        );

    \I__12080\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48579\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__48579\,
            I => \c0.n17162\
        );

    \I__12078\ : CascadeMux
    port map (
            O => \N__48576\,
            I => \c0.n17150_cascade_\
        );

    \I__12077\ : InMux
    port map (
            O => \N__48573\,
            I => \N__48567\
        );

    \I__12076\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48561\
        );

    \I__12075\ : InMux
    port map (
            O => \N__48571\,
            I => \N__48561\
        );

    \I__12074\ : InMux
    port map (
            O => \N__48570\,
            I => \N__48558\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__48567\,
            I => \N__48555\
        );

    \I__12072\ : InMux
    port map (
            O => \N__48566\,
            I => \N__48552\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__48561\,
            I => \N__48549\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__48558\,
            I => \N__48546\
        );

    \I__12069\ : Span4Mux_h
    port map (
            O => \N__48555\,
            I => \N__48543\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__48552\,
            I => \c0.data_out_9_1\
        );

    \I__12067\ : Odrv4
    port map (
            O => \N__48549\,
            I => \c0.data_out_9_1\
        );

    \I__12066\ : Odrv4
    port map (
            O => \N__48546\,
            I => \c0.data_out_9_1\
        );

    \I__12065\ : Odrv4
    port map (
            O => \N__48543\,
            I => \c0.data_out_9_1\
        );

    \I__12064\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48529\
        );

    \I__12063\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48526\
        );

    \I__12062\ : InMux
    port map (
            O => \N__48532\,
            I => \N__48523\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__48529\,
            I => \N__48518\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__48526\,
            I => \N__48518\
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__48523\,
            I => \N__48513\
        );

    \I__12058\ : Span4Mux_h
    port map (
            O => \N__48518\,
            I => \N__48513\
        );

    \I__12057\ : Odrv4
    port map (
            O => \N__48513\,
            I => \c0.data_out_9_5\
        );

    \I__12056\ : InMux
    port map (
            O => \N__48510\,
            I => \N__48507\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__48507\,
            I => \N__48504\
        );

    \I__12054\ : Span4Mux_h
    port map (
            O => \N__48504\,
            I => \N__48501\
        );

    \I__12053\ : Span4Mux_v
    port map (
            O => \N__48501\,
            I => \N__48497\
        );

    \I__12052\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48494\
        );

    \I__12051\ : Sp12to4
    port map (
            O => \N__48497\,
            I => \N__48489\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__48494\,
            I => \N__48489\
        );

    \I__12049\ : Span12Mux_h
    port map (
            O => \N__48489\,
            I => \N__48486\
        );

    \I__12048\ : Odrv12
    port map (
            O => \N__48486\,
            I => \c0.n17110\
        );

    \I__12047\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48477\
        );

    \I__12046\ : InMux
    port map (
            O => \N__48482\,
            I => \N__48477\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__48477\,
            I => \N__48474\
        );

    \I__12044\ : Sp12to4
    port map (
            O => \N__48474\,
            I => \N__48469\
        );

    \I__12043\ : InMux
    port map (
            O => \N__48473\,
            I => \N__48466\
        );

    \I__12042\ : InMux
    port map (
            O => \N__48472\,
            I => \N__48462\
        );

    \I__12041\ : Span12Mux_s5_v
    port map (
            O => \N__48469\,
            I => \N__48457\
        );

    \I__12040\ : LocalMux
    port map (
            O => \N__48466\,
            I => \N__48457\
        );

    \I__12039\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48454\
        );

    \I__12038\ : LocalMux
    port map (
            O => \N__48462\,
            I => data_out_8_4
        );

    \I__12037\ : Odrv12
    port map (
            O => \N__48457\,
            I => data_out_8_4
        );

    \I__12036\ : LocalMux
    port map (
            O => \N__48454\,
            I => data_out_8_4
        );

    \I__12035\ : InMux
    port map (
            O => \N__48447\,
            I => \N__48443\
        );

    \I__12034\ : InMux
    port map (
            O => \N__48446\,
            I => \N__48440\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__48443\,
            I => \N__48437\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__48440\,
            I => \N__48434\
        );

    \I__12031\ : Span4Mux_h
    port map (
            O => \N__48437\,
            I => \N__48431\
        );

    \I__12030\ : Odrv4
    port map (
            O => \N__48434\,
            I => \c0.data_out_10_7\
        );

    \I__12029\ : Odrv4
    port map (
            O => \N__48431\,
            I => \c0.data_out_10_7\
        );

    \I__12028\ : InMux
    port map (
            O => \N__48426\,
            I => \N__48422\
        );

    \I__12027\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48413\
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48406\
        );

    \I__12025\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48401\
        );

    \I__12024\ : InMux
    port map (
            O => \N__48420\,
            I => \N__48396\
        );

    \I__12023\ : InMux
    port map (
            O => \N__48419\,
            I => \N__48396\
        );

    \I__12022\ : CascadeMux
    port map (
            O => \N__48418\,
            I => \N__48393\
        );

    \I__12021\ : CascadeMux
    port map (
            O => \N__48417\,
            I => \N__48389\
        );

    \I__12020\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48385\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__48413\,
            I => \N__48376\
        );

    \I__12018\ : InMux
    port map (
            O => \N__48412\,
            I => \N__48373\
        );

    \I__12017\ : CascadeMux
    port map (
            O => \N__48411\,
            I => \N__48368\
        );

    \I__12016\ : CascadeMux
    port map (
            O => \N__48410\,
            I => \N__48365\
        );

    \I__12015\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48362\
        );

    \I__12014\ : Span4Mux_h
    port map (
            O => \N__48406\,
            I => \N__48359\
        );

    \I__12013\ : InMux
    port map (
            O => \N__48405\,
            I => \N__48356\
        );

    \I__12012\ : CascadeMux
    port map (
            O => \N__48404\,
            I => \N__48353\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__48401\,
            I => \N__48348\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__48396\,
            I => \N__48348\
        );

    \I__12009\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48343\
        );

    \I__12008\ : InMux
    port map (
            O => \N__48392\,
            I => \N__48343\
        );

    \I__12007\ : InMux
    port map (
            O => \N__48389\,
            I => \N__48340\
        );

    \I__12006\ : InMux
    port map (
            O => \N__48388\,
            I => \N__48337\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__48385\,
            I => \N__48334\
        );

    \I__12004\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48331\
        );

    \I__12003\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48328\
        );

    \I__12002\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48325\
        );

    \I__12001\ : InMux
    port map (
            O => \N__48381\,
            I => \N__48322\
        );

    \I__12000\ : InMux
    port map (
            O => \N__48380\,
            I => \N__48319\
        );

    \I__11999\ : CascadeMux
    port map (
            O => \N__48379\,
            I => \N__48316\
        );

    \I__11998\ : Span4Mux_v
    port map (
            O => \N__48376\,
            I => \N__48310\
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48307\
        );

    \I__11996\ : InMux
    port map (
            O => \N__48372\,
            I => \N__48304\
        );

    \I__11995\ : CascadeMux
    port map (
            O => \N__48371\,
            I => \N__48299\
        );

    \I__11994\ : InMux
    port map (
            O => \N__48368\,
            I => \N__48295\
        );

    \I__11993\ : InMux
    port map (
            O => \N__48365\,
            I => \N__48292\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__48362\,
            I => \N__48285\
        );

    \I__11991\ : Span4Mux_h
    port map (
            O => \N__48359\,
            I => \N__48285\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__48356\,
            I => \N__48285\
        );

    \I__11989\ : InMux
    port map (
            O => \N__48353\,
            I => \N__48282\
        );

    \I__11988\ : Span4Mux_h
    port map (
            O => \N__48348\,
            I => \N__48279\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__48343\,
            I => \N__48273\
        );

    \I__11986\ : LocalMux
    port map (
            O => \N__48340\,
            I => \N__48264\
        );

    \I__11985\ : LocalMux
    port map (
            O => \N__48337\,
            I => \N__48264\
        );

    \I__11984\ : Span4Mux_h
    port map (
            O => \N__48334\,
            I => \N__48264\
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__48331\,
            I => \N__48264\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__48328\,
            I => \N__48259\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__48325\,
            I => \N__48259\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__48322\,
            I => \N__48254\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__48319\,
            I => \N__48254\
        );

    \I__11978\ : InMux
    port map (
            O => \N__48316\,
            I => \N__48247\
        );

    \I__11977\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48247\
        );

    \I__11976\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48247\
        );

    \I__11975\ : InMux
    port map (
            O => \N__48313\,
            I => \N__48244\
        );

    \I__11974\ : Span4Mux_h
    port map (
            O => \N__48310\,
            I => \N__48241\
        );

    \I__11973\ : Span4Mux_v
    port map (
            O => \N__48307\,
            I => \N__48236\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__48304\,
            I => \N__48236\
        );

    \I__11971\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48233\
        );

    \I__11970\ : InMux
    port map (
            O => \N__48302\,
            I => \N__48230\
        );

    \I__11969\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48225\
        );

    \I__11968\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48225\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__48295\,
            I => \N__48220\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__48292\,
            I => \N__48220\
        );

    \I__11965\ : Span4Mux_v
    port map (
            O => \N__48285\,
            I => \N__48217\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__48282\,
            I => \N__48212\
        );

    \I__11963\ : Span4Mux_h
    port map (
            O => \N__48279\,
            I => \N__48212\
        );

    \I__11962\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48205\
        );

    \I__11961\ : InMux
    port map (
            O => \N__48277\,
            I => \N__48205\
        );

    \I__11960\ : InMux
    port map (
            O => \N__48276\,
            I => \N__48205\
        );

    \I__11959\ : Span4Mux_h
    port map (
            O => \N__48273\,
            I => \N__48198\
        );

    \I__11958\ : Span4Mux_v
    port map (
            O => \N__48264\,
            I => \N__48198\
        );

    \I__11957\ : Span4Mux_v
    port map (
            O => \N__48259\,
            I => \N__48198\
        );

    \I__11956\ : Span4Mux_h
    port map (
            O => \N__48254\,
            I => \N__48187\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__48247\,
            I => \N__48187\
        );

    \I__11954\ : LocalMux
    port map (
            O => \N__48244\,
            I => \N__48187\
        );

    \I__11953\ : Span4Mux_v
    port map (
            O => \N__48241\,
            I => \N__48187\
        );

    \I__11952\ : Span4Mux_h
    port map (
            O => \N__48236\,
            I => \N__48187\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__48233\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11950\ : LocalMux
    port map (
            O => \N__48230\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__48225\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11948\ : Odrv12
    port map (
            O => \N__48220\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11947\ : Odrv4
    port map (
            O => \N__48217\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11946\ : Odrv4
    port map (
            O => \N__48212\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__48205\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11944\ : Odrv4
    port map (
            O => \N__48198\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11943\ : Odrv4
    port map (
            O => \N__48187\,
            I => \UART_TRANSMITTER_state_2\
        );

    \I__11942\ : InMux
    port map (
            O => \N__48168\,
            I => \N__48161\
        );

    \I__11941\ : InMux
    port map (
            O => \N__48167\,
            I => \N__48158\
        );

    \I__11940\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48145\
        );

    \I__11939\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48145\
        );

    \I__11938\ : InMux
    port map (
            O => \N__48164\,
            I => \N__48141\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__48161\,
            I => \N__48138\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__48158\,
            I => \N__48135\
        );

    \I__11935\ : CascadeMux
    port map (
            O => \N__48157\,
            I => \N__48124\
        );

    \I__11934\ : InMux
    port map (
            O => \N__48156\,
            I => \N__48118\
        );

    \I__11933\ : CascadeMux
    port map (
            O => \N__48155\,
            I => \N__48115\
        );

    \I__11932\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48101\
        );

    \I__11931\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48101\
        );

    \I__11930\ : InMux
    port map (
            O => \N__48152\,
            I => \N__48101\
        );

    \I__11929\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48101\
        );

    \I__11928\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48096\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__48145\,
            I => \N__48093\
        );

    \I__11926\ : CascadeMux
    port map (
            O => \N__48144\,
            I => \N__48090\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__48141\,
            I => \N__48085\
        );

    \I__11924\ : Span4Mux_v
    port map (
            O => \N__48138\,
            I => \N__48082\
        );

    \I__11923\ : Span4Mux_v
    port map (
            O => \N__48135\,
            I => \N__48079\
        );

    \I__11922\ : InMux
    port map (
            O => \N__48134\,
            I => \N__48076\
        );

    \I__11921\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48073\
        );

    \I__11920\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48066\
        );

    \I__11919\ : InMux
    port map (
            O => \N__48131\,
            I => \N__48066\
        );

    \I__11918\ : InMux
    port map (
            O => \N__48130\,
            I => \N__48066\
        );

    \I__11917\ : InMux
    port map (
            O => \N__48129\,
            I => \N__48059\
        );

    \I__11916\ : InMux
    port map (
            O => \N__48128\,
            I => \N__48059\
        );

    \I__11915\ : InMux
    port map (
            O => \N__48127\,
            I => \N__48059\
        );

    \I__11914\ : InMux
    port map (
            O => \N__48124\,
            I => \N__48050\
        );

    \I__11913\ : InMux
    port map (
            O => \N__48123\,
            I => \N__48050\
        );

    \I__11912\ : InMux
    port map (
            O => \N__48122\,
            I => \N__48050\
        );

    \I__11911\ : InMux
    port map (
            O => \N__48121\,
            I => \N__48050\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__48047\
        );

    \I__11909\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48042\
        );

    \I__11908\ : InMux
    port map (
            O => \N__48114\,
            I => \N__48042\
        );

    \I__11907\ : InMux
    port map (
            O => \N__48113\,
            I => \N__48039\
        );

    \I__11906\ : InMux
    port map (
            O => \N__48112\,
            I => \N__48036\
        );

    \I__11905\ : InMux
    port map (
            O => \N__48111\,
            I => \N__48033\
        );

    \I__11904\ : InMux
    port map (
            O => \N__48110\,
            I => \N__48029\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__48026\
        );

    \I__11902\ : CascadeMux
    port map (
            O => \N__48100\,
            I => \N__48023\
        );

    \I__11901\ : CascadeMux
    port map (
            O => \N__48099\,
            I => \N__48017\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__48096\,
            I => \N__48014\
        );

    \I__11899\ : Span12Mux_s8_v
    port map (
            O => \N__48093\,
            I => \N__48011\
        );

    \I__11898\ : InMux
    port map (
            O => \N__48090\,
            I => \N__48008\
        );

    \I__11897\ : InMux
    port map (
            O => \N__48089\,
            I => \N__48003\
        );

    \I__11896\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48003\
        );

    \I__11895\ : Span4Mux_h
    port map (
            O => \N__48085\,
            I => \N__47996\
        );

    \I__11894\ : Span4Mux_h
    port map (
            O => \N__48082\,
            I => \N__47996\
        );

    \I__11893\ : Span4Mux_h
    port map (
            O => \N__48079\,
            I => \N__47996\
        );

    \I__11892\ : LocalMux
    port map (
            O => \N__48076\,
            I => \N__47993\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__48073\,
            I => \N__47990\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__48066\,
            I => \N__47987\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__48059\,
            I => \N__47978\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__48050\,
            I => \N__47978\
        );

    \I__11887\ : Span4Mux_h
    port map (
            O => \N__48047\,
            I => \N__47978\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__48042\,
            I => \N__47978\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__48039\,
            I => \N__47971\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__48036\,
            I => \N__47971\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__48033\,
            I => \N__47971\
        );

    \I__11882\ : InMux
    port map (
            O => \N__48032\,
            I => \N__47968\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__48029\,
            I => \N__47965\
        );

    \I__11880\ : Span4Mux_h
    port map (
            O => \N__48026\,
            I => \N__47962\
        );

    \I__11879\ : InMux
    port map (
            O => \N__48023\,
            I => \N__47959\
        );

    \I__11878\ : InMux
    port map (
            O => \N__48022\,
            I => \N__47956\
        );

    \I__11877\ : InMux
    port map (
            O => \N__48021\,
            I => \N__47953\
        );

    \I__11876\ : InMux
    port map (
            O => \N__48020\,
            I => \N__47948\
        );

    \I__11875\ : InMux
    port map (
            O => \N__48017\,
            I => \N__47948\
        );

    \I__11874\ : Sp12to4
    port map (
            O => \N__48014\,
            I => \N__47941\
        );

    \I__11873\ : Span12Mux_h
    port map (
            O => \N__48011\,
            I => \N__47941\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__48008\,
            I => \N__47941\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__48003\,
            I => \N__47938\
        );

    \I__11870\ : Span4Mux_v
    port map (
            O => \N__47996\,
            I => \N__47935\
        );

    \I__11869\ : Span4Mux_h
    port map (
            O => \N__47993\,
            I => \N__47924\
        );

    \I__11868\ : Span4Mux_s2_v
    port map (
            O => \N__47990\,
            I => \N__47924\
        );

    \I__11867\ : Span4Mux_h
    port map (
            O => \N__47987\,
            I => \N__47924\
        );

    \I__11866\ : Span4Mux_v
    port map (
            O => \N__47978\,
            I => \N__47924\
        );

    \I__11865\ : Span4Mux_s2_v
    port map (
            O => \N__47971\,
            I => \N__47924\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__47968\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11863\ : Odrv4
    port map (
            O => \N__47965\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11862\ : Odrv4
    port map (
            O => \N__47962\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__47959\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__47956\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__47953\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__47948\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11857\ : Odrv12
    port map (
            O => \N__47941\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11856\ : Odrv12
    port map (
            O => \N__47938\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11855\ : Odrv4
    port map (
            O => \N__47935\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11854\ : Odrv4
    port map (
            O => \N__47924\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__11853\ : CascadeMux
    port map (
            O => \N__47901\,
            I => \N__47898\
        );

    \I__11852\ : InMux
    port map (
            O => \N__47898\,
            I => \N__47895\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__47895\,
            I => \N__47891\
        );

    \I__11850\ : CascadeMux
    port map (
            O => \N__47894\,
            I => \N__47888\
        );

    \I__11849\ : Span12Mux_s4_v
    port map (
            O => \N__47891\,
            I => \N__47885\
        );

    \I__11848\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47882\
        );

    \I__11847\ : Odrv12
    port map (
            O => \N__47885\,
            I => rand_setpoint_25
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__47882\,
            I => rand_setpoint_25
        );

    \I__11845\ : InMux
    port map (
            O => \N__47877\,
            I => \N__47866\
        );

    \I__11844\ : InMux
    port map (
            O => \N__47876\,
            I => \N__47866\
        );

    \I__11843\ : InMux
    port map (
            O => \N__47875\,
            I => \N__47866\
        );

    \I__11842\ : InMux
    port map (
            O => \N__47874\,
            I => \N__47861\
        );

    \I__11841\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47861\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__47866\,
            I => \N__47858\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__47861\,
            I => \N__47853\
        );

    \I__11838\ : Span4Mux_h
    port map (
            O => \N__47858\,
            I => \N__47853\
        );

    \I__11837\ : Span4Mux_h
    port map (
            O => \N__47853\,
            I => \N__47850\
        );

    \I__11836\ : Odrv4
    port map (
            O => \N__47850\,
            I => data_out_5_1
        );

    \I__11835\ : CascadeMux
    port map (
            O => \N__47847\,
            I => \N__47843\
        );

    \I__11834\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47835\
        );

    \I__11833\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47822\
        );

    \I__11832\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47814\
        );

    \I__11831\ : InMux
    port map (
            O => \N__47841\,
            I => \N__47806\
        );

    \I__11830\ : InMux
    port map (
            O => \N__47840\,
            I => \N__47806\
        );

    \I__11829\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47797\
        );

    \I__11828\ : InMux
    port map (
            O => \N__47838\,
            I => \N__47797\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__47835\,
            I => \N__47788\
        );

    \I__11826\ : InMux
    port map (
            O => \N__47834\,
            I => \N__47782\
        );

    \I__11825\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47782\
        );

    \I__11824\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47777\
        );

    \I__11823\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47777\
        );

    \I__11822\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47772\
        );

    \I__11821\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47772\
        );

    \I__11820\ : InMux
    port map (
            O => \N__47828\,
            I => \N__47769\
        );

    \I__11819\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47764\
        );

    \I__11818\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47764\
        );

    \I__11817\ : CascadeMux
    port map (
            O => \N__47825\,
            I => \N__47761\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__47822\,
            I => \N__47758\
        );

    \I__11815\ : InMux
    port map (
            O => \N__47821\,
            I => \N__47755\
        );

    \I__11814\ : InMux
    port map (
            O => \N__47820\,
            I => \N__47752\
        );

    \I__11813\ : InMux
    port map (
            O => \N__47819\,
            I => \N__47749\
        );

    \I__11812\ : InMux
    port map (
            O => \N__47818\,
            I => \N__47744\
        );

    \I__11811\ : InMux
    port map (
            O => \N__47817\,
            I => \N__47744\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__47814\,
            I => \N__47741\
        );

    \I__11809\ : InMux
    port map (
            O => \N__47813\,
            I => \N__47733\
        );

    \I__11808\ : InMux
    port map (
            O => \N__47812\,
            I => \N__47733\
        );

    \I__11807\ : InMux
    port map (
            O => \N__47811\,
            I => \N__47733\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__47806\,
            I => \N__47730\
        );

    \I__11805\ : InMux
    port map (
            O => \N__47805\,
            I => \N__47723\
        );

    \I__11804\ : InMux
    port map (
            O => \N__47804\,
            I => \N__47723\
        );

    \I__11803\ : InMux
    port map (
            O => \N__47803\,
            I => \N__47723\
        );

    \I__11802\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47720\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__47797\,
            I => \N__47717\
        );

    \I__11800\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47714\
        );

    \I__11799\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47709\
        );

    \I__11798\ : InMux
    port map (
            O => \N__47794\,
            I => \N__47709\
        );

    \I__11797\ : InMux
    port map (
            O => \N__47793\,
            I => \N__47704\
        );

    \I__11796\ : InMux
    port map (
            O => \N__47792\,
            I => \N__47704\
        );

    \I__11795\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47701\
        );

    \I__11794\ : Span4Mux_h
    port map (
            O => \N__47788\,
            I => \N__47697\
        );

    \I__11793\ : InMux
    port map (
            O => \N__47787\,
            I => \N__47694\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__47782\,
            I => \N__47689\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__47777\,
            I => \N__47689\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__47772\,
            I => \N__47686\
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__47769\,
            I => \N__47681\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__47764\,
            I => \N__47681\
        );

    \I__11787\ : InMux
    port map (
            O => \N__47761\,
            I => \N__47678\
        );

    \I__11786\ : Span4Mux_h
    port map (
            O => \N__47758\,
            I => \N__47662\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__47755\,
            I => \N__47662\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__47752\,
            I => \N__47662\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__47749\,
            I => \N__47657\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__47744\,
            I => \N__47657\
        );

    \I__11781\ : Span4Mux_v
    port map (
            O => \N__47741\,
            I => \N__47654\
        );

    \I__11780\ : InMux
    port map (
            O => \N__47740\,
            I => \N__47650\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__47733\,
            I => \N__47637\
        );

    \I__11778\ : Span4Mux_h
    port map (
            O => \N__47730\,
            I => \N__47637\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__47723\,
            I => \N__47637\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__47720\,
            I => \N__47637\
        );

    \I__11775\ : Span4Mux_v
    port map (
            O => \N__47717\,
            I => \N__47637\
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__47714\,
            I => \N__47637\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__47709\,
            I => \N__47630\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__47704\,
            I => \N__47630\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__47701\,
            I => \N__47630\
        );

    \I__11770\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47627\
        );

    \I__11769\ : Span4Mux_v
    port map (
            O => \N__47697\,
            I => \N__47622\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__47694\,
            I => \N__47622\
        );

    \I__11767\ : Span4Mux_v
    port map (
            O => \N__47689\,
            I => \N__47613\
        );

    \I__11766\ : Span4Mux_h
    port map (
            O => \N__47686\,
            I => \N__47613\
        );

    \I__11765\ : Span4Mux_s2_v
    port map (
            O => \N__47681\,
            I => \N__47613\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__47678\,
            I => \N__47613\
        );

    \I__11763\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47608\
        );

    \I__11762\ : InMux
    port map (
            O => \N__47676\,
            I => \N__47608\
        );

    \I__11761\ : InMux
    port map (
            O => \N__47675\,
            I => \N__47599\
        );

    \I__11760\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47599\
        );

    \I__11759\ : InMux
    port map (
            O => \N__47673\,
            I => \N__47599\
        );

    \I__11758\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47599\
        );

    \I__11757\ : InMux
    port map (
            O => \N__47671\,
            I => \N__47596\
        );

    \I__11756\ : InMux
    port map (
            O => \N__47670\,
            I => \N__47591\
        );

    \I__11755\ : InMux
    port map (
            O => \N__47669\,
            I => \N__47591\
        );

    \I__11754\ : Span4Mux_v
    port map (
            O => \N__47662\,
            I => \N__47586\
        );

    \I__11753\ : Span4Mux_s3_v
    port map (
            O => \N__47657\,
            I => \N__47586\
        );

    \I__11752\ : Span4Mux_h
    port map (
            O => \N__47654\,
            I => \N__47583\
        );

    \I__11751\ : InMux
    port map (
            O => \N__47653\,
            I => \N__47580\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__47650\,
            I => \N__47575\
        );

    \I__11749\ : Span4Mux_h
    port map (
            O => \N__47637\,
            I => \N__47575\
        );

    \I__11748\ : Span4Mux_h
    port map (
            O => \N__47630\,
            I => \N__47566\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__47627\,
            I => \N__47566\
        );

    \I__11746\ : Span4Mux_v
    port map (
            O => \N__47622\,
            I => \N__47566\
        );

    \I__11745\ : Span4Mux_h
    port map (
            O => \N__47613\,
            I => \N__47566\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__47608\,
            I => byte_transmit_counter_0
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__47599\,
            I => byte_transmit_counter_0
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__47596\,
            I => byte_transmit_counter_0
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__47591\,
            I => byte_transmit_counter_0
        );

    \I__11740\ : Odrv4
    port map (
            O => \N__47586\,
            I => byte_transmit_counter_0
        );

    \I__11739\ : Odrv4
    port map (
            O => \N__47583\,
            I => byte_transmit_counter_0
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__47580\,
            I => byte_transmit_counter_0
        );

    \I__11737\ : Odrv4
    port map (
            O => \N__47575\,
            I => byte_transmit_counter_0
        );

    \I__11736\ : Odrv4
    port map (
            O => \N__47566\,
            I => byte_transmit_counter_0
        );

    \I__11735\ : InMux
    port map (
            O => \N__47547\,
            I => \N__47543\
        );

    \I__11734\ : InMux
    port map (
            O => \N__47546\,
            I => \N__47540\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__47543\,
            I => \N__47537\
        );

    \I__11732\ : LocalMux
    port map (
            O => \N__47540\,
            I => \N__47533\
        );

    \I__11731\ : Span4Mux_h
    port map (
            O => \N__47537\,
            I => \N__47530\
        );

    \I__11730\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47527\
        );

    \I__11729\ : Span4Mux_h
    port map (
            O => \N__47533\,
            I => \N__47524\
        );

    \I__11728\ : Odrv4
    port map (
            O => \N__47530\,
            I => \c0.data_out_10_4\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__47527\,
            I => \c0.data_out_10_4\
        );

    \I__11726\ : Odrv4
    port map (
            O => \N__47524\,
            I => \c0.data_out_10_4\
        );

    \I__11725\ : CascadeMux
    port map (
            O => \N__47517\,
            I => \c0.n8_adj_2198_cascade_\
        );

    \I__11724\ : InMux
    port map (
            O => \N__47514\,
            I => \N__47510\
        );

    \I__11723\ : InMux
    port map (
            O => \N__47513\,
            I => \N__47504\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__47510\,
            I => \N__47501\
        );

    \I__11721\ : InMux
    port map (
            O => \N__47509\,
            I => \N__47498\
        );

    \I__11720\ : InMux
    port map (
            O => \N__47508\,
            I => \N__47489\
        );

    \I__11719\ : InMux
    port map (
            O => \N__47507\,
            I => \N__47489\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__47504\,
            I => \N__47478\
        );

    \I__11717\ : Span4Mux_v
    port map (
            O => \N__47501\,
            I => \N__47473\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__47498\,
            I => \N__47473\
        );

    \I__11715\ : InMux
    port map (
            O => \N__47497\,
            I => \N__47470\
        );

    \I__11714\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47465\
        );

    \I__11713\ : InMux
    port map (
            O => \N__47495\,
            I => \N__47465\
        );

    \I__11712\ : InMux
    port map (
            O => \N__47494\,
            I => \N__47462\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__47489\,
            I => \N__47459\
        );

    \I__11710\ : InMux
    port map (
            O => \N__47488\,
            I => \N__47455\
        );

    \I__11709\ : InMux
    port map (
            O => \N__47487\,
            I => \N__47451\
        );

    \I__11708\ : InMux
    port map (
            O => \N__47486\,
            I => \N__47448\
        );

    \I__11707\ : InMux
    port map (
            O => \N__47485\,
            I => \N__47445\
        );

    \I__11706\ : InMux
    port map (
            O => \N__47484\,
            I => \N__47442\
        );

    \I__11705\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47439\
        );

    \I__11704\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47435\
        );

    \I__11703\ : InMux
    port map (
            O => \N__47481\,
            I => \N__47432\
        );

    \I__11702\ : Span4Mux_v
    port map (
            O => \N__47478\,
            I => \N__47428\
        );

    \I__11701\ : Span4Mux_h
    port map (
            O => \N__47473\,
            I => \N__47423\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__47470\,
            I => \N__47423\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__47465\,
            I => \N__47416\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__47462\,
            I => \N__47416\
        );

    \I__11697\ : Span4Mux_s2_v
    port map (
            O => \N__47459\,
            I => \N__47416\
        );

    \I__11696\ : InMux
    port map (
            O => \N__47458\,
            I => \N__47413\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__47455\,
            I => \N__47410\
        );

    \I__11694\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47407\
        );

    \I__11693\ : LocalMux
    port map (
            O => \N__47451\,
            I => \N__47404\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47395\
        );

    \I__11691\ : LocalMux
    port map (
            O => \N__47445\,
            I => \N__47395\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__47442\,
            I => \N__47395\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__47439\,
            I => \N__47395\
        );

    \I__11688\ : InMux
    port map (
            O => \N__47438\,
            I => \N__47392\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__47435\,
            I => \N__47387\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__47432\,
            I => \N__47387\
        );

    \I__11685\ : InMux
    port map (
            O => \N__47431\,
            I => \N__47384\
        );

    \I__11684\ : Span4Mux_h
    port map (
            O => \N__47428\,
            I => \N__47379\
        );

    \I__11683\ : Span4Mux_v
    port map (
            O => \N__47423\,
            I => \N__47379\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__47416\,
            I => \N__47376\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__47413\,
            I => \N__47365\
        );

    \I__11680\ : Span4Mux_v
    port map (
            O => \N__47410\,
            I => \N__47365\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__47407\,
            I => \N__47365\
        );

    \I__11678\ : Span4Mux_h
    port map (
            O => \N__47404\,
            I => \N__47365\
        );

    \I__11677\ : Span4Mux_v
    port map (
            O => \N__47395\,
            I => \N__47365\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__47392\,
            I => byte_transmit_counter_1
        );

    \I__11675\ : Odrv12
    port map (
            O => \N__47387\,
            I => byte_transmit_counter_1
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__47384\,
            I => byte_transmit_counter_1
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__47379\,
            I => byte_transmit_counter_1
        );

    \I__11672\ : Odrv4
    port map (
            O => \N__47376\,
            I => byte_transmit_counter_1
        );

    \I__11671\ : Odrv4
    port map (
            O => \N__47365\,
            I => byte_transmit_counter_1
        );

    \I__11670\ : CascadeMux
    port map (
            O => \N__47352\,
            I => \N__47349\
        );

    \I__11669\ : InMux
    port map (
            O => \N__47349\,
            I => \N__47346\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__47346\,
            I => \N__47343\
        );

    \I__11667\ : Span12Mux_h
    port map (
            O => \N__47343\,
            I => \N__47340\
        );

    \I__11666\ : Odrv12
    port map (
            O => \N__47340\,
            I => n10_adj_2430
        );

    \I__11665\ : InMux
    port map (
            O => \N__47337\,
            I => \N__47334\
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__47334\,
            I => \c0.n17209\
        );

    \I__11663\ : InMux
    port map (
            O => \N__47331\,
            I => \N__47328\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__47328\,
            I => \c0.n17297\
        );

    \I__11661\ : CascadeMux
    port map (
            O => \N__47325\,
            I => \c0.n17297_cascade_\
        );

    \I__11660\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47317\
        );

    \I__11659\ : InMux
    port map (
            O => \N__47321\,
            I => \N__47314\
        );

    \I__11658\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47310\
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__47317\,
            I => \N__47307\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__47314\,
            I => \N__47304\
        );

    \I__11655\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47301\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__47310\,
            I => \N__47297\
        );

    \I__11653\ : Span4Mux_h
    port map (
            O => \N__47307\,
            I => \N__47294\
        );

    \I__11652\ : Span4Mux_h
    port map (
            O => \N__47304\,
            I => \N__47289\
        );

    \I__11651\ : LocalMux
    port map (
            O => \N__47301\,
            I => \N__47289\
        );

    \I__11650\ : InMux
    port map (
            O => \N__47300\,
            I => \N__47286\
        );

    \I__11649\ : Odrv4
    port map (
            O => \N__47297\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__11648\ : Odrv4
    port map (
            O => \N__47294\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__11647\ : Odrv4
    port map (
            O => \N__47289\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__47286\,
            I => \c0.data_out_7__2__N_447\
        );

    \I__11645\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47274\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__47274\,
            I => \N__47271\
        );

    \I__11643\ : Span4Mux_h
    port map (
            O => \N__47271\,
            I => \N__47268\
        );

    \I__11642\ : Odrv4
    port map (
            O => \N__47268\,
            I => \c0.n14_adj_2176\
        );

    \I__11641\ : InMux
    port map (
            O => \N__47265\,
            I => \N__47260\
        );

    \I__11640\ : InMux
    port map (
            O => \N__47264\,
            I => \N__47257\
        );

    \I__11639\ : InMux
    port map (
            O => \N__47263\,
            I => \N__47253\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__47260\,
            I => \N__47250\
        );

    \I__11637\ : LocalMux
    port map (
            O => \N__47257\,
            I => \N__47247\
        );

    \I__11636\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47244\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__47253\,
            I => \N__47241\
        );

    \I__11634\ : Span4Mux_v
    port map (
            O => \N__47250\,
            I => \N__47234\
        );

    \I__11633\ : Span4Mux_h
    port map (
            O => \N__47247\,
            I => \N__47234\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__47244\,
            I => \N__47234\
        );

    \I__11631\ : Span4Mux_h
    port map (
            O => \N__47241\,
            I => \N__47231\
        );

    \I__11630\ : Span4Mux_v
    port map (
            O => \N__47234\,
            I => \N__47227\
        );

    \I__11629\ : Span4Mux_h
    port map (
            O => \N__47231\,
            I => \N__47224\
        );

    \I__11628\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47221\
        );

    \I__11627\ : Span4Mux_s2_v
    port map (
            O => \N__47227\,
            I => \N__47218\
        );

    \I__11626\ : Odrv4
    port map (
            O => \N__47224\,
            I => \c0.data_out_7_6\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__47221\,
            I => \c0.data_out_7_6\
        );

    \I__11624\ : Odrv4
    port map (
            O => \N__47218\,
            I => \c0.data_out_7_6\
        );

    \I__11623\ : CascadeMux
    port map (
            O => \N__47211\,
            I => \N__47208\
        );

    \I__11622\ : InMux
    port map (
            O => \N__47208\,
            I => \N__47205\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__47205\,
            I => \N__47202\
        );

    \I__11620\ : Odrv4
    port map (
            O => \N__47202\,
            I => \c0.n12_adj_2180\
        );

    \I__11619\ : CascadeMux
    port map (
            O => \N__47199\,
            I => \N__47196\
        );

    \I__11618\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47191\
        );

    \I__11617\ : CascadeMux
    port map (
            O => \N__47195\,
            I => \N__47188\
        );

    \I__11616\ : CascadeMux
    port map (
            O => \N__47194\,
            I => \N__47185\
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__47191\,
            I => \N__47182\
        );

    \I__11614\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47179\
        );

    \I__11613\ : InMux
    port map (
            O => \N__47185\,
            I => \N__47176\
        );

    \I__11612\ : Span4Mux_v
    port map (
            O => \N__47182\,
            I => \N__47173\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__47179\,
            I => \N__47168\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__47176\,
            I => \N__47168\
        );

    \I__11609\ : Odrv4
    port map (
            O => \N__47173\,
            I => data_out_10_0
        );

    \I__11608\ : Odrv4
    port map (
            O => \N__47168\,
            I => data_out_10_0
        );

    \I__11607\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47157\
        );

    \I__11606\ : InMux
    port map (
            O => \N__47162\,
            I => \N__47157\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__47157\,
            I => \N__47153\
        );

    \I__11604\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47150\
        );

    \I__11603\ : Span12Mux_h
    port map (
            O => \N__47153\,
            I => \N__47147\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__47150\,
            I => \N__47144\
        );

    \I__11601\ : Span12Mux_h
    port map (
            O => \N__47147\,
            I => \N__47141\
        );

    \I__11600\ : Span12Mux_v
    port map (
            O => \N__47144\,
            I => \N__47138\
        );

    \I__11599\ : Odrv12
    port map (
            O => \N__47141\,
            I => \c0.data_out_7_3\
        );

    \I__11598\ : Odrv12
    port map (
            O => \N__47138\,
            I => \c0.data_out_7_3\
        );

    \I__11597\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47128\
        );

    \I__11596\ : InMux
    port map (
            O => \N__47132\,
            I => \N__47125\
        );

    \I__11595\ : InMux
    port map (
            O => \N__47131\,
            I => \N__47121\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__47128\,
            I => \N__47116\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__47125\,
            I => \N__47113\
        );

    \I__11592\ : InMux
    port map (
            O => \N__47124\,
            I => \N__47110\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__47121\,
            I => \N__47107\
        );

    \I__11590\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47103\
        );

    \I__11589\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47100\
        );

    \I__11588\ : Span4Mux_v
    port map (
            O => \N__47116\,
            I => \N__47097\
        );

    \I__11587\ : Span4Mux_v
    port map (
            O => \N__47113\,
            I => \N__47092\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__47110\,
            I => \N__47092\
        );

    \I__11585\ : Span4Mux_v
    port map (
            O => \N__47107\,
            I => \N__47089\
        );

    \I__11584\ : InMux
    port map (
            O => \N__47106\,
            I => \N__47086\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__47103\,
            I => \N__47082\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__47100\,
            I => \N__47075\
        );

    \I__11581\ : Span4Mux_h
    port map (
            O => \N__47097\,
            I => \N__47075\
        );

    \I__11580\ : Span4Mux_h
    port map (
            O => \N__47092\,
            I => \N__47075\
        );

    \I__11579\ : Sp12to4
    port map (
            O => \N__47089\,
            I => \N__47070\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__47086\,
            I => \N__47070\
        );

    \I__11577\ : InMux
    port map (
            O => \N__47085\,
            I => \N__47067\
        );

    \I__11576\ : Odrv4
    port map (
            O => \N__47082\,
            I => \c0.data_out_5_3\
        );

    \I__11575\ : Odrv4
    port map (
            O => \N__47075\,
            I => \c0.data_out_5_3\
        );

    \I__11574\ : Odrv12
    port map (
            O => \N__47070\,
            I => \c0.data_out_5_3\
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__47067\,
            I => \c0.data_out_5_3\
        );

    \I__11572\ : InMux
    port map (
            O => \N__47058\,
            I => \N__47055\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__47052\
        );

    \I__11570\ : Odrv4
    port map (
            O => \N__47052\,
            I => \c0.n17180\
        );

    \I__11569\ : InMux
    port map (
            O => \N__47049\,
            I => \N__47045\
        );

    \I__11568\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47042\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__47045\,
            I => \N__47039\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__47042\,
            I => \N__47035\
        );

    \I__11565\ : Span4Mux_h
    port map (
            O => \N__47039\,
            I => \N__47032\
        );

    \I__11564\ : InMux
    port map (
            O => \N__47038\,
            I => \N__47029\
        );

    \I__11563\ : Span4Mux_h
    port map (
            O => \N__47035\,
            I => \N__47026\
        );

    \I__11562\ : Odrv4
    port map (
            O => \N__47032\,
            I => \c0.data_out_9_4\
        );

    \I__11561\ : LocalMux
    port map (
            O => \N__47029\,
            I => \c0.data_out_9_4\
        );

    \I__11560\ : Odrv4
    port map (
            O => \N__47026\,
            I => \c0.data_out_9_4\
        );

    \I__11559\ : CascadeMux
    port map (
            O => \N__47019\,
            I => \c0.n17162_cascade_\
        );

    \I__11558\ : InMux
    port map (
            O => \N__47016\,
            I => \N__47010\
        );

    \I__11557\ : InMux
    port map (
            O => \N__47015\,
            I => \N__47007\
        );

    \I__11556\ : InMux
    port map (
            O => \N__47014\,
            I => \N__47004\
        );

    \I__11555\ : InMux
    port map (
            O => \N__47013\,
            I => \N__47001\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__47010\,
            I => \N__46998\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__47007\,
            I => \N__46994\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__47004\,
            I => \N__46991\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__47001\,
            I => \N__46986\
        );

    \I__11550\ : Span4Mux_v
    port map (
            O => \N__46998\,
            I => \N__46986\
        );

    \I__11549\ : InMux
    port map (
            O => \N__46997\,
            I => \N__46983\
        );

    \I__11548\ : Span12Mux_v
    port map (
            O => \N__46994\,
            I => \N__46980\
        );

    \I__11547\ : Span4Mux_v
    port map (
            O => \N__46991\,
            I => \N__46977\
        );

    \I__11546\ : Span4Mux_h
    port map (
            O => \N__46986\,
            I => \N__46972\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__46983\,
            I => \N__46972\
        );

    \I__11544\ : Odrv12
    port map (
            O => \N__46980\,
            I => \c0.data_out_6_2\
        );

    \I__11543\ : Odrv4
    port map (
            O => \N__46977\,
            I => \c0.data_out_6_2\
        );

    \I__11542\ : Odrv4
    port map (
            O => \N__46972\,
            I => \c0.data_out_6_2\
        );

    \I__11541\ : CascadeMux
    port map (
            O => \N__46965\,
            I => \N__46962\
        );

    \I__11540\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46959\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__46959\,
            I => \N__46955\
        );

    \I__11538\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46952\
        );

    \I__11537\ : Odrv4
    port map (
            O => \N__46955\,
            I => \c0.n17197\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__46952\,
            I => \c0.n17197\
        );

    \I__11535\ : CascadeMux
    port map (
            O => \N__46947\,
            I => \c0.n10_adj_2196_cascade_\
        );

    \I__11534\ : InMux
    port map (
            O => \N__46944\,
            I => \N__46938\
        );

    \I__11533\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46938\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__46938\,
            I => \c0.n17261\
        );

    \I__11531\ : CEMux
    port map (
            O => \N__46935\,
            I => \N__46930\
        );

    \I__11530\ : CEMux
    port map (
            O => \N__46934\,
            I => \N__46927\
        );

    \I__11529\ : CEMux
    port map (
            O => \N__46933\,
            I => \N__46924\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__46930\,
            I => \N__46919\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__46927\,
            I => \N__46915\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__46924\,
            I => \N__46912\
        );

    \I__11525\ : CEMux
    port map (
            O => \N__46923\,
            I => \N__46909\
        );

    \I__11524\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46906\
        );

    \I__11523\ : Span4Mux_s3_h
    port map (
            O => \N__46919\,
            I => \N__46902\
        );

    \I__11522\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46899\
        );

    \I__11521\ : Span4Mux_h
    port map (
            O => \N__46915\,
            I => \N__46895\
        );

    \I__11520\ : Span4Mux_v
    port map (
            O => \N__46912\,
            I => \N__46890\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__46909\,
            I => \N__46890\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__46906\,
            I => \N__46887\
        );

    \I__11517\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46884\
        );

    \I__11516\ : Span4Mux_h
    port map (
            O => \N__46902\,
            I => \N__46881\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__46899\,
            I => \N__46878\
        );

    \I__11514\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46875\
        );

    \I__11513\ : Span4Mux_v
    port map (
            O => \N__46895\,
            I => \N__46870\
        );

    \I__11512\ : Span4Mux_h
    port map (
            O => \N__46890\,
            I => \N__46870\
        );

    \I__11511\ : Span4Mux_v
    port map (
            O => \N__46887\,
            I => \N__46867\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__46884\,
            I => \N__46864\
        );

    \I__11509\ : Span4Mux_h
    port map (
            O => \N__46881\,
            I => \N__46859\
        );

    \I__11508\ : Span4Mux_v
    port map (
            O => \N__46878\,
            I => \N__46859\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__46875\,
            I => \N__46856\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__46870\,
            I => \N__46853\
        );

    \I__11505\ : Span4Mux_h
    port map (
            O => \N__46867\,
            I => \N__46850\
        );

    \I__11504\ : Span12Mux_h
    port map (
            O => \N__46864\,
            I => \N__46847\
        );

    \I__11503\ : Span4Mux_h
    port map (
            O => \N__46859\,
            I => \N__46842\
        );

    \I__11502\ : Span4Mux_v
    port map (
            O => \N__46856\,
            I => \N__46842\
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__46853\,
            I => \c0.n10595\
        );

    \I__11500\ : Odrv4
    port map (
            O => \N__46850\,
            I => \c0.n10595\
        );

    \I__11499\ : Odrv12
    port map (
            O => \N__46847\,
            I => \c0.n10595\
        );

    \I__11498\ : Odrv4
    port map (
            O => \N__46842\,
            I => \c0.n10595\
        );

    \I__11497\ : InMux
    port map (
            O => \N__46833\,
            I => \N__46829\
        );

    \I__11496\ : CascadeMux
    port map (
            O => \N__46832\,
            I => \N__46826\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__46829\,
            I => \N__46821\
        );

    \I__11494\ : InMux
    port map (
            O => \N__46826\,
            I => \N__46818\
        );

    \I__11493\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46814\
        );

    \I__11492\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46811\
        );

    \I__11491\ : Span4Mux_v
    port map (
            O => \N__46821\,
            I => \N__46806\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__46818\,
            I => \N__46806\
        );

    \I__11489\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46803\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__46814\,
            I => \N__46798\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__46811\,
            I => \N__46798\
        );

    \I__11486\ : Span4Mux_h
    port map (
            O => \N__46806\,
            I => \N__46795\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__46803\,
            I => \c0.data_out_6_0\
        );

    \I__11484\ : Odrv12
    port map (
            O => \N__46798\,
            I => \c0.data_out_6_0\
        );

    \I__11483\ : Odrv4
    port map (
            O => \N__46795\,
            I => \c0.data_out_6_0\
        );

    \I__11482\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46785\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46781\
        );

    \I__11480\ : InMux
    port map (
            O => \N__46784\,
            I => \N__46778\
        );

    \I__11479\ : Odrv4
    port map (
            O => \N__46781\,
            I => \c0.n17129\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__46778\,
            I => \c0.n17129\
        );

    \I__11477\ : CascadeMux
    port map (
            O => \N__46773\,
            I => \c0.n10447_cascade_\
        );

    \I__11476\ : InMux
    port map (
            O => \N__46770\,
            I => \N__46767\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46763\
        );

    \I__11474\ : InMux
    port map (
            O => \N__46766\,
            I => \N__46760\
        );

    \I__11473\ : Span4Mux_v
    port map (
            O => \N__46763\,
            I => \N__46754\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__46760\,
            I => \N__46754\
        );

    \I__11471\ : InMux
    port map (
            O => \N__46759\,
            I => \N__46751\
        );

    \I__11470\ : Span4Mux_h
    port map (
            O => \N__46754\,
            I => \N__46747\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__46751\,
            I => \N__46744\
        );

    \I__11468\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46741\
        );

    \I__11467\ : Odrv4
    port map (
            O => \N__46747\,
            I => \c0.data_out_6_1\
        );

    \I__11466\ : Odrv4
    port map (
            O => \N__46744\,
            I => \c0.data_out_6_1\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__46741\,
            I => \c0.data_out_6_1\
        );

    \I__11464\ : CascadeMux
    port map (
            O => \N__46734\,
            I => \N__46731\
        );

    \I__11463\ : InMux
    port map (
            O => \N__46731\,
            I => \N__46728\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__46728\,
            I => \N__46723\
        );

    \I__11461\ : InMux
    port map (
            O => \N__46727\,
            I => \N__46720\
        );

    \I__11460\ : InMux
    port map (
            O => \N__46726\,
            I => \N__46717\
        );

    \I__11459\ : Span4Mux_h
    port map (
            O => \N__46723\,
            I => \N__46714\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46711\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__46717\,
            I => \c0.n10183\
        );

    \I__11456\ : Odrv4
    port map (
            O => \N__46714\,
            I => \c0.n10183\
        );

    \I__11455\ : Odrv12
    port map (
            O => \N__46711\,
            I => \c0.n10183\
        );

    \I__11454\ : InMux
    port map (
            O => \N__46704\,
            I => \N__46700\
        );

    \I__11453\ : InMux
    port map (
            O => \N__46703\,
            I => \N__46697\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__46700\,
            I => \N__46690\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__46697\,
            I => \N__46690\
        );

    \I__11450\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46687\
        );

    \I__11449\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46684\
        );

    \I__11448\ : Span4Mux_v
    port map (
            O => \N__46690\,
            I => \N__46681\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__46687\,
            I => \N__46678\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__46684\,
            I => \N__46675\
        );

    \I__11445\ : Span4Mux_h
    port map (
            O => \N__46681\,
            I => \N__46670\
        );

    \I__11444\ : Span4Mux_v
    port map (
            O => \N__46678\,
            I => \N__46670\
        );

    \I__11443\ : Span4Mux_h
    port map (
            O => \N__46675\,
            I => \N__46667\
        );

    \I__11442\ : Odrv4
    port map (
            O => \N__46670\,
            I => \c0.data_out_6_3\
        );

    \I__11441\ : Odrv4
    port map (
            O => \N__46667\,
            I => \c0.data_out_6_3\
        );

    \I__11440\ : CascadeMux
    port map (
            O => \N__46662\,
            I => \N__46659\
        );

    \I__11439\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46655\
        );

    \I__11438\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46652\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__46655\,
            I => \c0.n17222\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__46652\,
            I => \c0.n17222\
        );

    \I__11435\ : CascadeMux
    port map (
            O => \N__46647\,
            I => \N__46643\
        );

    \I__11434\ : CascadeMux
    port map (
            O => \N__46646\,
            I => \N__46640\
        );

    \I__11433\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46637\
        );

    \I__11432\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46634\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__46637\,
            I => \N__46631\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__46634\,
            I => \N__46628\
        );

    \I__11429\ : Span4Mux_v
    port map (
            O => \N__46631\,
            I => \N__46623\
        );

    \I__11428\ : Span4Mux_h
    port map (
            O => \N__46628\,
            I => \N__46620\
        );

    \I__11427\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46617\
        );

    \I__11426\ : InMux
    port map (
            O => \N__46626\,
            I => \N__46614\
        );

    \I__11425\ : Span4Mux_h
    port map (
            O => \N__46623\,
            I => \N__46611\
        );

    \I__11424\ : Sp12to4
    port map (
            O => \N__46620\,
            I => \N__46606\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46606\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__46614\,
            I => \c0.data_out_9_7\
        );

    \I__11421\ : Odrv4
    port map (
            O => \N__46611\,
            I => \c0.data_out_9_7\
        );

    \I__11420\ : Odrv12
    port map (
            O => \N__46606\,
            I => \c0.data_out_9_7\
        );

    \I__11419\ : CascadeMux
    port map (
            O => \N__46599\,
            I => \N__46596\
        );

    \I__11418\ : InMux
    port map (
            O => \N__46596\,
            I => \N__46593\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__46593\,
            I => \N__46590\
        );

    \I__11416\ : Span4Mux_h
    port map (
            O => \N__46590\,
            I => \N__46586\
        );

    \I__11415\ : InMux
    port map (
            O => \N__46589\,
            I => \N__46583\
        );

    \I__11414\ : Odrv4
    port map (
            O => \N__46586\,
            I => \c0.n17243\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__46583\,
            I => \c0.n17243\
        );

    \I__11412\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46575\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__46575\,
            I => \N__46571\
        );

    \I__11410\ : InMux
    port map (
            O => \N__46574\,
            I => \N__46568\
        );

    \I__11409\ : Span4Mux_h
    port map (
            O => \N__46571\,
            I => \N__46565\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__46568\,
            I => \N__46562\
        );

    \I__11407\ : Span4Mux_h
    port map (
            O => \N__46565\,
            I => \N__46559\
        );

    \I__11406\ : Odrv12
    port map (
            O => \N__46562\,
            I => \c0.n17264\
        );

    \I__11405\ : Odrv4
    port map (
            O => \N__46559\,
            I => \c0.n17264\
        );

    \I__11404\ : CascadeMux
    port map (
            O => \N__46554\,
            I => \c0.n10_adj_2191_cascade_\
        );

    \I__11403\ : InMux
    port map (
            O => \N__46551\,
            I => \N__46548\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__46548\,
            I => \N__46543\
        );

    \I__11401\ : InMux
    port map (
            O => \N__46547\,
            I => \N__46540\
        );

    \I__11400\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46537\
        );

    \I__11399\ : Odrv4
    port map (
            O => \N__46543\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__46540\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__46537\,
            I => \c0.tx.r_Clock_Count_7\
        );

    \I__11396\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46526\
        );

    \I__11395\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46523\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__46526\,
            I => data_out_3_7
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__46523\,
            I => data_out_3_7
        );

    \I__11392\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46512\
        );

    \I__11391\ : InMux
    port map (
            O => \N__46517\,
            I => \N__46512\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__46512\,
            I => data_out_2_7
        );

    \I__11389\ : InMux
    port map (
            O => \N__46509\,
            I => \N__46503\
        );

    \I__11388\ : InMux
    port map (
            O => \N__46508\,
            I => \N__46500\
        );

    \I__11387\ : InMux
    port map (
            O => \N__46507\,
            I => \N__46497\
        );

    \I__11386\ : InMux
    port map (
            O => \N__46506\,
            I => \N__46494\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__46503\,
            I => \N__46491\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__46500\,
            I => \N__46488\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__46497\,
            I => \N__46483\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__46494\,
            I => \N__46483\
        );

    \I__11381\ : Span4Mux_v
    port map (
            O => \N__46491\,
            I => \N__46480\
        );

    \I__11380\ : Span4Mux_v
    port map (
            O => \N__46488\,
            I => \N__46477\
        );

    \I__11379\ : Span12Mux_h
    port map (
            O => \N__46483\,
            I => \N__46473\
        );

    \I__11378\ : Span4Mux_h
    port map (
            O => \N__46480\,
            I => \N__46470\
        );

    \I__11377\ : Span4Mux_h
    port map (
            O => \N__46477\,
            I => \N__46467\
        );

    \I__11376\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46464\
        );

    \I__11375\ : Span12Mux_h
    port map (
            O => \N__46473\,
            I => \N__46461\
        );

    \I__11374\ : Sp12to4
    port map (
            O => \N__46470\,
            I => \N__46456\
        );

    \I__11373\ : Sp12to4
    port map (
            O => \N__46467\,
            I => \N__46456\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__46464\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__11371\ : Odrv12
    port map (
            O => \N__46461\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__11370\ : Odrv12
    port map (
            O => \N__46456\,
            I => \c0.data_out_7__3__N_441\
        );

    \I__11369\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46446\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__46446\,
            I => \N__46443\
        );

    \I__11367\ : Span4Mux_v
    port map (
            O => \N__46443\,
            I => \N__46440\
        );

    \I__11366\ : Odrv4
    port map (
            O => \N__46440\,
            I => \c0.n1\
        );

    \I__11365\ : CascadeMux
    port map (
            O => \N__46437\,
            I => \c0.n17747_cascade_\
        );

    \I__11364\ : InMux
    port map (
            O => \N__46434\,
            I => \N__46431\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__46431\,
            I => \c0.n2_adj_2156\
        );

    \I__11362\ : CascadeMux
    port map (
            O => \N__46428\,
            I => \c0.n18220_cascade_\
        );

    \I__11361\ : InMux
    port map (
            O => \N__46425\,
            I => \N__46422\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__46422\,
            I => \N__46419\
        );

    \I__11359\ : Odrv12
    port map (
            O => \N__46419\,
            I => \c0.n17607\
        );

    \I__11358\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46410\
        );

    \I__11357\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46407\
        );

    \I__11356\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46404\
        );

    \I__11355\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46397\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__46410\,
            I => \N__46392\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__46407\,
            I => \N__46392\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__46404\,
            I => \N__46389\
        );

    \I__11351\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46386\
        );

    \I__11350\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46383\
        );

    \I__11349\ : InMux
    port map (
            O => \N__46401\,
            I => \N__46380\
        );

    \I__11348\ : InMux
    port map (
            O => \N__46400\,
            I => \N__46376\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__46397\,
            I => \N__46372\
        );

    \I__11346\ : Span4Mux_v
    port map (
            O => \N__46392\,
            I => \N__46369\
        );

    \I__11345\ : Span4Mux_s2_v
    port map (
            O => \N__46389\,
            I => \N__46360\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__46386\,
            I => \N__46360\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__46383\,
            I => \N__46360\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__46380\,
            I => \N__46360\
        );

    \I__11341\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46357\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__46376\,
            I => \N__46354\
        );

    \I__11339\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46351\
        );

    \I__11338\ : Span4Mux_v
    port map (
            O => \N__46372\,
            I => \N__46346\
        );

    \I__11337\ : Span4Mux_h
    port map (
            O => \N__46369\,
            I => \N__46346\
        );

    \I__11336\ : Span4Mux_v
    port map (
            O => \N__46360\,
            I => \N__46343\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__46357\,
            I => byte_transmit_counter_3
        );

    \I__11334\ : Odrv12
    port map (
            O => \N__46354\,
            I => byte_transmit_counter_3
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__46351\,
            I => byte_transmit_counter_3
        );

    \I__11332\ : Odrv4
    port map (
            O => \N__46346\,
            I => byte_transmit_counter_3
        );

    \I__11331\ : Odrv4
    port map (
            O => \N__46343\,
            I => byte_transmit_counter_3
        );

    \I__11330\ : InMux
    port map (
            O => \N__46332\,
            I => \N__46329\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__46329\,
            I => n10_adj_2413
        );

    \I__11328\ : CascadeMux
    port map (
            O => \N__46326\,
            I => \n18223_cascade_\
        );

    \I__11327\ : InMux
    port map (
            O => \N__46323\,
            I => \N__46316\
        );

    \I__11326\ : InMux
    port map (
            O => \N__46322\,
            I => \N__46316\
        );

    \I__11325\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46310\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__46316\,
            I => \N__46307\
        );

    \I__11323\ : InMux
    port map (
            O => \N__46315\,
            I => \N__46300\
        );

    \I__11322\ : InMux
    port map (
            O => \N__46314\,
            I => \N__46300\
        );

    \I__11321\ : InMux
    port map (
            O => \N__46313\,
            I => \N__46300\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__46310\,
            I => \N__46285\
        );

    \I__11319\ : Span4Mux_h
    port map (
            O => \N__46307\,
            I => \N__46280\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__46300\,
            I => \N__46280\
        );

    \I__11317\ : InMux
    port map (
            O => \N__46299\,
            I => \N__46277\
        );

    \I__11316\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46274\
        );

    \I__11315\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46267\
        );

    \I__11314\ : InMux
    port map (
            O => \N__46296\,
            I => \N__46267\
        );

    \I__11313\ : InMux
    port map (
            O => \N__46295\,
            I => \N__46267\
        );

    \I__11312\ : InMux
    port map (
            O => \N__46294\,
            I => \N__46262\
        );

    \I__11311\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46262\
        );

    \I__11310\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46259\
        );

    \I__11309\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46256\
        );

    \I__11308\ : InMux
    port map (
            O => \N__46290\,
            I => \N__46247\
        );

    \I__11307\ : InMux
    port map (
            O => \N__46289\,
            I => \N__46244\
        );

    \I__11306\ : InMux
    port map (
            O => \N__46288\,
            I => \N__46241\
        );

    \I__11305\ : Span4Mux_s1_v
    port map (
            O => \N__46285\,
            I => \N__46234\
        );

    \I__11304\ : Span4Mux_v
    port map (
            O => \N__46280\,
            I => \N__46234\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__46277\,
            I => \N__46234\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__46274\,
            I => \N__46227\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__46267\,
            I => \N__46227\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__46262\,
            I => \N__46227\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__46259\,
            I => \N__46222\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__46256\,
            I => \N__46222\
        );

    \I__11297\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46219\
        );

    \I__11296\ : InMux
    port map (
            O => \N__46254\,
            I => \N__46216\
        );

    \I__11295\ : InMux
    port map (
            O => \N__46253\,
            I => \N__46211\
        );

    \I__11294\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46211\
        );

    \I__11293\ : InMux
    port map (
            O => \N__46251\,
            I => \N__46206\
        );

    \I__11292\ : InMux
    port map (
            O => \N__46250\,
            I => \N__46206\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__46247\,
            I => \N__46201\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__46244\,
            I => \N__46201\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__46241\,
            I => \N__46196\
        );

    \I__11288\ : Span4Mux_h
    port map (
            O => \N__46234\,
            I => \N__46196\
        );

    \I__11287\ : Span4Mux_v
    port map (
            O => \N__46227\,
            I => \N__46191\
        );

    \I__11286\ : Span4Mux_s3_v
    port map (
            O => \N__46222\,
            I => \N__46191\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__46219\,
            I => byte_transmit_counter_2
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__46216\,
            I => byte_transmit_counter_2
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__46211\,
            I => byte_transmit_counter_2
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__46206\,
            I => byte_transmit_counter_2
        );

    \I__11281\ : Odrv4
    port map (
            O => \N__46201\,
            I => byte_transmit_counter_2
        );

    \I__11280\ : Odrv4
    port map (
            O => \N__46196\,
            I => byte_transmit_counter_2
        );

    \I__11279\ : Odrv4
    port map (
            O => \N__46191\,
            I => byte_transmit_counter_2
        );

    \I__11278\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46173\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__46173\,
            I => \N__46170\
        );

    \I__11276\ : Span4Mux_h
    port map (
            O => \N__46170\,
            I => \N__46167\
        );

    \I__11275\ : Odrv4
    port map (
            O => \N__46167\,
            I => n10
        );

    \I__11274\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46161\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__46161\,
            I => \N__46158\
        );

    \I__11272\ : Odrv4
    port map (
            O => \N__46158\,
            I => n10960
        );

    \I__11271\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46150\
        );

    \I__11270\ : InMux
    port map (
            O => \N__46154\,
            I => \N__46147\
        );

    \I__11269\ : InMux
    port map (
            O => \N__46153\,
            I => \N__46144\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__46150\,
            I => \N__46137\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__46147\,
            I => \N__46137\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__46144\,
            I => \N__46137\
        );

    \I__11265\ : Odrv4
    port map (
            O => \N__46137\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__11264\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46131\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__46131\,
            I => \N__46128\
        );

    \I__11262\ : Odrv12
    port map (
            O => \N__46128\,
            I => n10994
        );

    \I__11261\ : InMux
    port map (
            O => \N__46125\,
            I => \N__46112\
        );

    \I__11260\ : InMux
    port map (
            O => \N__46124\,
            I => \N__46112\
        );

    \I__11259\ : InMux
    port map (
            O => \N__46123\,
            I => \N__46112\
        );

    \I__11258\ : InMux
    port map (
            O => \N__46122\,
            I => \N__46106\
        );

    \I__11257\ : InMux
    port map (
            O => \N__46121\,
            I => \N__46106\
        );

    \I__11256\ : InMux
    port map (
            O => \N__46120\,
            I => \N__46101\
        );

    \I__11255\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46101\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__46112\,
            I => \N__46098\
        );

    \I__11253\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46095\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__46106\,
            I => n5142
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__46101\,
            I => n5142
        );

    \I__11250\ : Odrv4
    port map (
            O => \N__46098\,
            I => n5142
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__46095\,
            I => n5142
        );

    \I__11248\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46081\
        );

    \I__11247\ : InMux
    port map (
            O => \N__46085\,
            I => \N__46078\
        );

    \I__11246\ : InMux
    port map (
            O => \N__46084\,
            I => \N__46075\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__46081\,
            I => \N__46070\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__46078\,
            I => \N__46070\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46067\
        );

    \I__11242\ : Span4Mux_h
    port map (
            O => \N__46070\,
            I => \N__46062\
        );

    \I__11241\ : Span4Mux_h
    port map (
            O => \N__46067\,
            I => \N__46062\
        );

    \I__11240\ : Odrv4
    port map (
            O => \N__46062\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__11239\ : InMux
    port map (
            O => \N__46059\,
            I => \c0.tx.n16120\
        );

    \I__11238\ : InMux
    port map (
            O => \N__46056\,
            I => \N__46052\
        );

    \I__11237\ : InMux
    port map (
            O => \N__46055\,
            I => \N__46048\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__46052\,
            I => \N__46045\
        );

    \I__11235\ : InMux
    port map (
            O => \N__46051\,
            I => \N__46042\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__46048\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__11233\ : Odrv4
    port map (
            O => \N__46045\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__46042\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__11231\ : CascadeMux
    port map (
            O => \N__46035\,
            I => \N__46032\
        );

    \I__11230\ : InMux
    port map (
            O => \N__46032\,
            I => \N__46029\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__46029\,
            I => n10963
        );

    \I__11228\ : InMux
    port map (
            O => \N__46026\,
            I => \c0.tx.n16121\
        );

    \I__11227\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46018\
        );

    \I__11226\ : InMux
    port map (
            O => \N__46022\,
            I => \N__46015\
        );

    \I__11225\ : InMux
    port map (
            O => \N__46021\,
            I => \N__46012\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__46018\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__46015\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__46012\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__11221\ : InMux
    port map (
            O => \N__46005\,
            I => \N__46002\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__46002\,
            I => \N__45999\
        );

    \I__11219\ : Odrv4
    port map (
            O => \N__45999\,
            I => n10966
        );

    \I__11218\ : InMux
    port map (
            O => \N__45996\,
            I => \c0.tx.n16122\
        );

    \I__11217\ : InMux
    port map (
            O => \N__45993\,
            I => \c0.tx.n16123\
        );

    \I__11216\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45987\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__45987\,
            I => \N__45982\
        );

    \I__11214\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45979\
        );

    \I__11213\ : InMux
    port map (
            O => \N__45985\,
            I => \N__45976\
        );

    \I__11212\ : Span4Mux_h
    port map (
            O => \N__45982\,
            I => \N__45973\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__45979\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__45976\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__11209\ : Odrv4
    port map (
            O => \N__45973\,
            I => \c0.tx.r_Clock_Count_8\
        );

    \I__11208\ : CascadeMux
    port map (
            O => \N__45966\,
            I => \N__45955\
        );

    \I__11207\ : CascadeMux
    port map (
            O => \N__45965\,
            I => \N__45952\
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__45964\,
            I => \N__45949\
        );

    \I__11205\ : CascadeMux
    port map (
            O => \N__45963\,
            I => \N__45946\
        );

    \I__11204\ : CascadeMux
    port map (
            O => \N__45962\,
            I => \N__45942\
        );

    \I__11203\ : CascadeMux
    port map (
            O => \N__45961\,
            I => \N__45937\
        );

    \I__11202\ : CascadeMux
    port map (
            O => \N__45960\,
            I => \N__45934\
        );

    \I__11201\ : CascadeMux
    port map (
            O => \N__45959\,
            I => \N__45931\
        );

    \I__11200\ : CascadeMux
    port map (
            O => \N__45958\,
            I => \N__45928\
        );

    \I__11199\ : InMux
    port map (
            O => \N__45955\,
            I => \N__45915\
        );

    \I__11198\ : InMux
    port map (
            O => \N__45952\,
            I => \N__45915\
        );

    \I__11197\ : InMux
    port map (
            O => \N__45949\,
            I => \N__45915\
        );

    \I__11196\ : InMux
    port map (
            O => \N__45946\,
            I => \N__45915\
        );

    \I__11195\ : InMux
    port map (
            O => \N__45945\,
            I => \N__45912\
        );

    \I__11194\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45909\
        );

    \I__11193\ : InMux
    port map (
            O => \N__45941\,
            I => \N__45904\
        );

    \I__11192\ : InMux
    port map (
            O => \N__45940\,
            I => \N__45904\
        );

    \I__11191\ : InMux
    port map (
            O => \N__45937\,
            I => \N__45895\
        );

    \I__11190\ : InMux
    port map (
            O => \N__45934\,
            I => \N__45895\
        );

    \I__11189\ : InMux
    port map (
            O => \N__45931\,
            I => \N__45895\
        );

    \I__11188\ : InMux
    port map (
            O => \N__45928\,
            I => \N__45895\
        );

    \I__11187\ : InMux
    port map (
            O => \N__45927\,
            I => \N__45891\
        );

    \I__11186\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45884\
        );

    \I__11185\ : InMux
    port map (
            O => \N__45925\,
            I => \N__45884\
        );

    \I__11184\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45884\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__45915\,
            I => \N__45881\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__45912\,
            I => \N__45872\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__45909\,
            I => \N__45872\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__45904\,
            I => \N__45872\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__45895\,
            I => \N__45872\
        );

    \I__11178\ : InMux
    port map (
            O => \N__45894\,
            I => \N__45869\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__45891\,
            I => \N__45866\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__45884\,
            I => \N__45859\
        );

    \I__11175\ : Span4Mux_v
    port map (
            O => \N__45881\,
            I => \N__45859\
        );

    \I__11174\ : Span4Mux_v
    port map (
            O => \N__45872\,
            I => \N__45859\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__45869\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__11172\ : Odrv4
    port map (
            O => \N__45866\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__11171\ : Odrv4
    port map (
            O => \N__45859\,
            I => \c0.tx.r_SM_Main_2\
        );

    \I__11170\ : InMux
    port map (
            O => \N__45852\,
            I => \bfn_16_29_0_\
        );

    \I__11169\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45846\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__45846\,
            I => n10972
        );

    \I__11167\ : CascadeMux
    port map (
            O => \N__45843\,
            I => \N__45840\
        );

    \I__11166\ : InMux
    port map (
            O => \N__45840\,
            I => \N__45833\
        );

    \I__11165\ : InMux
    port map (
            O => \N__45839\,
            I => \N__45830\
        );

    \I__11164\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45827\
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__45837\,
            I => \N__45824\
        );

    \I__11162\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45821\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__45833\,
            I => \N__45818\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45813\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__45827\,
            I => \N__45813\
        );

    \I__11158\ : InMux
    port map (
            O => \N__45824\,
            I => \N__45810\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__45821\,
            I => \N__45807\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__45818\,
            I => \N__45802\
        );

    \I__11155\ : Span4Mux_h
    port map (
            O => \N__45813\,
            I => \N__45802\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__45810\,
            I => \N__45797\
        );

    \I__11153\ : Span4Mux_h
    port map (
            O => \N__45807\,
            I => \N__45797\
        );

    \I__11152\ : Odrv4
    port map (
            O => \N__45802\,
            I => data_out_8_7
        );

    \I__11151\ : Odrv4
    port map (
            O => \N__45797\,
            I => data_out_8_7
        );

    \I__11150\ : InMux
    port map (
            O => \N__45792\,
            I => \N__45789\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__45789\,
            I => n10951
        );

    \I__11148\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45781\
        );

    \I__11147\ : InMux
    port map (
            O => \N__45785\,
            I => \N__45778\
        );

    \I__11146\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45775\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__45781\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__45778\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__45775\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__11142\ : InMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45762\
        );

    \I__11140\ : Odrv4
    port map (
            O => \N__45762\,
            I => n10969
        );

    \I__11139\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__45756\,
            I => n32
        );

    \I__11137\ : CascadeMux
    port map (
            O => \N__45753\,
            I => \n29_cascade_\
        );

    \I__11136\ : InMux
    port map (
            O => \N__45750\,
            I => \N__45747\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__45747\,
            I => n26
        );

    \I__11134\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45740\
        );

    \I__11133\ : InMux
    port map (
            O => \N__45743\,
            I => \N__45737\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__45740\,
            I => \N__45734\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__45737\,
            I => \N__45729\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__45734\,
            I => \N__45724\
        );

    \I__11129\ : InMux
    port map (
            O => \N__45733\,
            I => \N__45719\
        );

    \I__11128\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45719\
        );

    \I__11127\ : Span12Mux_h
    port map (
            O => \N__45729\,
            I => \N__45716\
        );

    \I__11126\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45711\
        );

    \I__11125\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45711\
        );

    \I__11124\ : Span4Mux_h
    port map (
            O => \N__45724\,
            I => \N__45708\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__45719\,
            I => \N__45705\
        );

    \I__11122\ : Odrv12
    port map (
            O => \N__45716\,
            I => \c0.data_out_5_2\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__45711\,
            I => \c0.data_out_5_2\
        );

    \I__11120\ : Odrv4
    port map (
            O => \N__45708\,
            I => \c0.data_out_5_2\
        );

    \I__11119\ : Odrv4
    port map (
            O => \N__45705\,
            I => \c0.data_out_5_2\
        );

    \I__11118\ : CascadeMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__11117\ : InMux
    port map (
            O => \N__45693\,
            I => \N__45690\
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__45690\,
            I => \N__45687\
        );

    \I__11115\ : Span4Mux_h
    port map (
            O => \N__45687\,
            I => \N__45684\
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__45684\,
            I => \c0.n10196\
        );

    \I__11113\ : CascadeMux
    port map (
            O => \N__45681\,
            I => \c0.n10196_cascade_\
        );

    \I__11112\ : InMux
    port map (
            O => \N__45678\,
            I => \N__45675\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__45675\,
            I => \N__45672\
        );

    \I__11110\ : Span4Mux_v
    port map (
            O => \N__45672\,
            I => \N__45667\
        );

    \I__11109\ : InMux
    port map (
            O => \N__45671\,
            I => \N__45662\
        );

    \I__11108\ : InMux
    port map (
            O => \N__45670\,
            I => \N__45662\
        );

    \I__11107\ : Odrv4
    port map (
            O => \N__45667\,
            I => \c0.data_out_10_3\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__45662\,
            I => \c0.data_out_10_3\
        );

    \I__11105\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45653\
        );

    \I__11104\ : InMux
    port map (
            O => \N__45656\,
            I => \N__45650\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__45653\,
            I => \N__45647\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__45650\,
            I => \N__45643\
        );

    \I__11101\ : Span4Mux_h
    port map (
            O => \N__45647\,
            I => \N__45640\
        );

    \I__11100\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45637\
        );

    \I__11099\ : Span4Mux_h
    port map (
            O => \N__45643\,
            I => \N__45634\
        );

    \I__11098\ : Span4Mux_v
    port map (
            O => \N__45640\,
            I => \N__45631\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__45637\,
            I => \N__45626\
        );

    \I__11096\ : Span4Mux_h
    port map (
            O => \N__45634\,
            I => \N__45626\
        );

    \I__11095\ : Odrv4
    port map (
            O => \N__45631\,
            I => \c0.data_out_6_4\
        );

    \I__11094\ : Odrv4
    port map (
            O => \N__45626\,
            I => \c0.data_out_6_4\
        );

    \I__11093\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45617\
        );

    \I__11092\ : InMux
    port map (
            O => \N__45620\,
            I => \N__45611\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__45617\,
            I => \N__45608\
        );

    \I__11090\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45605\
        );

    \I__11089\ : InMux
    port map (
            O => \N__45615\,
            I => \N__45600\
        );

    \I__11088\ : InMux
    port map (
            O => \N__45614\,
            I => \N__45600\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__45611\,
            I => data_out_8_5
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__45608\,
            I => data_out_8_5
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__45605\,
            I => data_out_8_5
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__45600\,
            I => data_out_8_5
        );

    \I__11083\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45587\
        );

    \I__11082\ : InMux
    port map (
            O => \N__45590\,
            I => \N__45584\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__45587\,
            I => \N__45579\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45579\
        );

    \I__11079\ : Odrv12
    port map (
            O => \N__45579\,
            I => \c0.n10392\
        );

    \I__11078\ : InMux
    port map (
            O => \N__45576\,
            I => \bfn_16_28_0_\
        );

    \I__11077\ : InMux
    port map (
            O => \N__45573\,
            I => \c0.tx.n16117\
        );

    \I__11076\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45565\
        );

    \I__11075\ : InMux
    port map (
            O => \N__45569\,
            I => \N__45562\
        );

    \I__11074\ : InMux
    port map (
            O => \N__45568\,
            I => \N__45559\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__45565\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__45562\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__45559\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__11070\ : InMux
    port map (
            O => \N__45552\,
            I => \N__45549\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__45549\,
            I => n10954
        );

    \I__11068\ : InMux
    port map (
            O => \N__45546\,
            I => \c0.tx.n16118\
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__45543\,
            I => \N__45538\
        );

    \I__11066\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45535\
        );

    \I__11065\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45532\
        );

    \I__11064\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45529\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__45535\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__45532\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__45529\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__11060\ : InMux
    port map (
            O => \N__45522\,
            I => \N__45519\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__45519\,
            I => n10957
        );

    \I__11058\ : InMux
    port map (
            O => \N__45516\,
            I => \c0.tx.n16119\
        );

    \I__11057\ : CascadeMux
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__11056\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45506\
        );

    \I__11055\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45503\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__45506\,
            I => \N__45500\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__45503\,
            I => \c0.n10179\
        );

    \I__11052\ : Odrv12
    port map (
            O => \N__45500\,
            I => \c0.n10179\
        );

    \I__11051\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45491\
        );

    \I__11050\ : InMux
    port map (
            O => \N__45494\,
            I => \N__45488\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__45491\,
            I => \N__45485\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__45488\,
            I => \N__45482\
        );

    \I__11047\ : Span4Mux_h
    port map (
            O => \N__45485\,
            I => \N__45479\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__45482\,
            I => \N__45476\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__45479\,
            I => \N__45473\
        );

    \I__11044\ : Odrv4
    port map (
            O => \N__45476\,
            I => \c0.n10188\
        );

    \I__11043\ : Odrv4
    port map (
            O => \N__45473\,
            I => \c0.n10188\
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__45468\,
            I => \c0.n17209_cascade_\
        );

    \I__11041\ : InMux
    port map (
            O => \N__45465\,
            I => \N__45460\
        );

    \I__11040\ : CascadeMux
    port map (
            O => \N__45464\,
            I => \N__45457\
        );

    \I__11039\ : InMux
    port map (
            O => \N__45463\,
            I => \N__45454\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__45460\,
            I => \N__45451\
        );

    \I__11037\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45448\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__45454\,
            I => \c0.data_out_10_2\
        );

    \I__11035\ : Odrv12
    port map (
            O => \N__45451\,
            I => \c0.data_out_10_2\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__45448\,
            I => \c0.data_out_10_2\
        );

    \I__11033\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45438\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__45438\,
            I => \c0.n6_adj_2216\
        );

    \I__11031\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45430\
        );

    \I__11030\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45425\
        );

    \I__11029\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45425\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__45430\,
            I => \c0.data_out_9_6\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__45425\,
            I => \c0.data_out_9_6\
        );

    \I__11026\ : InMux
    port map (
            O => \N__45420\,
            I => \N__45417\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__45417\,
            I => \c0.n17200\
        );

    \I__11024\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45410\
        );

    \I__11023\ : InMux
    port map (
            O => \N__45413\,
            I => \N__45407\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__45410\,
            I => \N__45402\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__45407\,
            I => \N__45399\
        );

    \I__11020\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45393\
        );

    \I__11019\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45393\
        );

    \I__11018\ : Span4Mux_h
    port map (
            O => \N__45402\,
            I => \N__45388\
        );

    \I__11017\ : Span4Mux_v
    port map (
            O => \N__45399\,
            I => \N__45388\
        );

    \I__11016\ : InMux
    port map (
            O => \N__45398\,
            I => \N__45385\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__45393\,
            I => \c0.data_out_8_0\
        );

    \I__11014\ : Odrv4
    port map (
            O => \N__45388\,
            I => \c0.data_out_8_0\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__45385\,
            I => \c0.data_out_8_0\
        );

    \I__11012\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45375\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__45375\,
            I => n8_adj_2445
        );

    \I__11010\ : InMux
    port map (
            O => \N__45372\,
            I => \N__45369\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__45369\,
            I => n6_adj_2446
        );

    \I__11008\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45363\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__45363\,
            I => \N__45360\
        );

    \I__11006\ : Span4Mux_h
    port map (
            O => \N__45360\,
            I => \N__45357\
        );

    \I__11005\ : Odrv4
    port map (
            O => \N__45357\,
            I => n23
        );

    \I__11004\ : InMux
    port map (
            O => \N__45354\,
            I => \N__45351\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__45351\,
            I => \N__45348\
        );

    \I__11002\ : Span4Mux_s1_v
    port map (
            O => \N__45348\,
            I => \N__45345\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__45345\,
            I => \N__45342\
        );

    \I__11000\ : Odrv4
    port map (
            O => \N__45342\,
            I => \c0.n17622\
        );

    \I__10999\ : InMux
    port map (
            O => \N__45339\,
            I => \N__45336\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__45336\,
            I => \c0.n18088\
        );

    \I__10997\ : CascadeMux
    port map (
            O => \N__45333\,
            I => \c0.n2_adj_2164_cascade_\
        );

    \I__10996\ : InMux
    port map (
            O => \N__45330\,
            I => \N__45327\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__45327\,
            I => n18091
        );

    \I__10994\ : InMux
    port map (
            O => \N__45324\,
            I => \N__45318\
        );

    \I__10993\ : InMux
    port map (
            O => \N__45323\,
            I => \N__45318\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__45318\,
            I => data_out_3_5
        );

    \I__10991\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45312\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__45312\,
            I => \N__45309\
        );

    \I__10989\ : Sp12to4
    port map (
            O => \N__45309\,
            I => \N__45305\
        );

    \I__10988\ : InMux
    port map (
            O => \N__45308\,
            I => \N__45302\
        );

    \I__10987\ : Span12Mux_v
    port map (
            O => \N__45305\,
            I => \N__45299\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__45302\,
            I => \c0.data_out_0_6\
        );

    \I__10985\ : Odrv12
    port map (
            O => \N__45299\,
            I => \c0.data_out_0_6\
        );

    \I__10984\ : CascadeMux
    port map (
            O => \N__45294\,
            I => \N__45290\
        );

    \I__10983\ : InMux
    port map (
            O => \N__45293\,
            I => \N__45287\
        );

    \I__10982\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45284\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__45287\,
            I => \N__45281\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__45284\,
            I => \N__45278\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__45281\,
            I => \N__45275\
        );

    \I__10978\ : Span4Mux_v
    port map (
            O => \N__45278\,
            I => \N__45272\
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__45275\,
            I => n4
        );

    \I__10976\ : Odrv4
    port map (
            O => \N__45272\,
            I => n4
        );

    \I__10975\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45264\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__45264\,
            I => \N__45255\
        );

    \I__10973\ : InMux
    port map (
            O => \N__45263\,
            I => \N__45252\
        );

    \I__10972\ : InMux
    port map (
            O => \N__45262\,
            I => \N__45247\
        );

    \I__10971\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45247\
        );

    \I__10970\ : InMux
    port map (
            O => \N__45260\,
            I => \N__45244\
        );

    \I__10969\ : InMux
    port map (
            O => \N__45259\,
            I => \N__45241\
        );

    \I__10968\ : InMux
    port map (
            O => \N__45258\,
            I => \N__45238\
        );

    \I__10967\ : Span4Mux_s1_v
    port map (
            O => \N__45255\,
            I => \N__45235\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__45252\,
            I => \N__45230\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45230\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__45227\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__45241\,
            I => \N__45224\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__45238\,
            I => \N__45221\
        );

    \I__10961\ : Sp12to4
    port map (
            O => \N__45235\,
            I => \N__45211\
        );

    \I__10960\ : Span12Mux_s2_v
    port map (
            O => \N__45230\,
            I => \N__45211\
        );

    \I__10959\ : Span4Mux_h
    port map (
            O => \N__45227\,
            I => \N__45208\
        );

    \I__10958\ : Span4Mux_v
    port map (
            O => \N__45224\,
            I => \N__45203\
        );

    \I__10957\ : Span4Mux_v
    port map (
            O => \N__45221\,
            I => \N__45203\
        );

    \I__10956\ : InMux
    port map (
            O => \N__45220\,
            I => \N__45200\
        );

    \I__10955\ : InMux
    port map (
            O => \N__45219\,
            I => \N__45191\
        );

    \I__10954\ : InMux
    port map (
            O => \N__45218\,
            I => \N__45191\
        );

    \I__10953\ : InMux
    port map (
            O => \N__45217\,
            I => \N__45191\
        );

    \I__10952\ : InMux
    port map (
            O => \N__45216\,
            I => \N__45191\
        );

    \I__10951\ : Span12Mux_v
    port map (
            O => \N__45211\,
            I => \N__45188\
        );

    \I__10950\ : Odrv4
    port map (
            O => \N__45208\,
            I => \r_Rx_Data\
        );

    \I__10949\ : Odrv4
    port map (
            O => \N__45203\,
            I => \r_Rx_Data\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__45200\,
            I => \r_Rx_Data\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__45191\,
            I => \r_Rx_Data\
        );

    \I__10946\ : Odrv12
    port map (
            O => \N__45188\,
            I => \r_Rx_Data\
        );

    \I__10945\ : InMux
    port map (
            O => \N__45177\,
            I => \N__45172\
        );

    \I__10944\ : InMux
    port map (
            O => \N__45176\,
            I => \N__45169\
        );

    \I__10943\ : InMux
    port map (
            O => \N__45175\,
            I => \N__45166\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__45172\,
            I => \N__45163\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__45169\,
            I => \N__45160\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__45166\,
            I => \N__45157\
        );

    \I__10939\ : Span4Mux_v
    port map (
            O => \N__45163\,
            I => \N__45153\
        );

    \I__10938\ : Span4Mux_h
    port map (
            O => \N__45160\,
            I => \N__45150\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__45157\,
            I => \N__45147\
        );

    \I__10936\ : InMux
    port map (
            O => \N__45156\,
            I => \N__45144\
        );

    \I__10935\ : Odrv4
    port map (
            O => \N__45153\,
            I => n9999
        );

    \I__10934\ : Odrv4
    port map (
            O => \N__45150\,
            I => n9999
        );

    \I__10933\ : Odrv4
    port map (
            O => \N__45147\,
            I => n9999
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__45144\,
            I => n9999
        );

    \I__10931\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45127\
        );

    \I__10930\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45124\
        );

    \I__10929\ : CascadeMux
    port map (
            O => \N__45133\,
            I => \N__45121\
        );

    \I__10928\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45113\
        );

    \I__10927\ : InMux
    port map (
            O => \N__45131\,
            I => \N__45113\
        );

    \I__10926\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45113\
        );

    \I__10925\ : LocalMux
    port map (
            O => \N__45127\,
            I => \N__45110\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__45124\,
            I => \N__45107\
        );

    \I__10923\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45104\
        );

    \I__10922\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45101\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45098\
        );

    \I__10920\ : Span4Mux_h
    port map (
            O => \N__45110\,
            I => \N__45094\
        );

    \I__10919\ : Span4Mux_v
    port map (
            O => \N__45107\,
            I => \N__45089\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__45104\,
            I => \N__45089\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__45101\,
            I => \N__45086\
        );

    \I__10916\ : Span4Mux_h
    port map (
            O => \N__45098\,
            I => \N__45083\
        );

    \I__10915\ : CascadeMux
    port map (
            O => \N__45097\,
            I => \N__45080\
        );

    \I__10914\ : Span4Mux_h
    port map (
            O => \N__45094\,
            I => \N__45077\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__45089\,
            I => \N__45074\
        );

    \I__10912\ : Span12Mux_h
    port map (
            O => \N__45086\,
            I => \N__45071\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__45083\,
            I => \N__45068\
        );

    \I__10910\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45065\
        );

    \I__10909\ : Odrv4
    port map (
            O => \N__45077\,
            I => rx_data_4
        );

    \I__10908\ : Odrv4
    port map (
            O => \N__45074\,
            I => rx_data_4
        );

    \I__10907\ : Odrv12
    port map (
            O => \N__45071\,
            I => rx_data_4
        );

    \I__10906\ : Odrv4
    port map (
            O => \N__45068\,
            I => rx_data_4
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__45065\,
            I => rx_data_4
        );

    \I__10904\ : InMux
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__45051\,
            I => \N__45047\
        );

    \I__10902\ : InMux
    port map (
            O => \N__45050\,
            I => \N__45044\
        );

    \I__10901\ : Span4Mux_h
    port map (
            O => \N__45047\,
            I => \N__45041\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__45044\,
            I => data_out_1_6
        );

    \I__10899\ : Odrv4
    port map (
            O => \N__45041\,
            I => data_out_1_6
        );

    \I__10898\ : InMux
    port map (
            O => \N__45036\,
            I => \N__45033\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__45033\,
            I => \N__45025\
        );

    \I__10896\ : InMux
    port map (
            O => \N__45032\,
            I => \N__45022\
        );

    \I__10895\ : InMux
    port map (
            O => \N__45031\,
            I => \N__45014\
        );

    \I__10894\ : InMux
    port map (
            O => \N__45030\,
            I => \N__45011\
        );

    \I__10893\ : InMux
    port map (
            O => \N__45029\,
            I => \N__45008\
        );

    \I__10892\ : InMux
    port map (
            O => \N__45028\,
            I => \N__45005\
        );

    \I__10891\ : Span4Mux_s2_v
    port map (
            O => \N__45025\,
            I => \N__45002\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__45022\,
            I => \N__44999\
        );

    \I__10889\ : InMux
    port map (
            O => \N__45021\,
            I => \N__44996\
        );

    \I__10888\ : InMux
    port map (
            O => \N__45020\,
            I => \N__44993\
        );

    \I__10887\ : InMux
    port map (
            O => \N__45019\,
            I => \N__44987\
        );

    \I__10886\ : InMux
    port map (
            O => \N__45018\,
            I => \N__44983\
        );

    \I__10885\ : CascadeMux
    port map (
            O => \N__45017\,
            I => \N__44979\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__45014\,
            I => \N__44972\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__45011\,
            I => \N__44967\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__45008\,
            I => \N__44967\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__45005\,
            I => \N__44964\
        );

    \I__10880\ : Span4Mux_h
    port map (
            O => \N__45002\,
            I => \N__44955\
        );

    \I__10879\ : Span4Mux_s2_v
    port map (
            O => \N__44999\,
            I => \N__44955\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__44996\,
            I => \N__44955\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__44993\,
            I => \N__44955\
        );

    \I__10876\ : InMux
    port map (
            O => \N__44992\,
            I => \N__44952\
        );

    \I__10875\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44949\
        );

    \I__10874\ : InMux
    port map (
            O => \N__44990\,
            I => \N__44946\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__44987\,
            I => \N__44942\
        );

    \I__10872\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44939\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__44983\,
            I => \N__44936\
        );

    \I__10870\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44933\
        );

    \I__10869\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44928\
        );

    \I__10868\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44925\
        );

    \I__10867\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44922\
        );

    \I__10866\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44919\
        );

    \I__10865\ : InMux
    port map (
            O => \N__44975\,
            I => \N__44916\
        );

    \I__10864\ : Span4Mux_v
    port map (
            O => \N__44972\,
            I => \N__44912\
        );

    \I__10863\ : Span4Mux_v
    port map (
            O => \N__44967\,
            I => \N__44907\
        );

    \I__10862\ : Span4Mux_v
    port map (
            O => \N__44964\,
            I => \N__44907\
        );

    \I__10861\ : Span4Mux_v
    port map (
            O => \N__44955\,
            I => \N__44898\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__44952\,
            I => \N__44898\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44898\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__44946\,
            I => \N__44898\
        );

    \I__10857\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44895\
        );

    \I__10856\ : Span4Mux_v
    port map (
            O => \N__44942\,
            I => \N__44892\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__44939\,
            I => \N__44889\
        );

    \I__10854\ : Span4Mux_h
    port map (
            O => \N__44936\,
            I => \N__44884\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__44933\,
            I => \N__44884\
        );

    \I__10852\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44881\
        );

    \I__10851\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44878\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__44928\,
            I => \N__44871\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__44925\,
            I => \N__44871\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__44922\,
            I => \N__44871\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__44919\,
            I => \N__44866\
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__44916\,
            I => \N__44866\
        );

    \I__10845\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44863\
        );

    \I__10844\ : Span4Mux_h
    port map (
            O => \N__44912\,
            I => \N__44859\
        );

    \I__10843\ : Span4Mux_h
    port map (
            O => \N__44907\,
            I => \N__44854\
        );

    \I__10842\ : Span4Mux_v
    port map (
            O => \N__44898\,
            I => \N__44854\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44851\
        );

    \I__10840\ : Span4Mux_h
    port map (
            O => \N__44892\,
            I => \N__44840\
        );

    \I__10839\ : Span4Mux_v
    port map (
            O => \N__44889\,
            I => \N__44840\
        );

    \I__10838\ : Span4Mux_h
    port map (
            O => \N__44884\,
            I => \N__44840\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__44881\,
            I => \N__44840\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__44878\,
            I => \N__44840\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__44871\,
            I => \N__44833\
        );

    \I__10834\ : Span4Mux_h
    port map (
            O => \N__44866\,
            I => \N__44833\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__44863\,
            I => \N__44833\
        );

    \I__10832\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44830\
        );

    \I__10831\ : Odrv4
    port map (
            O => \N__44859\,
            I => \c0.n9369\
        );

    \I__10830\ : Odrv4
    port map (
            O => \N__44854\,
            I => \c0.n9369\
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__44851\,
            I => \c0.n9369\
        );

    \I__10828\ : Odrv4
    port map (
            O => \N__44840\,
            I => \c0.n9369\
        );

    \I__10827\ : Odrv4
    port map (
            O => \N__44833\,
            I => \c0.n9369\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__44830\,
            I => \c0.n9369\
        );

    \I__10825\ : InMux
    port map (
            O => \N__44817\,
            I => \N__44814\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__44814\,
            I => \N__44808\
        );

    \I__10823\ : InMux
    port map (
            O => \N__44813\,
            I => \N__44805\
        );

    \I__10822\ : InMux
    port map (
            O => \N__44812\,
            I => \N__44802\
        );

    \I__10821\ : InMux
    port map (
            O => \N__44811\,
            I => \N__44795\
        );

    \I__10820\ : Span4Mux_v
    port map (
            O => \N__44808\,
            I => \N__44792\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__44805\,
            I => \N__44787\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__44802\,
            I => \N__44787\
        );

    \I__10817\ : InMux
    port map (
            O => \N__44801\,
            I => \N__44784\
        );

    \I__10816\ : InMux
    port map (
            O => \N__44800\,
            I => \N__44781\
        );

    \I__10815\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44778\
        );

    \I__10814\ : InMux
    port map (
            O => \N__44798\,
            I => \N__44773\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__44795\,
            I => \N__44769\
        );

    \I__10812\ : Span4Mux_h
    port map (
            O => \N__44792\,
            I => \N__44757\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__44787\,
            I => \N__44757\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__44784\,
            I => \N__44757\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__44781\,
            I => \N__44757\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__44778\,
            I => \N__44757\
        );

    \I__10807\ : InMux
    port map (
            O => \N__44777\,
            I => \N__44754\
        );

    \I__10806\ : InMux
    port map (
            O => \N__44776\,
            I => \N__44751\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__44773\,
            I => \N__44748\
        );

    \I__10804\ : InMux
    port map (
            O => \N__44772\,
            I => \N__44745\
        );

    \I__10803\ : Span4Mux_v
    port map (
            O => \N__44769\,
            I => \N__44742\
        );

    \I__10802\ : InMux
    port map (
            O => \N__44768\,
            I => \N__44739\
        );

    \I__10801\ : Span4Mux_v
    port map (
            O => \N__44757\,
            I => \N__44730\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__44754\,
            I => \N__44730\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__44751\,
            I => \N__44730\
        );

    \I__10798\ : Span4Mux_h
    port map (
            O => \N__44748\,
            I => \N__44725\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__44745\,
            I => \N__44725\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__44742\,
            I => \N__44719\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__44739\,
            I => \N__44719\
        );

    \I__10794\ : InMux
    port map (
            O => \N__44738\,
            I => \N__44715\
        );

    \I__10793\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44711\
        );

    \I__10792\ : Span4Mux_h
    port map (
            O => \N__44730\,
            I => \N__44706\
        );

    \I__10791\ : Span4Mux_v
    port map (
            O => \N__44725\,
            I => \N__44706\
        );

    \I__10790\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44703\
        );

    \I__10789\ : Span4Mux_v
    port map (
            O => \N__44719\,
            I => \N__44699\
        );

    \I__10788\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44696\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__44715\,
            I => \N__44693\
        );

    \I__10786\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44690\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__44711\,
            I => \N__44687\
        );

    \I__10784\ : Span4Mux_h
    port map (
            O => \N__44706\,
            I => \N__44682\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__44703\,
            I => \N__44682\
        );

    \I__10782\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44679\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__44699\,
            I => \N__44668\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__44696\,
            I => \N__44668\
        );

    \I__10779\ : Span4Mux_h
    port map (
            O => \N__44693\,
            I => \N__44663\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__44690\,
            I => \N__44663\
        );

    \I__10777\ : Span4Mux_v
    port map (
            O => \N__44687\,
            I => \N__44656\
        );

    \I__10776\ : Span4Mux_h
    port map (
            O => \N__44682\,
            I => \N__44656\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__44679\,
            I => \N__44656\
        );

    \I__10774\ : InMux
    port map (
            O => \N__44678\,
            I => \N__44653\
        );

    \I__10773\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44650\
        );

    \I__10772\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44647\
        );

    \I__10771\ : InMux
    port map (
            O => \N__44675\,
            I => \N__44644\
        );

    \I__10770\ : InMux
    port map (
            O => \N__44674\,
            I => \N__44641\
        );

    \I__10769\ : InMux
    port map (
            O => \N__44673\,
            I => \N__44638\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__44668\,
            I => \c0.n276\
        );

    \I__10767\ : Odrv4
    port map (
            O => \N__44663\,
            I => \c0.n276\
        );

    \I__10766\ : Odrv4
    port map (
            O => \N__44656\,
            I => \c0.n276\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__44653\,
            I => \c0.n276\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__44650\,
            I => \c0.n276\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__44647\,
            I => \c0.n276\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__44644\,
            I => \c0.n276\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__44641\,
            I => \c0.n276\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__44638\,
            I => \c0.n276\
        );

    \I__10759\ : CascadeMux
    port map (
            O => \N__44619\,
            I => \N__44612\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__44618\,
            I => \N__44607\
        );

    \I__10757\ : InMux
    port map (
            O => \N__44617\,
            I => \N__44596\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__44616\,
            I => \N__44593\
        );

    \I__10755\ : InMux
    port map (
            O => \N__44615\,
            I => \N__44590\
        );

    \I__10754\ : InMux
    port map (
            O => \N__44612\,
            I => \N__44587\
        );

    \I__10753\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44584\
        );

    \I__10752\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44580\
        );

    \I__10751\ : InMux
    port map (
            O => \N__44607\,
            I => \N__44577\
        );

    \I__10750\ : InMux
    port map (
            O => \N__44606\,
            I => \N__44574\
        );

    \I__10749\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44570\
        );

    \I__10748\ : CascadeMux
    port map (
            O => \N__44604\,
            I => \N__44567\
        );

    \I__10747\ : CascadeMux
    port map (
            O => \N__44603\,
            I => \N__44561\
        );

    \I__10746\ : InMux
    port map (
            O => \N__44602\,
            I => \N__44558\
        );

    \I__10745\ : InMux
    port map (
            O => \N__44601\,
            I => \N__44555\
        );

    \I__10744\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44552\
        );

    \I__10743\ : InMux
    port map (
            O => \N__44599\,
            I => \N__44549\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__44596\,
            I => \N__44546\
        );

    \I__10741\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44543\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__44590\,
            I => \N__44539\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__44587\,
            I => \N__44536\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__44584\,
            I => \N__44533\
        );

    \I__10737\ : InMux
    port map (
            O => \N__44583\,
            I => \N__44530\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__44580\,
            I => \N__44523\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__44577\,
            I => \N__44523\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__44574\,
            I => \N__44523\
        );

    \I__10733\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44520\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__44570\,
            I => \N__44517\
        );

    \I__10731\ : InMux
    port map (
            O => \N__44567\,
            I => \N__44514\
        );

    \I__10730\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44507\
        );

    \I__10729\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44504\
        );

    \I__10728\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44501\
        );

    \I__10727\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44498\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__44558\,
            I => \N__44493\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__44555\,
            I => \N__44493\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__44552\,
            I => \N__44486\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__44549\,
            I => \N__44486\
        );

    \I__10722\ : Span4Mux_h
    port map (
            O => \N__44546\,
            I => \N__44486\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__44543\,
            I => \N__44483\
        );

    \I__10720\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44480\
        );

    \I__10719\ : Span4Mux_h
    port map (
            O => \N__44539\,
            I => \N__44473\
        );

    \I__10718\ : Span4Mux_s3_v
    port map (
            O => \N__44536\,
            I => \N__44473\
        );

    \I__10717\ : Span4Mux_s3_v
    port map (
            O => \N__44533\,
            I => \N__44473\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__44530\,
            I => \N__44470\
        );

    \I__10715\ : Span4Mux_v
    port map (
            O => \N__44523\,
            I => \N__44467\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__44520\,
            I => \N__44460\
        );

    \I__10713\ : Span4Mux_h
    port map (
            O => \N__44517\,
            I => \N__44460\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__44514\,
            I => \N__44460\
        );

    \I__10711\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44457\
        );

    \I__10710\ : InMux
    port map (
            O => \N__44512\,
            I => \N__44454\
        );

    \I__10709\ : InMux
    port map (
            O => \N__44511\,
            I => \N__44451\
        );

    \I__10708\ : InMux
    port map (
            O => \N__44510\,
            I => \N__44448\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__44507\,
            I => \N__44445\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__44504\,
            I => \N__44442\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__44501\,
            I => \N__44437\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__44498\,
            I => \N__44437\
        );

    \I__10703\ : Span4Mux_h
    port map (
            O => \N__44493\,
            I => \N__44430\
        );

    \I__10702\ : Span4Mux_h
    port map (
            O => \N__44486\,
            I => \N__44430\
        );

    \I__10701\ : Span4Mux_h
    port map (
            O => \N__44483\,
            I => \N__44430\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__44480\,
            I => \N__44425\
        );

    \I__10699\ : Sp12to4
    port map (
            O => \N__44473\,
            I => \N__44425\
        );

    \I__10698\ : Span4Mux_h
    port map (
            O => \N__44470\,
            I => \N__44415\
        );

    \I__10697\ : Span4Mux_h
    port map (
            O => \N__44467\,
            I => \N__44415\
        );

    \I__10696\ : Span4Mux_v
    port map (
            O => \N__44460\,
            I => \N__44415\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__44457\,
            I => \N__44415\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__44454\,
            I => \N__44407\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__44451\,
            I => \N__44407\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__44448\,
            I => \N__44407\
        );

    \I__10691\ : Span4Mux_h
    port map (
            O => \N__44445\,
            I => \N__44400\
        );

    \I__10690\ : Span4Mux_h
    port map (
            O => \N__44442\,
            I => \N__44400\
        );

    \I__10689\ : Span4Mux_h
    port map (
            O => \N__44437\,
            I => \N__44400\
        );

    \I__10688\ : Sp12to4
    port map (
            O => \N__44430\,
            I => \N__44395\
        );

    \I__10687\ : Span12Mux_s10_h
    port map (
            O => \N__44425\,
            I => \N__44395\
        );

    \I__10686\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44392\
        );

    \I__10685\ : Span4Mux_h
    port map (
            O => \N__44415\,
            I => \N__44389\
        );

    \I__10684\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44386\
        );

    \I__10683\ : Odrv12
    port map (
            O => \N__44407\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__10682\ : Odrv4
    port map (
            O => \N__44400\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__10681\ : Odrv12
    port map (
            O => \N__44395\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__44392\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__10679\ : Odrv4
    port map (
            O => \N__44389\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__44386\,
            I => \FRAME_MATCHER_i_31__N_1275\
        );

    \I__10677\ : InMux
    port map (
            O => \N__44373\,
            I => \N__44366\
        );

    \I__10676\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44366\
        );

    \I__10675\ : CascadeMux
    port map (
            O => \N__44371\,
            I => \N__44363\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__44366\,
            I => \N__44360\
        );

    \I__10673\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44357\
        );

    \I__10672\ : Span4Mux_v
    port map (
            O => \N__44360\,
            I => \N__44354\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__44357\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__10670\ : Odrv4
    port map (
            O => \N__44354\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__10669\ : SRMux
    port map (
            O => \N__44349\,
            I => \N__44346\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44343\
        );

    \I__10667\ : Span4Mux_v
    port map (
            O => \N__44343\,
            I => \N__44340\
        );

    \I__10666\ : Span4Mux_h
    port map (
            O => \N__44340\,
            I => \N__44337\
        );

    \I__10665\ : Odrv4
    port map (
            O => \N__44337\,
            I => \c0.n16714\
        );

    \I__10664\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44328\
        );

    \I__10663\ : InMux
    port map (
            O => \N__44333\,
            I => \N__44328\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__44328\,
            I => data_out_1_7
        );

    \I__10661\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44322\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44319\
        );

    \I__10659\ : Span4Mux_v
    port map (
            O => \N__44319\,
            I => \N__44316\
        );

    \I__10658\ : Odrv4
    port map (
            O => \N__44316\,
            I => \c0.n8_adj_2352\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__44313\,
            I => \n5142_cascade_\
        );

    \I__10656\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44307\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__44307\,
            I => \N__44304\
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__44304\,
            I => \c0.tx.n6759\
        );

    \I__10653\ : InMux
    port map (
            O => \N__44301\,
            I => \N__44298\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__44298\,
            I => \c0.tx.n13702\
        );

    \I__10651\ : InMux
    port map (
            O => \N__44295\,
            I => \N__44292\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__44292\,
            I => \c0.tx_active_prev\
        );

    \I__10649\ : InMux
    port map (
            O => \N__44289\,
            I => \N__44282\
        );

    \I__10648\ : InMux
    port map (
            O => \N__44288\,
            I => \N__44279\
        );

    \I__10647\ : InMux
    port map (
            O => \N__44287\,
            I => \N__44274\
        );

    \I__10646\ : InMux
    port map (
            O => \N__44286\,
            I => \N__44274\
        );

    \I__10645\ : InMux
    port map (
            O => \N__44285\,
            I => \N__44271\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__44282\,
            I => \N__44268\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__44279\,
            I => \N__44265\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__44274\,
            I => \N__44262\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__44271\,
            I => \N__44259\
        );

    \I__10640\ : Span4Mux_s2_v
    port map (
            O => \N__44268\,
            I => \N__44256\
        );

    \I__10639\ : Span4Mux_h
    port map (
            O => \N__44265\,
            I => \N__44253\
        );

    \I__10638\ : Span4Mux_h
    port map (
            O => \N__44262\,
            I => \N__44250\
        );

    \I__10637\ : Span4Mux_h
    port map (
            O => \N__44259\,
            I => \N__44245\
        );

    \I__10636\ : Span4Mux_h
    port map (
            O => \N__44256\,
            I => \N__44245\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__44253\,
            I => \c0.data_out_5_5\
        );

    \I__10634\ : Odrv4
    port map (
            O => \N__44250\,
            I => \c0.data_out_5_5\
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__44245\,
            I => \c0.data_out_5_5\
        );

    \I__10632\ : InMux
    port map (
            O => \N__44238\,
            I => \N__44235\
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__10630\ : Span12Mux_s2_v
    port map (
            O => \N__44232\,
            I => \N__44229\
        );

    \I__10629\ : Odrv12
    port map (
            O => \N__44229\,
            I => \c0.n5_adj_2163\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__44226\,
            I => \c0.n17581_cascade_\
        );

    \I__10627\ : CascadeMux
    port map (
            O => \N__44223\,
            I => \N__44220\
        );

    \I__10626\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44217\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__44217\,
            I => n10_adj_2432
        );

    \I__10624\ : InMux
    port map (
            O => \N__44214\,
            I => \N__44209\
        );

    \I__10623\ : CascadeMux
    port map (
            O => \N__44213\,
            I => \N__44205\
        );

    \I__10622\ : CascadeMux
    port map (
            O => \N__44212\,
            I => \N__44200\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__44209\,
            I => \N__44197\
        );

    \I__10620\ : InMux
    port map (
            O => \N__44208\,
            I => \N__44194\
        );

    \I__10619\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44188\
        );

    \I__10618\ : InMux
    port map (
            O => \N__44204\,
            I => \N__44181\
        );

    \I__10617\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44181\
        );

    \I__10616\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44181\
        );

    \I__10615\ : Span4Mux_v
    port map (
            O => \N__44197\,
            I => \N__44173\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__44194\,
            I => \N__44173\
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__44193\,
            I => \N__44170\
        );

    \I__10612\ : CascadeMux
    port map (
            O => \N__44192\,
            I => \N__44167\
        );

    \I__10611\ : CascadeMux
    port map (
            O => \N__44191\,
            I => \N__44164\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__44188\,
            I => \N__44161\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__44181\,
            I => \N__44158\
        );

    \I__10608\ : InMux
    port map (
            O => \N__44180\,
            I => \N__44155\
        );

    \I__10607\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44152\
        );

    \I__10606\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44149\
        );

    \I__10605\ : Span4Mux_h
    port map (
            O => \N__44173\,
            I => \N__44146\
        );

    \I__10604\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44139\
        );

    \I__10603\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44139\
        );

    \I__10602\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44139\
        );

    \I__10601\ : Span4Mux_h
    port map (
            O => \N__44161\,
            I => \N__44134\
        );

    \I__10600\ : Span4Mux_v
    port map (
            O => \N__44158\,
            I => \N__44134\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__44155\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__44152\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__44149\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__10596\ : Odrv4
    port map (
            O => \N__44146\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__44139\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__10594\ : Odrv4
    port map (
            O => \N__44134\,
            I => \c0.tx.r_SM_Main_1\
        );

    \I__10593\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44118\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__44118\,
            I => \c0.tx.n10613\
        );

    \I__10591\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44112\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__44112\,
            I => \c0.tx.n12_adj_2134\
        );

    \I__10589\ : CascadeMux
    port map (
            O => \N__44109\,
            I => \c0.n8_cascade_\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__44106\,
            I => \N__44100\
        );

    \I__10587\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44094\
        );

    \I__10586\ : InMux
    port map (
            O => \N__44104\,
            I => \N__44091\
        );

    \I__10585\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44088\
        );

    \I__10584\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44085\
        );

    \I__10583\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44082\
        );

    \I__10582\ : CascadeMux
    port map (
            O => \N__44098\,
            I => \N__44079\
        );

    \I__10581\ : CascadeMux
    port map (
            O => \N__44097\,
            I => \N__44076\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__44094\,
            I => \N__44072\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44069\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__44088\,
            I => \N__44066\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__44085\,
            I => \N__44063\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44060\
        );

    \I__10575\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44055\
        );

    \I__10574\ : InMux
    port map (
            O => \N__44076\,
            I => \N__44055\
        );

    \I__10573\ : CascadeMux
    port map (
            O => \N__44075\,
            I => \N__44052\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__44072\,
            I => \N__44049\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__44069\,
            I => \N__44044\
        );

    \I__10570\ : Span4Mux_h
    port map (
            O => \N__44066\,
            I => \N__44044\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__44063\,
            I => \N__44039\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__44060\,
            I => \N__44039\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__44055\,
            I => \N__44036\
        );

    \I__10566\ : InMux
    port map (
            O => \N__44052\,
            I => \N__44033\
        );

    \I__10565\ : Odrv4
    port map (
            O => \N__44049\,
            I => n9257
        );

    \I__10564\ : Odrv4
    port map (
            O => \N__44044\,
            I => n9257
        );

    \I__10563\ : Odrv4
    port map (
            O => \N__44039\,
            I => n9257
        );

    \I__10562\ : Odrv12
    port map (
            O => \N__44036\,
            I => n9257
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__44033\,
            I => n9257
        );

    \I__10560\ : InMux
    port map (
            O => \N__44022\,
            I => \N__44019\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__44019\,
            I => \c0.n65_adj_2192\
        );

    \I__10558\ : InMux
    port map (
            O => \N__44016\,
            I => \N__44011\
        );

    \I__10557\ : InMux
    port map (
            O => \N__44015\,
            I => \N__44008\
        );

    \I__10556\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44005\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__44011\,
            I => \N__44000\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__44008\,
            I => \N__43993\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__44005\,
            I => \N__43993\
        );

    \I__10552\ : CascadeMux
    port map (
            O => \N__44004\,
            I => \N__43990\
        );

    \I__10551\ : CascadeMux
    port map (
            O => \N__44003\,
            I => \N__43987\
        );

    \I__10550\ : Span4Mux_h
    port map (
            O => \N__44000\,
            I => \N__43982\
        );

    \I__10549\ : InMux
    port map (
            O => \N__43999\,
            I => \N__43977\
        );

    \I__10548\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43977\
        );

    \I__10547\ : Span4Mux_h
    port map (
            O => \N__43993\,
            I => \N__43974\
        );

    \I__10546\ : InMux
    port map (
            O => \N__43990\,
            I => \N__43965\
        );

    \I__10545\ : InMux
    port map (
            O => \N__43987\,
            I => \N__43965\
        );

    \I__10544\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43965\
        );

    \I__10543\ : InMux
    port map (
            O => \N__43985\,
            I => \N__43965\
        );

    \I__10542\ : Odrv4
    port map (
            O => \N__43982\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__43977\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__10540\ : Odrv4
    port map (
            O => \N__43974\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__43965\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__10538\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43953\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__43953\,
            I => \N__43947\
        );

    \I__10536\ : InMux
    port map (
            O => \N__43952\,
            I => \N__43942\
        );

    \I__10535\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43942\
        );

    \I__10534\ : InMux
    port map (
            O => \N__43950\,
            I => \N__43939\
        );

    \I__10533\ : Span4Mux_v
    port map (
            O => \N__43947\,
            I => \N__43933\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__43942\,
            I => \N__43930\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__43939\,
            I => \N__43927\
        );

    \I__10530\ : InMux
    port map (
            O => \N__43938\,
            I => \N__43924\
        );

    \I__10529\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43919\
        );

    \I__10528\ : InMux
    port map (
            O => \N__43936\,
            I => \N__43919\
        );

    \I__10527\ : Odrv4
    port map (
            O => \N__43933\,
            I => \c0.tx.n83\
        );

    \I__10526\ : Odrv12
    port map (
            O => \N__43930\,
            I => \c0.tx.n83\
        );

    \I__10525\ : Odrv12
    port map (
            O => \N__43927\,
            I => \c0.tx.n83\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__43924\,
            I => \c0.tx.n83\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__43919\,
            I => \c0.tx.n83\
        );

    \I__10522\ : InMux
    port map (
            O => \N__43908\,
            I => \N__43905\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__43905\,
            I => \N__43902\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__43902\,
            I => n10_adj_2422
        );

    \I__10519\ : CascadeMux
    port map (
            O => \N__43899\,
            I => \c0.tx.n77_cascade_\
        );

    \I__10518\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43893\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__43893\,
            I => \N__43890\
        );

    \I__10516\ : Odrv4
    port map (
            O => \N__43890\,
            I => \c0.tx.n12\
        );

    \I__10515\ : IoInMux
    port map (
            O => \N__43887\,
            I => \N__43884\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__43884\,
            I => \N__43881\
        );

    \I__10513\ : IoSpan4Mux
    port map (
            O => \N__43881\,
            I => \N__43877\
        );

    \I__10512\ : InMux
    port map (
            O => \N__43880\,
            I => \N__43874\
        );

    \I__10511\ : Span4Mux_s3_v
    port map (
            O => \N__43877\,
            I => \N__43871\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__43874\,
            I => \N__43868\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__43871\,
            I => \N__43863\
        );

    \I__10508\ : Span4Mux_h
    port map (
            O => \N__43868\,
            I => \N__43863\
        );

    \I__10507\ : Span4Mux_h
    port map (
            O => \N__43863\,
            I => \N__43859\
        );

    \I__10506\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43856\
        );

    \I__10505\ : Odrv4
    port map (
            O => \N__43859\,
            I => tx_o
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__43856\,
            I => tx_o
        );

    \I__10503\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43848\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__43848\,
            I => \c0.tx.n10\
        );

    \I__10501\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43837\
        );

    \I__10500\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43831\
        );

    \I__10499\ : InMux
    port map (
            O => \N__43843\,
            I => \N__43831\
        );

    \I__10498\ : CascadeMux
    port map (
            O => \N__43842\,
            I => \N__43828\
        );

    \I__10497\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43825\
        );

    \I__10496\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43822\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__43837\,
            I => \N__43819\
        );

    \I__10494\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43816\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43810\
        );

    \I__10492\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43807\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__43825\,
            I => \N__43804\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43801\
        );

    \I__10489\ : Span4Mux_s2_v
    port map (
            O => \N__43819\,
            I => \N__43796\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__43816\,
            I => \N__43796\
        );

    \I__10487\ : InMux
    port map (
            O => \N__43815\,
            I => \N__43793\
        );

    \I__10486\ : InMux
    port map (
            O => \N__43814\,
            I => \N__43788\
        );

    \I__10485\ : InMux
    port map (
            O => \N__43813\,
            I => \N__43788\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__43810\,
            I => \N__43785\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__43807\,
            I => \N__43778\
        );

    \I__10482\ : Span4Mux_v
    port map (
            O => \N__43804\,
            I => \N__43778\
        );

    \I__10481\ : Span4Mux_h
    port map (
            O => \N__43801\,
            I => \N__43778\
        );

    \I__10480\ : Span4Mux_v
    port map (
            O => \N__43796\,
            I => \N__43775\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__43793\,
            I => byte_transmit_counter_4
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__43788\,
            I => byte_transmit_counter_4
        );

    \I__10477\ : Odrv4
    port map (
            O => \N__43785\,
            I => byte_transmit_counter_4
        );

    \I__10476\ : Odrv4
    port map (
            O => \N__43778\,
            I => byte_transmit_counter_4
        );

    \I__10475\ : Odrv4
    port map (
            O => \N__43775\,
            I => byte_transmit_counter_4
        );

    \I__10474\ : InMux
    port map (
            O => \N__43764\,
            I => \N__43761\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__43761\,
            I => n10_adj_2443
        );

    \I__10472\ : InMux
    port map (
            O => \N__43758\,
            I => \N__43754\
        );

    \I__10471\ : InMux
    port map (
            O => \N__43757\,
            I => \N__43751\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__43754\,
            I => \N__43748\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__43751\,
            I => \r_Tx_Data_6\
        );

    \I__10468\ : Odrv4
    port map (
            O => \N__43748\,
            I => \r_Tx_Data_6\
        );

    \I__10467\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43740\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__43740\,
            I => \N__43737\
        );

    \I__10465\ : Span4Mux_v
    port map (
            O => \N__43737\,
            I => \N__43733\
        );

    \I__10464\ : CascadeMux
    port map (
            O => \N__43736\,
            I => \N__43730\
        );

    \I__10463\ : Span4Mux_h
    port map (
            O => \N__43733\,
            I => \N__43727\
        );

    \I__10462\ : InMux
    port map (
            O => \N__43730\,
            I => \N__43724\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__43727\,
            I => rand_setpoint_5
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__43724\,
            I => rand_setpoint_5
        );

    \I__10459\ : CascadeMux
    port map (
            O => \N__43719\,
            I => \N__43712\
        );

    \I__10458\ : CascadeMux
    port map (
            O => \N__43718\,
            I => \N__43709\
        );

    \I__10457\ : InMux
    port map (
            O => \N__43717\,
            I => \N__43706\
        );

    \I__10456\ : CascadeMux
    port map (
            O => \N__43716\,
            I => \N__43703\
        );

    \I__10455\ : CascadeMux
    port map (
            O => \N__43715\,
            I => \N__43700\
        );

    \I__10454\ : InMux
    port map (
            O => \N__43712\,
            I => \N__43697\
        );

    \I__10453\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43694\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__43706\,
            I => \N__43690\
        );

    \I__10451\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43687\
        );

    \I__10450\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43684\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__43697\,
            I => \N__43681\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__43694\,
            I => \N__43678\
        );

    \I__10447\ : InMux
    port map (
            O => \N__43693\,
            I => \N__43675\
        );

    \I__10446\ : Span4Mux_h
    port map (
            O => \N__43690\,
            I => \N__43668\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__43687\,
            I => \N__43668\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__43684\,
            I => \N__43668\
        );

    \I__10443\ : Span4Mux_v
    port map (
            O => \N__43681\,
            I => \N__43665\
        );

    \I__10442\ : Span4Mux_h
    port map (
            O => \N__43678\,
            I => \N__43662\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__43675\,
            I => \N__43657\
        );

    \I__10440\ : Span4Mux_v
    port map (
            O => \N__43668\,
            I => \N__43657\
        );

    \I__10439\ : Odrv4
    port map (
            O => \N__43665\,
            I => n2594
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__43662\,
            I => n2594
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__43657\,
            I => n2594
        );

    \I__10436\ : CascadeMux
    port map (
            O => \N__43650\,
            I => \N__43647\
        );

    \I__10435\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43643\
        );

    \I__10434\ : CascadeMux
    port map (
            O => \N__43646\,
            I => \N__43640\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__43643\,
            I => \N__43637\
        );

    \I__10432\ : InMux
    port map (
            O => \N__43640\,
            I => \N__43634\
        );

    \I__10431\ : Odrv12
    port map (
            O => \N__43637\,
            I => rand_setpoint_13
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__43634\,
            I => rand_setpoint_13
        );

    \I__10429\ : InMux
    port map (
            O => \N__43629\,
            I => \N__43626\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__43626\,
            I => \N__43621\
        );

    \I__10427\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43616\
        );

    \I__10426\ : InMux
    port map (
            O => \N__43624\,
            I => \N__43616\
        );

    \I__10425\ : Span12Mux_s6_v
    port map (
            O => \N__43621\,
            I => \N__43613\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__43616\,
            I => \c0.data_out_7_5\
        );

    \I__10423\ : Odrv12
    port map (
            O => \N__43613\,
            I => \c0.data_out_7_5\
        );

    \I__10422\ : CascadeMux
    port map (
            O => \N__43608\,
            I => \N__43605\
        );

    \I__10421\ : InMux
    port map (
            O => \N__43605\,
            I => \N__43602\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__43602\,
            I => \N__43598\
        );

    \I__10419\ : InMux
    port map (
            O => \N__43601\,
            I => \N__43595\
        );

    \I__10418\ : Span4Mux_h
    port map (
            O => \N__43598\,
            I => \N__43592\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__43595\,
            I => \r_Tx_Data_7\
        );

    \I__10416\ : Odrv4
    port map (
            O => \N__43592\,
            I => \r_Tx_Data_7\
        );

    \I__10415\ : InMux
    port map (
            O => \N__43587\,
            I => \N__43584\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__43584\,
            I => \N__43581\
        );

    \I__10413\ : Span4Mux_h
    port map (
            O => \N__43581\,
            I => \N__43578\
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__43578\,
            I => \c0.data_out_1_1\
        );

    \I__10411\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43571\
        );

    \I__10410\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43568\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__43571\,
            I => data_out_0_1
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__43568\,
            I => data_out_0_1
        );

    \I__10407\ : InMux
    port map (
            O => \N__43563\,
            I => \N__43560\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__43560\,
            I => n1_adj_2449
        );

    \I__10405\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43554\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__43554\,
            I => \c0.n12630\
        );

    \I__10403\ : InMux
    port map (
            O => \N__43551\,
            I => \N__43546\
        );

    \I__10402\ : InMux
    port map (
            O => \N__43550\,
            I => \N__43543\
        );

    \I__10401\ : InMux
    port map (
            O => \N__43549\,
            I => \N__43540\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__43546\,
            I => \c0.data_out_7_0\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__43543\,
            I => \c0.data_out_7_0\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__43540\,
            I => \c0.data_out_7_0\
        );

    \I__10397\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43530\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__43530\,
            I => \N__43526\
        );

    \I__10395\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43523\
        );

    \I__10394\ : Odrv4
    port map (
            O => \N__43526\,
            I => \c0.n10395\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__43523\,
            I => \c0.n10395\
        );

    \I__10392\ : CascadeMux
    port map (
            O => \N__43518\,
            I => \c0.n10_adj_2189_cascade_\
        );

    \I__10391\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43512\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__43512\,
            I => \N__43508\
        );

    \I__10389\ : InMux
    port map (
            O => \N__43511\,
            I => \N__43505\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__43508\,
            I => \N__43502\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__43505\,
            I => \r_Tx_Data_0\
        );

    \I__10386\ : Odrv4
    port map (
            O => \N__43502\,
            I => \r_Tx_Data_0\
        );

    \I__10385\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43494\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__43494\,
            I => \c0.n8_adj_2157\
        );

    \I__10383\ : InMux
    port map (
            O => \N__43491\,
            I => \N__43488\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__43488\,
            I => \c0.n15_adj_2177\
        );

    \I__10381\ : CascadeMux
    port map (
            O => \N__43485\,
            I => \N__43482\
        );

    \I__10380\ : InMux
    port map (
            O => \N__43482\,
            I => \N__43479\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__43479\,
            I => \N__43476\
        );

    \I__10378\ : Span4Mux_v
    port map (
            O => \N__43476\,
            I => \N__43473\
        );

    \I__10377\ : Odrv4
    port map (
            O => \N__43473\,
            I => \c0.n17270\
        );

    \I__10376\ : InMux
    port map (
            O => \N__43470\,
            I => \N__43466\
        );

    \I__10375\ : InMux
    port map (
            O => \N__43469\,
            I => \N__43462\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__43466\,
            I => \N__43459\
        );

    \I__10373\ : InMux
    port map (
            O => \N__43465\,
            I => \N__43456\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__43462\,
            I => \N__43453\
        );

    \I__10371\ : Span4Mux_v
    port map (
            O => \N__43459\,
            I => \N__43450\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__43456\,
            I => \N__43447\
        );

    \I__10369\ : Span12Mux_v
    port map (
            O => \N__43453\,
            I => \N__43444\
        );

    \I__10368\ : Span4Mux_h
    port map (
            O => \N__43450\,
            I => \N__43441\
        );

    \I__10367\ : Span4Mux_h
    port map (
            O => \N__43447\,
            I => \N__43438\
        );

    \I__10366\ : Odrv12
    port map (
            O => \N__43444\,
            I => \c0.data_out_7_2\
        );

    \I__10365\ : Odrv4
    port map (
            O => \N__43441\,
            I => \c0.data_out_7_2\
        );

    \I__10364\ : Odrv4
    port map (
            O => \N__43438\,
            I => \c0.data_out_7_2\
        );

    \I__10363\ : InMux
    port map (
            O => \N__43431\,
            I => \N__43428\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__43428\,
            I => \c0.n10316\
        );

    \I__10361\ : InMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__43422\,
            I => \c0.n17201\
        );

    \I__10359\ : CascadeMux
    port map (
            O => \N__43419\,
            I => \c0.n10316_cascade_\
        );

    \I__10358\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43410\
        );

    \I__10357\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43410\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__43410\,
            I => \c0.n17177\
        );

    \I__10355\ : InMux
    port map (
            O => \N__43407\,
            I => \N__43403\
        );

    \I__10354\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43400\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__43403\,
            I => \N__43395\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__43400\,
            I => \N__43392\
        );

    \I__10351\ : InMux
    port map (
            O => \N__43399\,
            I => \N__43387\
        );

    \I__10350\ : InMux
    port map (
            O => \N__43398\,
            I => \N__43387\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__43395\,
            I => \N__43383\
        );

    \I__10348\ : Span4Mux_v
    port map (
            O => \N__43392\,
            I => \N__43378\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__43387\,
            I => \N__43378\
        );

    \I__10346\ : InMux
    port map (
            O => \N__43386\,
            I => \N__43375\
        );

    \I__10345\ : Span4Mux_v
    port map (
            O => \N__43383\,
            I => \N__43372\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__43378\,
            I => \N__43369\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__43375\,
            I => data_out_8_6
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__43372\,
            I => data_out_8_6
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__43369\,
            I => data_out_8_6
        );

    \I__10340\ : InMux
    port map (
            O => \N__43362\,
            I => \N__43353\
        );

    \I__10339\ : InMux
    port map (
            O => \N__43361\,
            I => \N__43353\
        );

    \I__10338\ : InMux
    port map (
            O => \N__43360\,
            I => \N__43350\
        );

    \I__10337\ : InMux
    port map (
            O => \N__43359\,
            I => \N__43345\
        );

    \I__10336\ : InMux
    port map (
            O => \N__43358\,
            I => \N__43345\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__43353\,
            I => \N__43342\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__43350\,
            I => \N__43337\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__43345\,
            I => \N__43337\
        );

    \I__10332\ : Span4Mux_v
    port map (
            O => \N__43342\,
            I => \N__43334\
        );

    \I__10331\ : Span4Mux_v
    port map (
            O => \N__43337\,
            I => \N__43331\
        );

    \I__10330\ : Sp12to4
    port map (
            O => \N__43334\,
            I => \N__43326\
        );

    \I__10329\ : Sp12to4
    port map (
            O => \N__43331\,
            I => \N__43326\
        );

    \I__10328\ : Span12Mux_h
    port map (
            O => \N__43326\,
            I => \N__43323\
        );

    \I__10327\ : Odrv12
    port map (
            O => \N__43323\,
            I => \c0.data_out_6__1__N_537\
        );

    \I__10326\ : InMux
    port map (
            O => \N__43320\,
            I => \N__43317\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__43317\,
            I => \N__43314\
        );

    \I__10324\ : Span4Mux_v
    port map (
            O => \N__43314\,
            I => \N__43310\
        );

    \I__10323\ : InMux
    port map (
            O => \N__43313\,
            I => \N__43305\
        );

    \I__10322\ : Sp12to4
    port map (
            O => \N__43310\,
            I => \N__43302\
        );

    \I__10321\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43297\
        );

    \I__10320\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43297\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__43305\,
            I => \c0.data_out_7_7\
        );

    \I__10318\ : Odrv12
    port map (
            O => \N__43302\,
            I => \c0.data_out_7_7\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__43297\,
            I => \c0.data_out_7_7\
        );

    \I__10316\ : InMux
    port map (
            O => \N__43290\,
            I => \N__43287\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__43287\,
            I => n10_adj_2483
        );

    \I__10314\ : InMux
    port map (
            O => \N__43284\,
            I => \N__43281\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__43281\,
            I => \N__43277\
        );

    \I__10312\ : InMux
    port map (
            O => \N__43280\,
            I => \N__43274\
        );

    \I__10311\ : Span4Mux_v
    port map (
            O => \N__43277\,
            I => \N__43271\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__43274\,
            I => \c0.data_out_3_6\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__43271\,
            I => \c0.data_out_3_6\
        );

    \I__10308\ : CascadeMux
    port map (
            O => \N__43266\,
            I => \N__43261\
        );

    \I__10307\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43256\
        );

    \I__10306\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43256\
        );

    \I__10305\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43253\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__43256\,
            I => \N__43250\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__43253\,
            I => \N__43245\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__43250\,
            I => \N__43245\
        );

    \I__10301\ : Odrv4
    port map (
            O => \N__43245\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__10300\ : SRMux
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__43239\,
            I => \N__43236\
        );

    \I__10298\ : Span4Mux_v
    port map (
            O => \N__43236\,
            I => \N__43233\
        );

    \I__10297\ : Odrv4
    port map (
            O => \N__43233\,
            I => \c0.n16690\
        );

    \I__10296\ : CascadeMux
    port map (
            O => \N__43230\,
            I => \N__43226\
        );

    \I__10295\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43222\
        );

    \I__10294\ : InMux
    port map (
            O => \N__43226\,
            I => \N__43219\
        );

    \I__10293\ : InMux
    port map (
            O => \N__43225\,
            I => \N__43216\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__43222\,
            I => \N__43211\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__43219\,
            I => \N__43211\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__43216\,
            I => \N__43206\
        );

    \I__10289\ : Span4Mux_v
    port map (
            O => \N__43211\,
            I => \N__43206\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__43206\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__10287\ : SRMux
    port map (
            O => \N__43203\,
            I => \N__43200\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__43200\,
            I => \N__43197\
        );

    \I__10285\ : Span4Mux_h
    port map (
            O => \N__43197\,
            I => \N__43194\
        );

    \I__10284\ : Odrv4
    port map (
            O => \N__43194\,
            I => \c0.n16702\
        );

    \I__10283\ : InMux
    port map (
            O => \N__43191\,
            I => \N__43187\
        );

    \I__10282\ : CascadeMux
    port map (
            O => \N__43190\,
            I => \N__43184\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__43187\,
            I => \N__43180\
        );

    \I__10280\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43177\
        );

    \I__10279\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43174\
        );

    \I__10278\ : Span4Mux_h
    port map (
            O => \N__43180\,
            I => \N__43171\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__43177\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__43174\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__10275\ : Odrv4
    port map (
            O => \N__43171\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__10274\ : SRMux
    port map (
            O => \N__43164\,
            I => \N__43161\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__43161\,
            I => \c0.n8_adj_2330\
        );

    \I__10272\ : InMux
    port map (
            O => \N__43158\,
            I => \N__43154\
        );

    \I__10271\ : CascadeMux
    port map (
            O => \N__43157\,
            I => \N__43151\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__43154\,
            I => \N__43147\
        );

    \I__10269\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43144\
        );

    \I__10268\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43141\
        );

    \I__10267\ : Span4Mux_h
    port map (
            O => \N__43147\,
            I => \N__43138\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__43144\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__43141\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__43138\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__10263\ : SRMux
    port map (
            O => \N__43131\,
            I => \N__43128\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__43128\,
            I => \N__43125\
        );

    \I__10261\ : Span4Mux_v
    port map (
            O => \N__43125\,
            I => \N__43122\
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__43122\,
            I => \c0.n16686\
        );

    \I__10259\ : CascadeMux
    port map (
            O => \N__43119\,
            I => \N__43115\
        );

    \I__10258\ : InMux
    port map (
            O => \N__43118\,
            I => \N__43111\
        );

    \I__10257\ : InMux
    port map (
            O => \N__43115\,
            I => \N__43108\
        );

    \I__10256\ : CascadeMux
    port map (
            O => \N__43114\,
            I => \N__43105\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__43111\,
            I => \N__43100\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__43108\,
            I => \N__43100\
        );

    \I__10253\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43097\
        );

    \I__10252\ : Span4Mux_h
    port map (
            O => \N__43100\,
            I => \N__43094\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__43097\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__10250\ : Odrv4
    port map (
            O => \N__43094\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__10249\ : SRMux
    port map (
            O => \N__43089\,
            I => \N__43086\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__43086\,
            I => \N__43083\
        );

    \I__10247\ : Odrv4
    port map (
            O => \N__43083\,
            I => \c0.n16688\
        );

    \I__10246\ : CascadeMux
    port map (
            O => \N__43080\,
            I => \c0.n68_cascade_\
        );

    \I__10245\ : InMux
    port map (
            O => \N__43077\,
            I => \N__43072\
        );

    \I__10244\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43069\
        );

    \I__10243\ : InMux
    port map (
            O => \N__43075\,
            I => \N__43066\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__43072\,
            I => \tx_transmit_N_1947_7\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__43069\,
            I => \tx_transmit_N_1947_7\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__43066\,
            I => \tx_transmit_N_1947_7\
        );

    \I__10239\ : SRMux
    port map (
            O => \N__43059\,
            I => \N__43056\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__43056\,
            I => \N__43053\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__43053\,
            I => \c0.n4650\
        );

    \I__10236\ : InMux
    port map (
            O => \N__43050\,
            I => \N__43047\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__43047\,
            I => \N__43044\
        );

    \I__10234\ : Span4Mux_h
    port map (
            O => \N__43044\,
            I => \N__43035\
        );

    \I__10233\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43030\
        );

    \I__10232\ : InMux
    port map (
            O => \N__43042\,
            I => \N__43030\
        );

    \I__10231\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43027\
        );

    \I__10230\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43022\
        );

    \I__10229\ : InMux
    port map (
            O => \N__43039\,
            I => \N__43022\
        );

    \I__10228\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43019\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__43035\,
            I => \tx_transmit_N_1947_3\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__43030\,
            I => \tx_transmit_N_1947_3\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__43027\,
            I => \tx_transmit_N_1947_3\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__43022\,
            I => \tx_transmit_N_1947_3\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__43019\,
            I => \tx_transmit_N_1947_3\
        );

    \I__10222\ : InMux
    port map (
            O => \N__43008\,
            I => \N__43005\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__43005\,
            I => \c0.n59\
        );

    \I__10220\ : CascadeMux
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__10219\ : InMux
    port map (
            O => \N__42999\,
            I => \N__42996\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__42996\,
            I => \c0.n65\
        );

    \I__10217\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42990\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__42990\,
            I => \N__42986\
        );

    \I__10215\ : CascadeMux
    port map (
            O => \N__42989\,
            I => \N__42982\
        );

    \I__10214\ : Span4Mux_h
    port map (
            O => \N__42986\,
            I => \N__42979\
        );

    \I__10213\ : InMux
    port map (
            O => \N__42985\,
            I => \N__42976\
        );

    \I__10212\ : InMux
    port map (
            O => \N__42982\,
            I => \N__42973\
        );

    \I__10211\ : Odrv4
    port map (
            O => \N__42979\,
            I => \tx_transmit_N_1947_4\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__42976\,
            I => \tx_transmit_N_1947_4\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__42973\,
            I => \tx_transmit_N_1947_4\
        );

    \I__10208\ : CascadeMux
    port map (
            O => \N__42966\,
            I => \N__42963\
        );

    \I__10207\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42958\
        );

    \I__10206\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42955\
        );

    \I__10205\ : InMux
    port map (
            O => \N__42961\,
            I => \N__42952\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__42958\,
            I => \tx_transmit_N_1947_5\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__42955\,
            I => \tx_transmit_N_1947_5\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__42952\,
            I => \tx_transmit_N_1947_5\
        );

    \I__10201\ : InMux
    port map (
            O => \N__42945\,
            I => \N__42942\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__42942\,
            I => \N__42939\
        );

    \I__10199\ : Span4Mux_h
    port map (
            O => \N__42939\,
            I => \N__42936\
        );

    \I__10198\ : Span4Mux_v
    port map (
            O => \N__42936\,
            I => \N__42931\
        );

    \I__10197\ : InMux
    port map (
            O => \N__42935\,
            I => \N__42928\
        );

    \I__10196\ : InMux
    port map (
            O => \N__42934\,
            I => \N__42925\
        );

    \I__10195\ : Odrv4
    port map (
            O => \N__42931\,
            I => \tx_transmit_N_1947_6\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__42928\,
            I => \tx_transmit_N_1947_6\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__42925\,
            I => \tx_transmit_N_1947_6\
        );

    \I__10192\ : InMux
    port map (
            O => \N__42918\,
            I => \N__42915\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__42915\,
            I => \c0.n17404\
        );

    \I__10190\ : InMux
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__42909\,
            I => \N__42906\
        );

    \I__10188\ : Span4Mux_h
    port map (
            O => \N__42906\,
            I => \N__42902\
        );

    \I__10187\ : InMux
    port map (
            O => \N__42905\,
            I => \N__42899\
        );

    \I__10186\ : Odrv4
    port map (
            O => \N__42902\,
            I => \tx_transmit_N_1947_1\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__42899\,
            I => \tx_transmit_N_1947_1\
        );

    \I__10184\ : InMux
    port map (
            O => \N__42894\,
            I => \N__42891\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__42891\,
            I => \N__42888\
        );

    \I__10182\ : Span4Mux_v
    port map (
            O => \N__42888\,
            I => \N__42884\
        );

    \I__10181\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42881\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__42884\,
            I => \tx_transmit_N_1947_0\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__42881\,
            I => \tx_transmit_N_1947_0\
        );

    \I__10178\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42871\
        );

    \I__10177\ : InMux
    port map (
            O => \N__42875\,
            I => \N__42868\
        );

    \I__10176\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42865\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42862\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__42868\,
            I => \c0.n13662\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__42865\,
            I => \c0.n13662\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__42862\,
            I => \c0.n13662\
        );

    \I__10171\ : CascadeMux
    port map (
            O => \N__42855\,
            I => \c0.n13662_cascade_\
        );

    \I__10170\ : InMux
    port map (
            O => \N__42852\,
            I => \N__42849\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__42849\,
            I => \N__42846\
        );

    \I__10168\ : Span4Mux_h
    port map (
            O => \N__42846\,
            I => \N__42838\
        );

    \I__10167\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42835\
        );

    \I__10166\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42832\
        );

    \I__10165\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42825\
        );

    \I__10164\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42825\
        );

    \I__10163\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42825\
        );

    \I__10162\ : Odrv4
    port map (
            O => \N__42838\,
            I => \tx_transmit_N_1947_2\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__42835\,
            I => \tx_transmit_N_1947_2\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__42832\,
            I => \tx_transmit_N_1947_2\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__42825\,
            I => \tx_transmit_N_1947_2\
        );

    \I__10158\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42813\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__42813\,
            I => \N__42810\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__42810\,
            I => \c0.n13726\
        );

    \I__10155\ : SRMux
    port map (
            O => \N__42807\,
            I => \N__42803\
        );

    \I__10154\ : SRMux
    port map (
            O => \N__42806\,
            I => \N__42800\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__42803\,
            I => \N__42797\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__42800\,
            I => \N__42794\
        );

    \I__10151\ : Sp12to4
    port map (
            O => \N__42797\,
            I => \N__42790\
        );

    \I__10150\ : Span4Mux_h
    port map (
            O => \N__42794\,
            I => \N__42787\
        );

    \I__10149\ : SRMux
    port map (
            O => \N__42793\,
            I => \N__42784\
        );

    \I__10148\ : Span12Mux_s8_h
    port map (
            O => \N__42790\,
            I => \N__42781\
        );

    \I__10147\ : Span4Mux_h
    port map (
            O => \N__42787\,
            I => \N__42778\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__42784\,
            I => \N__42775\
        );

    \I__10145\ : Odrv12
    port map (
            O => \N__42781\,
            I => \c0.n10815\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__42778\,
            I => \c0.n10815\
        );

    \I__10143\ : Odrv12
    port map (
            O => \N__42775\,
            I => \c0.n10815\
        );

    \I__10142\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42765\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__42765\,
            I => \N__42762\
        );

    \I__10140\ : Span4Mux_h
    port map (
            O => \N__42762\,
            I => \N__42758\
        );

    \I__10139\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42755\
        );

    \I__10138\ : Span4Mux_v
    port map (
            O => \N__42758\,
            I => \N__42752\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__42755\,
            I => data_out_0_3
        );

    \I__10136\ : Odrv4
    port map (
            O => \N__42752\,
            I => data_out_0_3
        );

    \I__10135\ : InMux
    port map (
            O => \N__42747\,
            I => \c0.n16110\
        );

    \I__10134\ : InMux
    port map (
            O => \N__42744\,
            I => \c0.n16111\
        );

    \I__10133\ : InMux
    port map (
            O => \N__42741\,
            I => \c0.n16112\
        );

    \I__10132\ : InMux
    port map (
            O => \N__42738\,
            I => \c0.n16113\
        );

    \I__10131\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42731\
        );

    \I__10130\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42728\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__42731\,
            I => byte_transmit_counter_5
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__42728\,
            I => byte_transmit_counter_5
        );

    \I__10127\ : InMux
    port map (
            O => \N__42723\,
            I => \c0.n16114\
        );

    \I__10126\ : InMux
    port map (
            O => \N__42720\,
            I => \N__42717\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__42717\,
            I => \N__42713\
        );

    \I__10124\ : InMux
    port map (
            O => \N__42716\,
            I => \N__42710\
        );

    \I__10123\ : Span4Mux_v
    port map (
            O => \N__42713\,
            I => \N__42707\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__42710\,
            I => byte_transmit_counter_6
        );

    \I__10121\ : Odrv4
    port map (
            O => \N__42707\,
            I => byte_transmit_counter_6
        );

    \I__10120\ : InMux
    port map (
            O => \N__42702\,
            I => \c0.n16115\
        );

    \I__10119\ : InMux
    port map (
            O => \N__42699\,
            I => \N__42695\
        );

    \I__10118\ : InMux
    port map (
            O => \N__42698\,
            I => \N__42692\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__42695\,
            I => byte_transmit_counter_7
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__42692\,
            I => byte_transmit_counter_7
        );

    \I__10115\ : InMux
    port map (
            O => \N__42687\,
            I => \c0.n16116\
        );

    \I__10114\ : CascadeMux
    port map (
            O => \N__42684\,
            I => \n5_adj_2448_cascade_\
        );

    \I__10113\ : CascadeMux
    port map (
            O => \N__42681\,
            I => \n31_cascade_\
        );

    \I__10112\ : InMux
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__42675\,
            I => n22
        );

    \I__10110\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42667\
        );

    \I__10109\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42662\
        );

    \I__10108\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42662\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__42667\,
            I => n9524
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__42662\,
            I => n9524
        );

    \I__10105\ : InMux
    port map (
            O => \N__42657\,
            I => \N__42650\
        );

    \I__10104\ : InMux
    port map (
            O => \N__42656\,
            I => \N__42650\
        );

    \I__10103\ : InMux
    port map (
            O => \N__42655\,
            I => \N__42647\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__42650\,
            I => n450
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__42647\,
            I => n450
        );

    \I__10100\ : InMux
    port map (
            O => \N__42642\,
            I => \N__42637\
        );

    \I__10099\ : CascadeMux
    port map (
            O => \N__42641\,
            I => \N__42633\
        );

    \I__10098\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42630\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42627\
        );

    \I__10096\ : CascadeMux
    port map (
            O => \N__42636\,
            I => \N__42621\
        );

    \I__10095\ : InMux
    port map (
            O => \N__42633\,
            I => \N__42618\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__42630\,
            I => \N__42615\
        );

    \I__10093\ : Span4Mux_h
    port map (
            O => \N__42627\,
            I => \N__42612\
        );

    \I__10092\ : InMux
    port map (
            O => \N__42626\,
            I => \N__42607\
        );

    \I__10091\ : InMux
    port map (
            O => \N__42625\,
            I => \N__42607\
        );

    \I__10090\ : InMux
    port map (
            O => \N__42624\,
            I => \N__42602\
        );

    \I__10089\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42602\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__42618\,
            I => \r_Bit_Index_1\
        );

    \I__10087\ : Odrv4
    port map (
            O => \N__42615\,
            I => \r_Bit_Index_1\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__42612\,
            I => \r_Bit_Index_1\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__42607\,
            I => \r_Bit_Index_1\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__42602\,
            I => \r_Bit_Index_1\
        );

    \I__10083\ : CascadeMux
    port map (
            O => \N__42591\,
            I => \N__42588\
        );

    \I__10082\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42585\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__42585\,
            I => \N__42580\
        );

    \I__10080\ : InMux
    port map (
            O => \N__42584\,
            I => \N__42575\
        );

    \I__10079\ : InMux
    port map (
            O => \N__42583\,
            I => \N__42572\
        );

    \I__10078\ : Span4Mux_h
    port map (
            O => \N__42580\,
            I => \N__42569\
        );

    \I__10077\ : InMux
    port map (
            O => \N__42579\,
            I => \N__42564\
        );

    \I__10076\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42564\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__42575\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__42572\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__10073\ : Odrv4
    port map (
            O => \N__42569\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__42564\,
            I => \c0.tx.r_Bit_Index_0\
        );

    \I__10071\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42551\
        );

    \I__10070\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42547\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__42551\,
            I => \N__42543\
        );

    \I__10068\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42540\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__42547\,
            I => \N__42537\
        );

    \I__10066\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42534\
        );

    \I__10065\ : Span4Mux_h
    port map (
            O => \N__42543\,
            I => \N__42531\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__42540\,
            I => \r_Bit_Index_2\
        );

    \I__10063\ : Odrv4
    port map (
            O => \N__42537\,
            I => \r_Bit_Index_2\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__42534\,
            I => \r_Bit_Index_2\
        );

    \I__10061\ : Odrv4
    port map (
            O => \N__42531\,
            I => \r_Bit_Index_2\
        );

    \I__10060\ : CascadeMux
    port map (
            O => \N__42522\,
            I => \c0.tx.n17673_cascade_\
        );

    \I__10059\ : CascadeMux
    port map (
            O => \N__42519\,
            I => \N__42515\
        );

    \I__10058\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42512\
        );

    \I__10057\ : InMux
    port map (
            O => \N__42515\,
            I => \N__42509\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__42512\,
            I => \N__42506\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__42509\,
            I => \N__42503\
        );

    \I__10054\ : Span4Mux_h
    port map (
            O => \N__42506\,
            I => \N__42500\
        );

    \I__10053\ : Span4Mux_h
    port map (
            O => \N__42503\,
            I => \N__42497\
        );

    \I__10052\ : Odrv4
    port map (
            O => \N__42500\,
            I => \c0.n10326\
        );

    \I__10051\ : Odrv4
    port map (
            O => \N__42497\,
            I => \c0.n10326\
        );

    \I__10050\ : InMux
    port map (
            O => \N__42492\,
            I => \N__42489\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__42489\,
            I => \N__42486\
        );

    \I__10048\ : Span4Mux_h
    port map (
            O => \N__42486\,
            I => \N__42483\
        );

    \I__10047\ : Span4Mux_h
    port map (
            O => \N__42483\,
            I => \N__42480\
        );

    \I__10046\ : Odrv4
    port map (
            O => \N__42480\,
            I => \c0.n17126\
        );

    \I__10045\ : CascadeMux
    port map (
            O => \N__42477\,
            I => \c0.n17126_cascade_\
        );

    \I__10044\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42471\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__42471\,
            I => \N__42468\
        );

    \I__10042\ : Span4Mux_h
    port map (
            O => \N__42468\,
            I => \N__42465\
        );

    \I__10041\ : Odrv4
    port map (
            O => \N__42465\,
            I => \c0.n17651\
        );

    \I__10040\ : CascadeMux
    port map (
            O => \N__42462\,
            I => \N__42457\
        );

    \I__10039\ : CascadeMux
    port map (
            O => \N__42461\,
            I => \N__42453\
        );

    \I__10038\ : InMux
    port map (
            O => \N__42460\,
            I => \N__42449\
        );

    \I__10037\ : InMux
    port map (
            O => \N__42457\,
            I => \N__42443\
        );

    \I__10036\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42438\
        );

    \I__10035\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42438\
        );

    \I__10034\ : CascadeMux
    port map (
            O => \N__42452\,
            I => \N__42435\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__42449\,
            I => \N__42432\
        );

    \I__10032\ : CascadeMux
    port map (
            O => \N__42448\,
            I => \N__42429\
        );

    \I__10031\ : CascadeMux
    port map (
            O => \N__42447\,
            I => \N__42426\
        );

    \I__10030\ : CascadeMux
    port map (
            O => \N__42446\,
            I => \N__42423\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__42443\,
            I => \N__42418\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__42438\,
            I => \N__42418\
        );

    \I__10027\ : InMux
    port map (
            O => \N__42435\,
            I => \N__42415\
        );

    \I__10026\ : Span4Mux_v
    port map (
            O => \N__42432\,
            I => \N__42412\
        );

    \I__10025\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42405\
        );

    \I__10024\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42405\
        );

    \I__10023\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42405\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__42418\,
            I => \N__42402\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__42415\,
            I => \N__42399\
        );

    \I__10020\ : Span4Mux_v
    port map (
            O => \N__42412\,
            I => \N__42396\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__42405\,
            I => \N__42393\
        );

    \I__10018\ : Span4Mux_v
    port map (
            O => \N__42402\,
            I => \N__42390\
        );

    \I__10017\ : Span4Mux_h
    port map (
            O => \N__42399\,
            I => \N__42387\
        );

    \I__10016\ : Span4Mux_h
    port map (
            O => \N__42396\,
            I => \N__42382\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__42393\,
            I => \N__42382\
        );

    \I__10014\ : Span4Mux_h
    port map (
            O => \N__42390\,
            I => \N__42377\
        );

    \I__10013\ : Span4Mux_v
    port map (
            O => \N__42387\,
            I => \N__42377\
        );

    \I__10012\ : Span4Mux_v
    port map (
            O => \N__42382\,
            I => \N__42374\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__42377\,
            I => n10705
        );

    \I__10010\ : Odrv4
    port map (
            O => \N__42374\,
            I => n10705
        );

    \I__10009\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42358\
        );

    \I__10008\ : InMux
    port map (
            O => \N__42368\,
            I => \N__42358\
        );

    \I__10007\ : InMux
    port map (
            O => \N__42367\,
            I => \N__42358\
        );

    \I__10006\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42355\
        );

    \I__10005\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42352\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__42358\,
            I => \N__42345\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__42355\,
            I => \N__42345\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__42352\,
            I => \N__42342\
        );

    \I__10001\ : InMux
    port map (
            O => \N__42351\,
            I => \N__42339\
        );

    \I__10000\ : InMux
    port map (
            O => \N__42350\,
            I => \N__42336\
        );

    \I__9999\ : Odrv4
    port map (
            O => \N__42345\,
            I => n10_adj_2444
        );

    \I__9998\ : Odrv4
    port map (
            O => \N__42342\,
            I => n10_adj_2444
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__42339\,
            I => n10_adj_2444
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__42336\,
            I => n10_adj_2444
        );

    \I__9995\ : CascadeMux
    port map (
            O => \N__42327\,
            I => \n18187_cascade_\
        );

    \I__9994\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42320\
        );

    \I__9993\ : InMux
    port map (
            O => \N__42323\,
            I => \N__42317\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__42320\,
            I => \N__42312\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__42317\,
            I => \N__42312\
        );

    \I__9990\ : Odrv4
    port map (
            O => \N__42312\,
            I => \c0.data_out_6_6\
        );

    \I__9989\ : CascadeMux
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__9988\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42303\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__42303\,
            I => \c0.n5_adj_2159\
        );

    \I__9986\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42297\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__9984\ : Span4Mux_h
    port map (
            O => \N__42294\,
            I => \N__42290\
        );

    \I__9983\ : CascadeMux
    port map (
            O => \N__42293\,
            I => \N__42287\
        );

    \I__9982\ : Span4Mux_h
    port map (
            O => \N__42290\,
            I => \N__42284\
        );

    \I__9981\ : InMux
    port map (
            O => \N__42287\,
            I => \N__42281\
        );

    \I__9980\ : Odrv4
    port map (
            O => \N__42284\,
            I => rand_setpoint_30
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__42281\,
            I => rand_setpoint_30
        );

    \I__9978\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42273\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__42273\,
            I => \c0.n17698\
        );

    \I__9976\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42267\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__42267\,
            I => \c0.n17612\
        );

    \I__9974\ : CascadeMux
    port map (
            O => \N__42264\,
            I => \N__42261\
        );

    \I__9973\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42258\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__42258\,
            I => \N__42255\
        );

    \I__9971\ : Span4Mux_v
    port map (
            O => \N__42255\,
            I => \N__42252\
        );

    \I__9970\ : Span4Mux_h
    port map (
            O => \N__42252\,
            I => \N__42249\
        );

    \I__9969\ : Odrv4
    port map (
            O => \N__42249\,
            I => \c0.n17626\
        );

    \I__9968\ : CascadeMux
    port map (
            O => \N__42246\,
            I => \N__42243\
        );

    \I__9967\ : InMux
    port map (
            O => \N__42243\,
            I => \N__42240\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__42240\,
            I => \N__42237\
        );

    \I__9965\ : Span4Mux_h
    port map (
            O => \N__42237\,
            I => \N__42234\
        );

    \I__9964\ : Odrv4
    port map (
            O => \N__42234\,
            I => n25
        );

    \I__9963\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42228\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__42228\,
            I => \N__42225\
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__42225\,
            I => n28
        );

    \I__9960\ : SRMux
    port map (
            O => \N__42222\,
            I => \N__42219\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__42219\,
            I => \c0.n16704\
        );

    \I__9958\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42213\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__42213\,
            I => \N__42210\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__42210\,
            I => \c0.n3_adj_2193\
        );

    \I__9955\ : CascadeMux
    port map (
            O => \N__42207\,
            I => \N__42204\
        );

    \I__9954\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42201\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__42201\,
            I => \N__42198\
        );

    \I__9952\ : Span4Mux_h
    port map (
            O => \N__42198\,
            I => \N__42195\
        );

    \I__9951\ : Odrv4
    port map (
            O => \N__42195\,
            I => n10_adj_2431
        );

    \I__9950\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42189\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__42189\,
            I => \N__42186\
        );

    \I__9948\ : Span4Mux_v
    port map (
            O => \N__42186\,
            I => \N__42183\
        );

    \I__9947\ : Span4Mux_h
    port map (
            O => \N__42183\,
            I => \N__42180\
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__42180\,
            I => \c0.n6_adj_2221\
        );

    \I__9945\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42171\
        );

    \I__9944\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42171\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__42171\,
            I => \c0.n17147\
        );

    \I__9942\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42164\
        );

    \I__9941\ : CascadeMux
    port map (
            O => \N__42167\,
            I => \N__42161\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__42164\,
            I => \N__42158\
        );

    \I__9939\ : InMux
    port map (
            O => \N__42161\,
            I => \N__42155\
        );

    \I__9938\ : Odrv12
    port map (
            O => \N__42158\,
            I => rand_setpoint_8
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__42155\,
            I => rand_setpoint_8
        );

    \I__9936\ : InMux
    port map (
            O => \N__42150\,
            I => \N__42147\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__42147\,
            I => \c0.n17653\
        );

    \I__9934\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42140\
        );

    \I__9933\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42137\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__42140\,
            I => \N__42133\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__42137\,
            I => \N__42130\
        );

    \I__9930\ : InMux
    port map (
            O => \N__42136\,
            I => \N__42126\
        );

    \I__9929\ : Span4Mux_h
    port map (
            O => \N__42133\,
            I => \N__42123\
        );

    \I__9928\ : Span4Mux_v
    port map (
            O => \N__42130\,
            I => \N__42120\
        );

    \I__9927\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42117\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__42126\,
            I => data_out_8_1
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__42123\,
            I => data_out_8_1
        );

    \I__9924\ : Odrv4
    port map (
            O => \N__42120\,
            I => data_out_8_1
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__42117\,
            I => data_out_8_1
        );

    \I__9922\ : InMux
    port map (
            O => \N__42108\,
            I => \N__42105\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__42105\,
            I => \N__42102\
        );

    \I__9920\ : Odrv12
    port map (
            O => \N__42102\,
            I => \c0.n1_adj_2160\
        );

    \I__9919\ : CascadeMux
    port map (
            O => \N__42099\,
            I => \c0.n18184_cascade_\
        );

    \I__9918\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42090\
        );

    \I__9917\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42087\
        );

    \I__9916\ : InMux
    port map (
            O => \N__42094\,
            I => \N__42081\
        );

    \I__9915\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42078\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__42090\,
            I => \N__42075\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__42087\,
            I => \N__42072\
        );

    \I__9912\ : InMux
    port map (
            O => \N__42086\,
            I => \N__42069\
        );

    \I__9911\ : InMux
    port map (
            O => \N__42085\,
            I => \N__42066\
        );

    \I__9910\ : InMux
    port map (
            O => \N__42084\,
            I => \N__42063\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__42081\,
            I => \N__42060\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__42078\,
            I => \N__42057\
        );

    \I__9907\ : Span4Mux_v
    port map (
            O => \N__42075\,
            I => \N__42054\
        );

    \I__9906\ : Span4Mux_v
    port map (
            O => \N__42072\,
            I => \N__42050\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__42069\,
            I => \N__42047\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42044\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__42063\,
            I => \N__42041\
        );

    \I__9902\ : Span4Mux_h
    port map (
            O => \N__42060\,
            I => \N__42035\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__42057\,
            I => \N__42035\
        );

    \I__9900\ : Sp12to4
    port map (
            O => \N__42054\,
            I => \N__42032\
        );

    \I__9899\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42029\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__42050\,
            I => \N__42024\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__42047\,
            I => \N__42024\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__42044\,
            I => \N__42019\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__42041\,
            I => \N__42019\
        );

    \I__9894\ : InMux
    port map (
            O => \N__42040\,
            I => \N__42016\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__42035\,
            I => \N__42011\
        );

    \I__9892\ : Span12Mux_h
    port map (
            O => \N__42032\,
            I => \N__42006\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__42029\,
            I => \N__42006\
        );

    \I__9890\ : Span4Mux_h
    port map (
            O => \N__42024\,
            I => \N__42003\
        );

    \I__9889\ : Span4Mux_v
    port map (
            O => \N__42019\,
            I => \N__42000\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__42016\,
            I => \N__41997\
        );

    \I__9887\ : InMux
    port map (
            O => \N__42015\,
            I => \N__41994\
        );

    \I__9886\ : InMux
    port map (
            O => \N__42014\,
            I => \N__41991\
        );

    \I__9885\ : Odrv4
    port map (
            O => \N__42011\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9884\ : Odrv12
    port map (
            O => \N__42006\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9883\ : Odrv4
    port map (
            O => \N__42003\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__42000\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__41997\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__41994\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__41991\,
            I => \FRAME_MATCHER_i_31__N_1272\
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__41976\,
            I => \N__41973\
        );

    \I__9877\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41969\
        );

    \I__9876\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41964\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__41969\,
            I => \N__41961\
        );

    \I__9874\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41958\
        );

    \I__9873\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41953\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__41964\,
            I => \N__41950\
        );

    \I__9871\ : Span4Mux_h
    port map (
            O => \N__41961\,
            I => \N__41947\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__41958\,
            I => \N__41943\
        );

    \I__9869\ : InMux
    port map (
            O => \N__41957\,
            I => \N__41938\
        );

    \I__9868\ : InMux
    port map (
            O => \N__41956\,
            I => \N__41938\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__41953\,
            I => \N__41935\
        );

    \I__9866\ : Span4Mux_v
    port map (
            O => \N__41950\,
            I => \N__41932\
        );

    \I__9865\ : Span4Mux_v
    port map (
            O => \N__41947\,
            I => \N__41929\
        );

    \I__9864\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41926\
        );

    \I__9863\ : Span4Mux_h
    port map (
            O => \N__41943\,
            I => \N__41919\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__41938\,
            I => \N__41919\
        );

    \I__9861\ : Span4Mux_v
    port map (
            O => \N__41935\,
            I => \N__41919\
        );

    \I__9860\ : Span4Mux_v
    port map (
            O => \N__41932\,
            I => \N__41916\
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__41929\,
            I => n488
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__41926\,
            I => n488
        );

    \I__9857\ : Odrv4
    port map (
            O => \N__41919\,
            I => n488
        );

    \I__9856\ : Odrv4
    port map (
            O => \N__41916\,
            I => n488
        );

    \I__9855\ : InMux
    port map (
            O => \N__41907\,
            I => \N__41892\
        );

    \I__9854\ : InMux
    port map (
            O => \N__41906\,
            I => \N__41892\
        );

    \I__9853\ : InMux
    port map (
            O => \N__41905\,
            I => \N__41892\
        );

    \I__9852\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41892\
        );

    \I__9851\ : InMux
    port map (
            O => \N__41903\,
            I => \N__41892\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__41892\,
            I => \N__41855\
        );

    \I__9849\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41825\
        );

    \I__9848\ : InMux
    port map (
            O => \N__41890\,
            I => \N__41825\
        );

    \I__9847\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41825\
        );

    \I__9846\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41825\
        );

    \I__9845\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41825\
        );

    \I__9844\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41814\
        );

    \I__9843\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41814\
        );

    \I__9842\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41814\
        );

    \I__9841\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41814\
        );

    \I__9840\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41814\
        );

    \I__9839\ : InMux
    port map (
            O => \N__41881\,
            I => \N__41801\
        );

    \I__9838\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41801\
        );

    \I__9837\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41801\
        );

    \I__9836\ : InMux
    port map (
            O => \N__41878\,
            I => \N__41801\
        );

    \I__9835\ : InMux
    port map (
            O => \N__41877\,
            I => \N__41801\
        );

    \I__9834\ : InMux
    port map (
            O => \N__41876\,
            I => \N__41801\
        );

    \I__9833\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41794\
        );

    \I__9832\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41794\
        );

    \I__9831\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41794\
        );

    \I__9830\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41779\
        );

    \I__9829\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41779\
        );

    \I__9828\ : InMux
    port map (
            O => \N__41870\,
            I => \N__41779\
        );

    \I__9827\ : InMux
    port map (
            O => \N__41869\,
            I => \N__41779\
        );

    \I__9826\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41779\
        );

    \I__9825\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41779\
        );

    \I__9824\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41779\
        );

    \I__9823\ : InMux
    port map (
            O => \N__41865\,
            I => \N__41766\
        );

    \I__9822\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41766\
        );

    \I__9821\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41766\
        );

    \I__9820\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41766\
        );

    \I__9819\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41766\
        );

    \I__9818\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41766\
        );

    \I__9817\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41760\
        );

    \I__9816\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41760\
        );

    \I__9815\ : Span4Mux_v
    port map (
            O => \N__41855\,
            I => \N__41757\
        );

    \I__9814\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41742\
        );

    \I__9813\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41742\
        );

    \I__9812\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41742\
        );

    \I__9811\ : InMux
    port map (
            O => \N__41851\,
            I => \N__41742\
        );

    \I__9810\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41742\
        );

    \I__9809\ : InMux
    port map (
            O => \N__41849\,
            I => \N__41742\
        );

    \I__9808\ : InMux
    port map (
            O => \N__41848\,
            I => \N__41742\
        );

    \I__9807\ : InMux
    port map (
            O => \N__41847\,
            I => \N__41730\
        );

    \I__9806\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41730\
        );

    \I__9805\ : InMux
    port map (
            O => \N__41845\,
            I => \N__41730\
        );

    \I__9804\ : InMux
    port map (
            O => \N__41844\,
            I => \N__41730\
        );

    \I__9803\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41730\
        );

    \I__9802\ : InMux
    port map (
            O => \N__41842\,
            I => \N__41715\
        );

    \I__9801\ : InMux
    port map (
            O => \N__41841\,
            I => \N__41715\
        );

    \I__9800\ : InMux
    port map (
            O => \N__41840\,
            I => \N__41715\
        );

    \I__9799\ : InMux
    port map (
            O => \N__41839\,
            I => \N__41715\
        );

    \I__9798\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41715\
        );

    \I__9797\ : InMux
    port map (
            O => \N__41837\,
            I => \N__41715\
        );

    \I__9796\ : InMux
    port map (
            O => \N__41836\,
            I => \N__41715\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__41825\,
            I => \N__41704\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__41814\,
            I => \N__41704\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__41801\,
            I => \N__41704\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__41794\,
            I => \N__41704\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__41779\,
            I => \N__41704\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__41766\,
            I => \N__41701\
        );

    \I__9789\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41697\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__41760\,
            I => \N__41694\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__41757\,
            I => \N__41689\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__41742\,
            I => \N__41689\
        );

    \I__9785\ : InMux
    port map (
            O => \N__41741\,
            I => \N__41686\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__41730\,
            I => \N__41683\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__41715\,
            I => \N__41676\
        );

    \I__9782\ : Span4Mux_v
    port map (
            O => \N__41704\,
            I => \N__41676\
        );

    \I__9781\ : Span4Mux_h
    port map (
            O => \N__41701\,
            I => \N__41676\
        );

    \I__9780\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41665\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41662\
        );

    \I__9778\ : Span4Mux_h
    port map (
            O => \N__41694\,
            I => \N__41657\
        );

    \I__9777\ : Span4Mux_v
    port map (
            O => \N__41689\,
            I => \N__41657\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__41686\,
            I => \N__41654\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__41683\,
            I => \N__41649\
        );

    \I__9774\ : Span4Mux_h
    port map (
            O => \N__41676\,
            I => \N__41649\
        );

    \I__9773\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41636\
        );

    \I__9772\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41636\
        );

    \I__9771\ : InMux
    port map (
            O => \N__41673\,
            I => \N__41636\
        );

    \I__9770\ : InMux
    port map (
            O => \N__41672\,
            I => \N__41636\
        );

    \I__9769\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41636\
        );

    \I__9768\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41636\
        );

    \I__9767\ : InMux
    port map (
            O => \N__41669\,
            I => \N__41633\
        );

    \I__9766\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41630\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__41665\,
            I => \c0.n13146\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__41662\,
            I => \c0.n13146\
        );

    \I__9763\ : Odrv4
    port map (
            O => \N__41657\,
            I => \c0.n13146\
        );

    \I__9762\ : Odrv4
    port map (
            O => \N__41654\,
            I => \c0.n13146\
        );

    \I__9761\ : Odrv4
    port map (
            O => \N__41649\,
            I => \c0.n13146\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__41636\,
            I => \c0.n13146\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__41633\,
            I => \c0.n13146\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__41630\,
            I => \c0.n13146\
        );

    \I__9757\ : CascadeMux
    port map (
            O => \N__41613\,
            I => \N__41610\
        );

    \I__9756\ : InMux
    port map (
            O => \N__41610\,
            I => \N__41607\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__41607\,
            I => \N__41602\
        );

    \I__9754\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41599\
        );

    \I__9753\ : InMux
    port map (
            O => \N__41605\,
            I => \N__41596\
        );

    \I__9752\ : Span4Mux_v
    port map (
            O => \N__41602\,
            I => \N__41593\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__41599\,
            I => \N__41589\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__41596\,
            I => \N__41586\
        );

    \I__9749\ : Span4Mux_h
    port map (
            O => \N__41593\,
            I => \N__41583\
        );

    \I__9748\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41580\
        );

    \I__9747\ : Span4Mux_v
    port map (
            O => \N__41589\,
            I => \N__41577\
        );

    \I__9746\ : Sp12to4
    port map (
            O => \N__41586\,
            I => \N__41570\
        );

    \I__9745\ : Sp12to4
    port map (
            O => \N__41583\,
            I => \N__41570\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__41580\,
            I => \N__41570\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__41577\,
            I => \N__41567\
        );

    \I__9742\ : Span12Mux_h
    port map (
            O => \N__41570\,
            I => \N__41564\
        );

    \I__9741\ : Odrv4
    port map (
            O => \N__41567\,
            I => n4408
        );

    \I__9740\ : Odrv12
    port map (
            O => \N__41564\,
            I => n4408
        );

    \I__9739\ : CascadeMux
    port map (
            O => \N__41559\,
            I => \c0.n276_cascade_\
        );

    \I__9738\ : InMux
    port map (
            O => \N__41556\,
            I => \N__41553\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__41553\,
            I => \N__41549\
        );

    \I__9736\ : InMux
    port map (
            O => \N__41552\,
            I => \N__41546\
        );

    \I__9735\ : Span12Mux_h
    port map (
            O => \N__41549\,
            I => \N__41542\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__41546\,
            I => \N__41539\
        );

    \I__9733\ : InMux
    port map (
            O => \N__41545\,
            I => \N__41536\
        );

    \I__9732\ : Odrv12
    port map (
            O => \N__41542\,
            I => \c0.n4_adj_2135\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__41539\,
            I => \c0.n4_adj_2135\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__41536\,
            I => \c0.n4_adj_2135\
        );

    \I__9729\ : CascadeMux
    port map (
            O => \N__41529\,
            I => \c0.n4_adj_2135_cascade_\
        );

    \I__9728\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41519\
        );

    \I__9727\ : InMux
    port map (
            O => \N__41525\,
            I => \N__41519\
        );

    \I__9726\ : InMux
    port map (
            O => \N__41524\,
            I => \N__41516\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__41519\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__41516\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__9723\ : SRMux
    port map (
            O => \N__41511\,
            I => \N__41508\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__41508\,
            I => \N__41505\
        );

    \I__9721\ : Span4Mux_h
    port map (
            O => \N__41505\,
            I => \N__41502\
        );

    \I__9720\ : Odrv4
    port map (
            O => \N__41502\,
            I => \c0.n16700\
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__41499\,
            I => \N__41495\
        );

    \I__9718\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41482\
        );

    \I__9717\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41482\
        );

    \I__9716\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41482\
        );

    \I__9715\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41482\
        );

    \I__9714\ : CascadeMux
    port map (
            O => \N__41492\,
            I => \N__41479\
        );

    \I__9713\ : CascadeMux
    port map (
            O => \N__41491\,
            I => \N__41475\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__41482\,
            I => \N__41469\
        );

    \I__9711\ : InMux
    port map (
            O => \N__41479\,
            I => \N__41458\
        );

    \I__9710\ : InMux
    port map (
            O => \N__41478\,
            I => \N__41458\
        );

    \I__9709\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41458\
        );

    \I__9708\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41458\
        );

    \I__9707\ : InMux
    port map (
            O => \N__41473\,
            I => \N__41458\
        );

    \I__9706\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41454\
        );

    \I__9705\ : Span4Mux_h
    port map (
            O => \N__41469\,
            I => \N__41449\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__41458\,
            I => \N__41449\
        );

    \I__9703\ : InMux
    port map (
            O => \N__41457\,
            I => \N__41446\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__41454\,
            I => \N__41442\
        );

    \I__9701\ : Span4Mux_h
    port map (
            O => \N__41449\,
            I => \N__41437\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__41446\,
            I => \N__41437\
        );

    \I__9699\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41434\
        );

    \I__9698\ : Odrv4
    port map (
            O => \N__41442\,
            I => \c0.n9334\
        );

    \I__9697\ : Odrv4
    port map (
            O => \N__41437\,
            I => \c0.n9334\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__41434\,
            I => \c0.n9334\
        );

    \I__9695\ : CascadeMux
    port map (
            O => \N__41427\,
            I => \N__41424\
        );

    \I__9694\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41414\
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__41423\,
            I => \N__41411\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__41422\,
            I => \N__41408\
        );

    \I__9691\ : CascadeMux
    port map (
            O => \N__41421\,
            I => \N__41404\
        );

    \I__9690\ : CascadeMux
    port map (
            O => \N__41420\,
            I => \N__41401\
        );

    \I__9689\ : CascadeMux
    port map (
            O => \N__41419\,
            I => \N__41397\
        );

    \I__9688\ : CascadeMux
    port map (
            O => \N__41418\,
            I => \N__41393\
        );

    \I__9687\ : CascadeMux
    port map (
            O => \N__41417\,
            I => \N__41390\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41386\
        );

    \I__9685\ : InMux
    port map (
            O => \N__41411\,
            I => \N__41383\
        );

    \I__9684\ : InMux
    port map (
            O => \N__41408\,
            I => \N__41374\
        );

    \I__9683\ : InMux
    port map (
            O => \N__41407\,
            I => \N__41374\
        );

    \I__9682\ : InMux
    port map (
            O => \N__41404\,
            I => \N__41374\
        );

    \I__9681\ : InMux
    port map (
            O => \N__41401\,
            I => \N__41374\
        );

    \I__9680\ : InMux
    port map (
            O => \N__41400\,
            I => \N__41363\
        );

    \I__9679\ : InMux
    port map (
            O => \N__41397\,
            I => \N__41363\
        );

    \I__9678\ : InMux
    port map (
            O => \N__41396\,
            I => \N__41363\
        );

    \I__9677\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41363\
        );

    \I__9676\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41363\
        );

    \I__9675\ : InMux
    port map (
            O => \N__41389\,
            I => \N__41359\
        );

    \I__9674\ : Span4Mux_h
    port map (
            O => \N__41386\,
            I => \N__41354\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__41383\,
            I => \N__41354\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__41374\,
            I => \N__41349\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__41363\,
            I => \N__41349\
        );

    \I__9670\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41346\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__41359\,
            I => n44
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__41354\,
            I => n44
        );

    \I__9667\ : Odrv4
    port map (
            O => \N__41349\,
            I => n44
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__41346\,
            I => n44
        );

    \I__9665\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41323\
        );

    \I__9664\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41323\
        );

    \I__9663\ : InMux
    port map (
            O => \N__41335\,
            I => \N__41323\
        );

    \I__9662\ : InMux
    port map (
            O => \N__41334\,
            I => \N__41323\
        );

    \I__9661\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41315\
        );

    \I__9660\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41312\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41309\
        );

    \I__9658\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41298\
        );

    \I__9657\ : InMux
    port map (
            O => \N__41321\,
            I => \N__41298\
        );

    \I__9656\ : InMux
    port map (
            O => \N__41320\,
            I => \N__41298\
        );

    \I__9655\ : InMux
    port map (
            O => \N__41319\,
            I => \N__41298\
        );

    \I__9654\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41298\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__41315\,
            I => \N__41293\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__41312\,
            I => \N__41290\
        );

    \I__9651\ : Span4Mux_h
    port map (
            O => \N__41309\,
            I => \N__41285\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__41298\,
            I => \N__41285\
        );

    \I__9649\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41282\
        );

    \I__9648\ : InMux
    port map (
            O => \N__41296\,
            I => \N__41279\
        );

    \I__9647\ : Odrv4
    port map (
            O => \N__41293\,
            I => \c0.n17069\
        );

    \I__9646\ : Odrv4
    port map (
            O => \N__41290\,
            I => \c0.n17069\
        );

    \I__9645\ : Odrv4
    port map (
            O => \N__41285\,
            I => \c0.n17069\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__41282\,
            I => \c0.n17069\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__41279\,
            I => \c0.n17069\
        );

    \I__9642\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41265\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__41265\,
            I => \N__41260\
        );

    \I__9640\ : CascadeMux
    port map (
            O => \N__41264\,
            I => \N__41257\
        );

    \I__9639\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41254\
        );

    \I__9638\ : Span4Mux_v
    port map (
            O => \N__41260\,
            I => \N__41251\
        );

    \I__9637\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41248\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__41254\,
            I => \N__41245\
        );

    \I__9635\ : Span4Mux_h
    port map (
            O => \N__41251\,
            I => \N__41242\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__41248\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__41245\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__9632\ : Odrv4
    port map (
            O => \N__41242\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__9631\ : CascadeMux
    port map (
            O => \N__41235\,
            I => \N__41232\
        );

    \I__9630\ : InMux
    port map (
            O => \N__41232\,
            I => \N__41229\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__41229\,
            I => \N__41224\
        );

    \I__9628\ : InMux
    port map (
            O => \N__41228\,
            I => \N__41221\
        );

    \I__9627\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41218\
        );

    \I__9626\ : Span4Mux_h
    port map (
            O => \N__41224\,
            I => \N__41215\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__41221\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__41218\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__41215\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__9622\ : SRMux
    port map (
            O => \N__41208\,
            I => \N__41205\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__41205\,
            I => \N__41202\
        );

    \I__9620\ : Span4Mux_v
    port map (
            O => \N__41202\,
            I => \N__41199\
        );

    \I__9619\ : Span4Mux_h
    port map (
            O => \N__41199\,
            I => \N__41196\
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__41196\,
            I => \c0.n16658\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__41193\,
            I => \N__41189\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__41192\,
            I => \N__41185\
        );

    \I__9615\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41182\
        );

    \I__9614\ : InMux
    port map (
            O => \N__41188\,
            I => \N__41179\
        );

    \I__9613\ : InMux
    port map (
            O => \N__41185\,
            I => \N__41176\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__41182\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__41179\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__41176\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__9609\ : SRMux
    port map (
            O => \N__41169\,
            I => \N__41166\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__41166\,
            I => \N__41163\
        );

    \I__9607\ : Span4Mux_h
    port map (
            O => \N__41163\,
            I => \N__41160\
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__41160\,
            I => \c0.n16710\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__41157\,
            I => \N__41153\
        );

    \I__9604\ : InMux
    port map (
            O => \N__41156\,
            I => \N__41150\
        );

    \I__9603\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41146\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__41150\,
            I => \N__41141\
        );

    \I__9601\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41138\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__41146\,
            I => \N__41135\
        );

    \I__9599\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41132\
        );

    \I__9598\ : InMux
    port map (
            O => \N__41144\,
            I => \N__41129\
        );

    \I__9597\ : Span4Mux_h
    port map (
            O => \N__41141\,
            I => \N__41126\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__41138\,
            I => \N__41123\
        );

    \I__9595\ : Span12Mux_v
    port map (
            O => \N__41135\,
            I => \N__41118\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__41132\,
            I => \N__41118\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__41129\,
            I => data_out_frame2_13_4
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__41126\,
            I => data_out_frame2_13_4
        );

    \I__9591\ : Odrv12
    port map (
            O => \N__41123\,
            I => data_out_frame2_13_4
        );

    \I__9590\ : Odrv12
    port map (
            O => \N__41118\,
            I => data_out_frame2_13_4
        );

    \I__9589\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41102\
        );

    \I__9588\ : InMux
    port map (
            O => \N__41108\,
            I => \N__41099\
        );

    \I__9587\ : InMux
    port map (
            O => \N__41107\,
            I => \N__41093\
        );

    \I__9586\ : InMux
    port map (
            O => \N__41106\,
            I => \N__41093\
        );

    \I__9585\ : CascadeMux
    port map (
            O => \N__41105\,
            I => \N__41090\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__41102\,
            I => \N__41087\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__41099\,
            I => \N__41084\
        );

    \I__9582\ : InMux
    port map (
            O => \N__41098\,
            I => \N__41081\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41078\
        );

    \I__9580\ : InMux
    port map (
            O => \N__41090\,
            I => \N__41075\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__41087\,
            I => \N__41072\
        );

    \I__9578\ : Span4Mux_v
    port map (
            O => \N__41084\,
            I => \N__41065\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__41081\,
            I => \N__41065\
        );

    \I__9576\ : Span4Mux_v
    port map (
            O => \N__41078\,
            I => \N__41065\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__41075\,
            I => \N__41060\
        );

    \I__9574\ : Span4Mux_h
    port map (
            O => \N__41072\,
            I => \N__41060\
        );

    \I__9573\ : Odrv4
    port map (
            O => \N__41065\,
            I => data_out_frame2_9_0
        );

    \I__9572\ : Odrv4
    port map (
            O => \N__41060\,
            I => data_out_frame2_9_0
        );

    \I__9571\ : CascadeMux
    port map (
            O => \N__41055\,
            I => \N__41052\
        );

    \I__9570\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41049\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__41049\,
            I => \N__41046\
        );

    \I__9568\ : Span4Mux_v
    port map (
            O => \N__41046\,
            I => \N__41043\
        );

    \I__9567\ : Span4Mux_h
    port map (
            O => \N__41043\,
            I => \N__41040\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__41040\,
            I => \N__41037\
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__41037\,
            I => \c0.n17315\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__41034\,
            I => \N__41027\
        );

    \I__9563\ : InMux
    port map (
            O => \N__41033\,
            I => \N__41024\
        );

    \I__9562\ : InMux
    port map (
            O => \N__41032\,
            I => \N__41021\
        );

    \I__9561\ : InMux
    port map (
            O => \N__41031\,
            I => \N__41018\
        );

    \I__9560\ : InMux
    port map (
            O => \N__41030\,
            I => \N__41015\
        );

    \I__9559\ : InMux
    port map (
            O => \N__41027\,
            I => \N__41012\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__41024\,
            I => \N__41009\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__41021\,
            I => \N__41006\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__41018\,
            I => \N__41003\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41000\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__41012\,
            I => \c0.data_in_frame_0_0\
        );

    \I__9553\ : Odrv12
    port map (
            O => \N__41009\,
            I => \c0.data_in_frame_0_0\
        );

    \I__9552\ : Odrv4
    port map (
            O => \N__41006\,
            I => \c0.data_in_frame_0_0\
        );

    \I__9551\ : Odrv4
    port map (
            O => \N__41003\,
            I => \c0.data_in_frame_0_0\
        );

    \I__9550\ : Odrv4
    port map (
            O => \N__41000\,
            I => \c0.data_in_frame_0_0\
        );

    \I__9549\ : CascadeMux
    port map (
            O => \N__40989\,
            I => \N__40985\
        );

    \I__9548\ : InMux
    port map (
            O => \N__40988\,
            I => \N__40979\
        );

    \I__9547\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40979\
        );

    \I__9546\ : CascadeMux
    port map (
            O => \N__40984\,
            I => \N__40975\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40972\
        );

    \I__9544\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40969\
        );

    \I__9543\ : InMux
    port map (
            O => \N__40975\,
            I => \N__40966\
        );

    \I__9542\ : Span4Mux_h
    port map (
            O => \N__40972\,
            I => \N__40963\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__40969\,
            I => \N__40960\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__40966\,
            I => \c0.data_in_frame_1_7\
        );

    \I__9539\ : Odrv4
    port map (
            O => \N__40963\,
            I => \c0.data_in_frame_1_7\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__40960\,
            I => \c0.data_in_frame_1_7\
        );

    \I__9537\ : InMux
    port map (
            O => \N__40953\,
            I => \N__40947\
        );

    \I__9536\ : InMux
    port map (
            O => \N__40952\,
            I => \N__40947\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__40947\,
            I => \N__40944\
        );

    \I__9534\ : Span4Mux_h
    port map (
            O => \N__40944\,
            I => \N__40941\
        );

    \I__9533\ : Odrv4
    port map (
            O => \N__40941\,
            I => \c0.n17213\
        );

    \I__9532\ : CascadeMux
    port map (
            O => \N__40938\,
            I => \N__40935\
        );

    \I__9531\ : InMux
    port map (
            O => \N__40935\,
            I => \N__40930\
        );

    \I__9530\ : CascadeMux
    port map (
            O => \N__40934\,
            I => \N__40926\
        );

    \I__9529\ : InMux
    port map (
            O => \N__40933\,
            I => \N__40922\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__40930\,
            I => \N__40919\
        );

    \I__9527\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40914\
        );

    \I__9526\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40914\
        );

    \I__9525\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40911\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__40922\,
            I => \N__40908\
        );

    \I__9523\ : Span4Mux_v
    port map (
            O => \N__40919\,
            I => \N__40903\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__40914\,
            I => \N__40903\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__40911\,
            I => data_out_frame2_8_5
        );

    \I__9520\ : Odrv12
    port map (
            O => \N__40908\,
            I => data_out_frame2_8_5
        );

    \I__9519\ : Odrv4
    port map (
            O => \N__40903\,
            I => data_out_frame2_8_5
        );

    \I__9518\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40893\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__40893\,
            I => \N__40888\
        );

    \I__9516\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40885\
        );

    \I__9515\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40882\
        );

    \I__9514\ : Span4Mux_v
    port map (
            O => \N__40888\,
            I => \N__40879\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__40885\,
            I => \N__40876\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__40882\,
            I => \N__40873\
        );

    \I__9511\ : Span4Mux_h
    port map (
            O => \N__40879\,
            I => \N__40868\
        );

    \I__9510\ : Span4Mux_v
    port map (
            O => \N__40876\,
            I => \N__40868\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__40873\,
            I => \N__40865\
        );

    \I__9508\ : Span4Mux_h
    port map (
            O => \N__40868\,
            I => \N__40858\
        );

    \I__9507\ : Span4Mux_h
    port map (
            O => \N__40865\,
            I => \N__40858\
        );

    \I__9506\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40855\
        );

    \I__9505\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40852\
        );

    \I__9504\ : Sp12to4
    port map (
            O => \N__40858\,
            I => \N__40849\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__40855\,
            I => data_out_frame2_6_6
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__40852\,
            I => data_out_frame2_6_6
        );

    \I__9501\ : Odrv12
    port map (
            O => \N__40849\,
            I => data_out_frame2_6_6
        );

    \I__9500\ : CascadeMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__9499\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40836\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__40836\,
            I => \N__40833\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__40833\,
            I => \N__40830\
        );

    \I__9496\ : Sp12to4
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__9495\ : Span12Mux_s5_h
    port map (
            O => \N__40827\,
            I => \N__40824\
        );

    \I__9494\ : Odrv12
    port map (
            O => \N__40824\,
            I => \c0.n10472\
        );

    \I__9493\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40815\
        );

    \I__9492\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40815\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__40815\,
            I => \N__40811\
        );

    \I__9490\ : InMux
    port map (
            O => \N__40814\,
            I => \N__40808\
        );

    \I__9489\ : Span4Mux_v
    port map (
            O => \N__40811\,
            I => \N__40802\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__40808\,
            I => \N__40802\
        );

    \I__9487\ : InMux
    port map (
            O => \N__40807\,
            I => \N__40799\
        );

    \I__9486\ : Span4Mux_h
    port map (
            O => \N__40802\,
            I => \N__40789\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__40799\,
            I => \N__40786\
        );

    \I__9484\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40773\
        );

    \I__9483\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40773\
        );

    \I__9482\ : InMux
    port map (
            O => \N__40796\,
            I => \N__40773\
        );

    \I__9481\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40773\
        );

    \I__9480\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40773\
        );

    \I__9479\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40773\
        );

    \I__9478\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40770\
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__40789\,
            I => \c0.n15821\
        );

    \I__9476\ : Odrv4
    port map (
            O => \N__40786\,
            I => \c0.n15821\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__40773\,
            I => \c0.n15821\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__40770\,
            I => \c0.n15821\
        );

    \I__9473\ : CascadeMux
    port map (
            O => \N__40761\,
            I => \N__40756\
        );

    \I__9472\ : CascadeMux
    port map (
            O => \N__40760\,
            I => \N__40753\
        );

    \I__9471\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40750\
        );

    \I__9470\ : InMux
    port map (
            O => \N__40756\,
            I => \N__40747\
        );

    \I__9469\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40744\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__40750\,
            I => \N__40741\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__40747\,
            I => \N__40738\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__40744\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__40741\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__40738\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__9463\ : SRMux
    port map (
            O => \N__40731\,
            I => \N__40728\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__40728\,
            I => \N__40725\
        );

    \I__9461\ : Span4Mux_h
    port map (
            O => \N__40725\,
            I => \N__40722\
        );

    \I__9460\ : Odrv4
    port map (
            O => \N__40722\,
            I => \c0.n8_adj_2329\
        );

    \I__9459\ : InMux
    port map (
            O => \N__40719\,
            I => \N__40715\
        );

    \I__9458\ : InMux
    port map (
            O => \N__40718\,
            I => \N__40712\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__40715\,
            I => \N__40706\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__40712\,
            I => \N__40706\
        );

    \I__9455\ : CascadeMux
    port map (
            O => \N__40711\,
            I => \N__40703\
        );

    \I__9454\ : Span4Mux_h
    port map (
            O => \N__40706\,
            I => \N__40699\
        );

    \I__9453\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40694\
        );

    \I__9452\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40694\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__40699\,
            I => \c0.n8_adj_2385\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__40694\,
            I => \c0.n8_adj_2385\
        );

    \I__9449\ : InMux
    port map (
            O => \N__40689\,
            I => \N__40686\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__40686\,
            I => \N__40683\
        );

    \I__9447\ : Odrv12
    port map (
            O => \N__40683\,
            I => \c0.n46\
        );

    \I__9446\ : CascadeMux
    port map (
            O => \N__40680\,
            I => \N__40677\
        );

    \I__9445\ : InMux
    port map (
            O => \N__40677\,
            I => \N__40674\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__40674\,
            I => \N__40669\
        );

    \I__9443\ : InMux
    port map (
            O => \N__40673\,
            I => \N__40664\
        );

    \I__9442\ : InMux
    port map (
            O => \N__40672\,
            I => \N__40664\
        );

    \I__9441\ : Span4Mux_h
    port map (
            O => \N__40669\,
            I => \N__40660\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__40664\,
            I => \N__40657\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__40663\,
            I => \N__40654\
        );

    \I__9438\ : Sp12to4
    port map (
            O => \N__40660\,
            I => \N__40651\
        );

    \I__9437\ : Span4Mux_h
    port map (
            O => \N__40657\,
            I => \N__40648\
        );

    \I__9436\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40645\
        );

    \I__9435\ : Span12Mux_v
    port map (
            O => \N__40651\,
            I => \N__40642\
        );

    \I__9434\ : Span4Mux_h
    port map (
            O => \N__40648\,
            I => \N__40639\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__40645\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9432\ : Odrv12
    port map (
            O => \N__40642\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__40639\,
            I => \c0.data_out_frame2_0_0\
        );

    \I__9430\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40629\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__40629\,
            I => \c0.n17490\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__40626\,
            I => \N__40620\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__40625\,
            I => \N__40615\
        );

    \I__9426\ : CascadeMux
    port map (
            O => \N__40624\,
            I => \N__40611\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__40623\,
            I => \N__40607\
        );

    \I__9424\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40601\
        );

    \I__9423\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40601\
        );

    \I__9422\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40595\
        );

    \I__9421\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40592\
        );

    \I__9420\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40587\
        );

    \I__9419\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40587\
        );

    \I__9418\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40584\
        );

    \I__9417\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40579\
        );

    \I__9416\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40579\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__40601\,
            I => \N__40574\
        );

    \I__9414\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40571\
        );

    \I__9413\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40568\
        );

    \I__9412\ : InMux
    port map (
            O => \N__40598\,
            I => \N__40564\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__40595\,
            I => \N__40561\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__40592\,
            I => \N__40558\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__40587\,
            I => \N__40553\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__40584\,
            I => \N__40553\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__40579\,
            I => \N__40550\
        );

    \I__9406\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40545\
        );

    \I__9405\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40545\
        );

    \I__9404\ : Span4Mux_v
    port map (
            O => \N__40574\,
            I => \N__40538\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__40571\,
            I => \N__40538\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__40568\,
            I => \N__40538\
        );

    \I__9401\ : InMux
    port map (
            O => \N__40567\,
            I => \N__40535\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__40564\,
            I => \N__40528\
        );

    \I__9399\ : Span4Mux_v
    port map (
            O => \N__40561\,
            I => \N__40528\
        );

    \I__9398\ : Span4Mux_v
    port map (
            O => \N__40558\,
            I => \N__40528\
        );

    \I__9397\ : Span4Mux_h
    port map (
            O => \N__40553\,
            I => \N__40525\
        );

    \I__9396\ : Span4Mux_v
    port map (
            O => \N__40550\,
            I => \N__40518\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__40545\,
            I => \N__40518\
        );

    \I__9394\ : Span4Mux_v
    port map (
            O => \N__40538\,
            I => \N__40518\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__40535\,
            I => \c0.n15171\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__40528\,
            I => \c0.n15171\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__40525\,
            I => \c0.n15171\
        );

    \I__9390\ : Odrv4
    port map (
            O => \N__40518\,
            I => \c0.n15171\
        );

    \I__9389\ : CascadeMux
    port map (
            O => \N__40509\,
            I => \N__40506\
        );

    \I__9388\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40496\
        );

    \I__9387\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40493\
        );

    \I__9386\ : InMux
    port map (
            O => \N__40504\,
            I => \N__40490\
        );

    \I__9385\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40487\
        );

    \I__9384\ : CascadeMux
    port map (
            O => \N__40502\,
            I => \N__40484\
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__40501\,
            I => \N__40481\
        );

    \I__9382\ : InMux
    port map (
            O => \N__40500\,
            I => \N__40478\
        );

    \I__9381\ : InMux
    port map (
            O => \N__40499\,
            I => \N__40475\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__40496\,
            I => \N__40472\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__40493\,
            I => \N__40467\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__40490\,
            I => \N__40467\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__40487\,
            I => \N__40464\
        );

    \I__9376\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40461\
        );

    \I__9375\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40458\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__40478\,
            I => \N__40455\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__40475\,
            I => \N__40450\
        );

    \I__9372\ : Span4Mux_h
    port map (
            O => \N__40472\,
            I => \N__40450\
        );

    \I__9371\ : Span4Mux_v
    port map (
            O => \N__40467\,
            I => \N__40445\
        );

    \I__9370\ : Span4Mux_v
    port map (
            O => \N__40464\,
            I => \N__40445\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__40461\,
            I => rx_data_7
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__40458\,
            I => rx_data_7
        );

    \I__9367\ : Odrv12
    port map (
            O => \N__40455\,
            I => rx_data_7
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__40450\,
            I => rx_data_7
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__40445\,
            I => rx_data_7
        );

    \I__9364\ : CascadeMux
    port map (
            O => \N__40434\,
            I => \N__40415\
        );

    \I__9363\ : CascadeMux
    port map (
            O => \N__40433\,
            I => \N__40412\
        );

    \I__9362\ : InMux
    port map (
            O => \N__40432\,
            I => \N__40403\
        );

    \I__9361\ : InMux
    port map (
            O => \N__40431\,
            I => \N__40400\
        );

    \I__9360\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40397\
        );

    \I__9359\ : InMux
    port map (
            O => \N__40429\,
            I => \N__40390\
        );

    \I__9358\ : InMux
    port map (
            O => \N__40428\,
            I => \N__40390\
        );

    \I__9357\ : InMux
    port map (
            O => \N__40427\,
            I => \N__40390\
        );

    \I__9356\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40387\
        );

    \I__9355\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40382\
        );

    \I__9354\ : InMux
    port map (
            O => \N__40424\,
            I => \N__40382\
        );

    \I__9353\ : InMux
    port map (
            O => \N__40423\,
            I => \N__40379\
        );

    \I__9352\ : InMux
    port map (
            O => \N__40422\,
            I => \N__40374\
        );

    \I__9351\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40374\
        );

    \I__9350\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40367\
        );

    \I__9349\ : InMux
    port map (
            O => \N__40419\,
            I => \N__40367\
        );

    \I__9348\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40367\
        );

    \I__9347\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40358\
        );

    \I__9346\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40358\
        );

    \I__9345\ : InMux
    port map (
            O => \N__40411\,
            I => \N__40358\
        );

    \I__9344\ : InMux
    port map (
            O => \N__40410\,
            I => \N__40358\
        );

    \I__9343\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40349\
        );

    \I__9342\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40349\
        );

    \I__9341\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40349\
        );

    \I__9340\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40349\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__40403\,
            I => \N__40346\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__40400\,
            I => \N__40341\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__40397\,
            I => \N__40341\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__40390\,
            I => \N__40338\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__40387\,
            I => \c0.n17076\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__40382\,
            I => \c0.n17076\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__40379\,
            I => \c0.n17076\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__40374\,
            I => \c0.n17076\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__40367\,
            I => \c0.n17076\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__40358\,
            I => \c0.n17076\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__40349\,
            I => \c0.n17076\
        );

    \I__9328\ : Odrv4
    port map (
            O => \N__40346\,
            I => \c0.n17076\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__40341\,
            I => \c0.n17076\
        );

    \I__9326\ : Odrv4
    port map (
            O => \N__40338\,
            I => \c0.n17076\
        );

    \I__9325\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40310\
        );

    \I__9324\ : InMux
    port map (
            O => \N__40316\,
            I => \N__40305\
        );

    \I__9323\ : InMux
    port map (
            O => \N__40315\,
            I => \N__40305\
        );

    \I__9322\ : InMux
    port map (
            O => \N__40314\,
            I => \N__40300\
        );

    \I__9321\ : InMux
    port map (
            O => \N__40313\,
            I => \N__40300\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__40310\,
            I => \c0.n26_adj_2174\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__40305\,
            I => \c0.n26_adj_2174\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__40300\,
            I => \c0.n26_adj_2174\
        );

    \I__9317\ : CascadeMux
    port map (
            O => \N__40293\,
            I => \c0.n17487_cascade_\
        );

    \I__9316\ : InMux
    port map (
            O => \N__40290\,
            I => \N__40287\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__40287\,
            I => \N__40283\
        );

    \I__9314\ : InMux
    port map (
            O => \N__40286\,
            I => \N__40280\
        );

    \I__9313\ : Span4Mux_v
    port map (
            O => \N__40283\,
            I => \N__40277\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__40280\,
            I => \N__40274\
        );

    \I__9311\ : Span4Mux_h
    port map (
            O => \N__40277\,
            I => \N__40267\
        );

    \I__9310\ : Span4Mux_h
    port map (
            O => \N__40274\,
            I => \N__40267\
        );

    \I__9309\ : InMux
    port map (
            O => \N__40273\,
            I => \N__40264\
        );

    \I__9308\ : InMux
    port map (
            O => \N__40272\,
            I => \N__40261\
        );

    \I__9307\ : Span4Mux_h
    port map (
            O => \N__40267\,
            I => \N__40258\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__40264\,
            I => \N__40255\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__40261\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__40258\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__9303\ : Odrv12
    port map (
            O => \N__40255\,
            I => \c0.data_out_frame2_0_1\
        );

    \I__9302\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40240\
        );

    \I__9301\ : InMux
    port map (
            O => \N__40247\,
            I => \N__40236\
        );

    \I__9300\ : InMux
    port map (
            O => \N__40246\,
            I => \N__40227\
        );

    \I__9299\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40227\
        );

    \I__9298\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40227\
        );

    \I__9297\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40224\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__40240\,
            I => \N__40221\
        );

    \I__9295\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40216\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__40236\,
            I => \N__40213\
        );

    \I__9293\ : InMux
    port map (
            O => \N__40235\,
            I => \N__40208\
        );

    \I__9292\ : InMux
    port map (
            O => \N__40234\,
            I => \N__40208\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__40227\,
            I => \N__40203\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__40224\,
            I => \N__40203\
        );

    \I__9289\ : Span4Mux_h
    port map (
            O => \N__40221\,
            I => \N__40200\
        );

    \I__9288\ : CascadeMux
    port map (
            O => \N__40220\,
            I => \N__40194\
        );

    \I__9287\ : InMux
    port map (
            O => \N__40219\,
            I => \N__40189\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__40216\,
            I => \N__40186\
        );

    \I__9285\ : Span4Mux_h
    port map (
            O => \N__40213\,
            I => \N__40181\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__40208\,
            I => \N__40181\
        );

    \I__9283\ : Span4Mux_v
    port map (
            O => \N__40203\,
            I => \N__40176\
        );

    \I__9282\ : Span4Mux_h
    port map (
            O => \N__40200\,
            I => \N__40176\
        );

    \I__9281\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40171\
        );

    \I__9280\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40171\
        );

    \I__9279\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40168\
        );

    \I__9278\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40161\
        );

    \I__9277\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40161\
        );

    \I__9276\ : InMux
    port map (
            O => \N__40192\,
            I => \N__40161\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__40189\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__40186\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9273\ : Odrv4
    port map (
            O => \N__40181\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9272\ : Odrv4
    port map (
            O => \N__40176\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__40171\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__40168\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__40161\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__9268\ : CascadeMux
    port map (
            O => \N__40146\,
            I => \N__40137\
        );

    \I__9267\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40134\
        );

    \I__9266\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40129\
        );

    \I__9265\ : InMux
    port map (
            O => \N__40143\,
            I => \N__40129\
        );

    \I__9264\ : InMux
    port map (
            O => \N__40142\,
            I => \N__40126\
        );

    \I__9263\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40121\
        );

    \I__9262\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40121\
        );

    \I__9261\ : InMux
    port map (
            O => \N__40137\,
            I => \N__40118\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__40134\,
            I => \c0.n12491\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__40129\,
            I => \c0.n12491\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__40126\,
            I => \c0.n12491\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__40121\,
            I => \c0.n12491\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__40118\,
            I => \c0.n12491\
        );

    \I__9255\ : CascadeMux
    port map (
            O => \N__40107\,
            I => \c0.n17690_cascade_\
        );

    \I__9254\ : InMux
    port map (
            O => \N__40104\,
            I => \N__40100\
        );

    \I__9253\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40097\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__40097\,
            I => \N__40090\
        );

    \I__9250\ : Span4Mux_v
    port map (
            O => \N__40094\,
            I => \N__40086\
        );

    \I__9249\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40083\
        );

    \I__9248\ : Span4Mux_h
    port map (
            O => \N__40090\,
            I => \N__40080\
        );

    \I__9247\ : CascadeMux
    port map (
            O => \N__40089\,
            I => \N__40076\
        );

    \I__9246\ : Sp12to4
    port map (
            O => \N__40086\,
            I => \N__40071\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__40083\,
            I => \N__40071\
        );

    \I__9244\ : Span4Mux_h
    port map (
            O => \N__40080\,
            I => \N__40068\
        );

    \I__9243\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40063\
        );

    \I__9242\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40063\
        );

    \I__9241\ : Span12Mux_s5_h
    port map (
            O => \N__40071\,
            I => \N__40060\
        );

    \I__9240\ : Span4Mux_h
    port map (
            O => \N__40068\,
            I => \N__40057\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__40063\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__9238\ : Odrv12
    port map (
            O => \N__40060\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__40057\,
            I => \c0.data_out_frame2_0_2\
        );

    \I__9236\ : InMux
    port map (
            O => \N__40050\,
            I => \N__40046\
        );

    \I__9235\ : InMux
    port map (
            O => \N__40049\,
            I => \N__40043\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__40046\,
            I => \N__40040\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__40043\,
            I => \N__40037\
        );

    \I__9232\ : Span4Mux_h
    port map (
            O => \N__40040\,
            I => \N__40034\
        );

    \I__9231\ : Span4Mux_h
    port map (
            O => \N__40037\,
            I => \N__40031\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__40034\,
            I => \c0.data_in_frame_5_2\
        );

    \I__9229\ : Odrv4
    port map (
            O => \N__40031\,
            I => \c0.data_in_frame_5_2\
        );

    \I__9228\ : InMux
    port map (
            O => \N__40026\,
            I => \N__40023\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__40023\,
            I => \N__40016\
        );

    \I__9226\ : InMux
    port map (
            O => \N__40022\,
            I => \N__40011\
        );

    \I__9225\ : InMux
    port map (
            O => \N__40021\,
            I => \N__40011\
        );

    \I__9224\ : InMux
    port map (
            O => \N__40020\,
            I => \N__40006\
        );

    \I__9223\ : InMux
    port map (
            O => \N__40019\,
            I => \N__40006\
        );

    \I__9222\ : Odrv12
    port map (
            O => \N__40016\,
            I => \c0.data_in_frame_1_0\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__40011\,
            I => \c0.data_in_frame_1_0\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40006\,
            I => \c0.data_in_frame_1_0\
        );

    \I__9219\ : InMux
    port map (
            O => \N__39999\,
            I => \N__39995\
        );

    \I__9218\ : CascadeMux
    port map (
            O => \N__39998\,
            I => \N__39990\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__39995\,
            I => \N__39987\
        );

    \I__9216\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39984\
        );

    \I__9215\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39980\
        );

    \I__9214\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39977\
        );

    \I__9213\ : Span4Mux_h
    port map (
            O => \N__39987\,
            I => \N__39972\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__39984\,
            I => \N__39972\
        );

    \I__9211\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39969\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__39980\,
            I => \N__39966\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__39977\,
            I => \c0.data_in_frame_1_1\
        );

    \I__9208\ : Odrv4
    port map (
            O => \N__39972\,
            I => \c0.data_in_frame_1_1\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__39969\,
            I => \c0.data_in_frame_1_1\
        );

    \I__9206\ : Odrv4
    port map (
            O => \N__39966\,
            I => \c0.data_in_frame_1_1\
        );

    \I__9205\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39954\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__39954\,
            I => \c0.n17102\
        );

    \I__9203\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39948\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__39948\,
            I => \N__39940\
        );

    \I__9201\ : InMux
    port map (
            O => \N__39947\,
            I => \N__39937\
        );

    \I__9200\ : InMux
    port map (
            O => \N__39946\,
            I => \N__39929\
        );

    \I__9199\ : InMux
    port map (
            O => \N__39945\,
            I => \N__39929\
        );

    \I__9198\ : InMux
    port map (
            O => \N__39944\,
            I => \N__39924\
        );

    \I__9197\ : InMux
    port map (
            O => \N__39943\,
            I => \N__39924\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__39940\,
            I => \N__39921\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__39937\,
            I => \N__39918\
        );

    \I__9194\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39915\
        );

    \I__9193\ : InMux
    port map (
            O => \N__39935\,
            I => \N__39910\
        );

    \I__9192\ : InMux
    port map (
            O => \N__39934\,
            I => \N__39910\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39905\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__39924\,
            I => \N__39905\
        );

    \I__9189\ : Sp12to4
    port map (
            O => \N__39921\,
            I => \N__39902\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__39918\,
            I => \N__39899\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__39915\,
            I => \N__39896\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__39910\,
            I => \N__39893\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__39905\,
            I => \N__39890\
        );

    \I__9184\ : Odrv12
    port map (
            O => \N__39902\,
            I => \c0.n5815\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__39899\,
            I => \c0.n5815\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__39896\,
            I => \c0.n5815\
        );

    \I__9181\ : Odrv4
    port map (
            O => \N__39893\,
            I => \c0.n5815\
        );

    \I__9180\ : Odrv4
    port map (
            O => \N__39890\,
            I => \c0.n5815\
        );

    \I__9179\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39871\
        );

    \I__9178\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39866\
        );

    \I__9177\ : InMux
    port map (
            O => \N__39877\,
            I => \N__39866\
        );

    \I__9176\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39863\
        );

    \I__9175\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39860\
        );

    \I__9174\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39857\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__39871\,
            I => \c0.n4494\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__39866\,
            I => \c0.n4494\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__39863\,
            I => \c0.n4494\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__39860\,
            I => \c0.n4494\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__39857\,
            I => \c0.n4494\
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__39846\,
            I => \N__39841\
        );

    \I__9167\ : CascadeMux
    port map (
            O => \N__39845\,
            I => \N__39838\
        );

    \I__9166\ : CascadeMux
    port map (
            O => \N__39844\,
            I => \N__39832\
        );

    \I__9165\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39828\
        );

    \I__9164\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39821\
        );

    \I__9163\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39818\
        );

    \I__9162\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39815\
        );

    \I__9161\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39812\
        );

    \I__9160\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39807\
        );

    \I__9159\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39807\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__39828\,
            I => \N__39804\
        );

    \I__9157\ : InMux
    port map (
            O => \N__39827\,
            I => \N__39795\
        );

    \I__9156\ : InMux
    port map (
            O => \N__39826\,
            I => \N__39795\
        );

    \I__9155\ : InMux
    port map (
            O => \N__39825\,
            I => \N__39795\
        );

    \I__9154\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39795\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__39821\,
            I => \N__39792\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__39818\,
            I => \N__39789\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39782\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__39812\,
            I => \N__39782\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__39807\,
            I => \N__39782\
        );

    \I__9148\ : Span4Mux_h
    port map (
            O => \N__39804\,
            I => \N__39779\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__39795\,
            I => \N__39776\
        );

    \I__9146\ : Span4Mux_h
    port map (
            O => \N__39792\,
            I => \N__39773\
        );

    \I__9145\ : Span4Mux_v
    port map (
            O => \N__39789\,
            I => \N__39768\
        );

    \I__9144\ : Span4Mux_v
    port map (
            O => \N__39782\,
            I => \N__39768\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__39779\,
            I => \c0.n5817\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__39776\,
            I => \c0.n5817\
        );

    \I__9141\ : Odrv4
    port map (
            O => \N__39773\,
            I => \c0.n5817\
        );

    \I__9140\ : Odrv4
    port map (
            O => \N__39768\,
            I => \c0.n5817\
        );

    \I__9139\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39755\
        );

    \I__9138\ : InMux
    port map (
            O => \N__39758\,
            I => \N__39750\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__39755\,
            I => \N__39747\
        );

    \I__9136\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39742\
        );

    \I__9135\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39742\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__39750\,
            I => \N__39739\
        );

    \I__9133\ : Span12Mux_h
    port map (
            O => \N__39747\,
            I => \N__39734\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__39742\,
            I => \N__39734\
        );

    \I__9131\ : Odrv12
    port map (
            O => \N__39739\,
            I => n31_adj_2415
        );

    \I__9130\ : Odrv12
    port map (
            O => \N__39734\,
            I => n31_adj_2415
        );

    \I__9129\ : CascadeMux
    port map (
            O => \N__39729\,
            I => \N__39726\
        );

    \I__9128\ : InMux
    port map (
            O => \N__39726\,
            I => \N__39719\
        );

    \I__9127\ : InMux
    port map (
            O => \N__39725\,
            I => \N__39719\
        );

    \I__9126\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39716\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__39719\,
            I => \c0.n18202\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__39716\,
            I => \c0.n18202\
        );

    \I__9123\ : InMux
    port map (
            O => \N__39711\,
            I => \N__39708\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__39708\,
            I => \N__39705\
        );

    \I__9121\ : Odrv12
    port map (
            O => \N__39705\,
            I => \c0.n17712\
        );

    \I__9120\ : InMux
    port map (
            O => \N__39702\,
            I => \N__39698\
        );

    \I__9119\ : CascadeMux
    port map (
            O => \N__39701\,
            I => \N__39694\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39690\
        );

    \I__9117\ : CascadeMux
    port map (
            O => \N__39697\,
            I => \N__39687\
        );

    \I__9116\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39684\
        );

    \I__9115\ : CascadeMux
    port map (
            O => \N__39693\,
            I => \N__39680\
        );

    \I__9114\ : Sp12to4
    port map (
            O => \N__39690\,
            I => \N__39675\
        );

    \I__9113\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39672\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__39684\,
            I => \N__39669\
        );

    \I__9111\ : CascadeMux
    port map (
            O => \N__39683\,
            I => \N__39666\
        );

    \I__9110\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39663\
        );

    \I__9109\ : CascadeMux
    port map (
            O => \N__39679\,
            I => \N__39660\
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__39678\,
            I => \N__39657\
        );

    \I__9107\ : Span12Mux_v
    port map (
            O => \N__39675\,
            I => \N__39652\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__39672\,
            I => \N__39652\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__39669\,
            I => \N__39649\
        );

    \I__9104\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39646\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__39663\,
            I => \N__39643\
        );

    \I__9102\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39640\
        );

    \I__9101\ : InMux
    port map (
            O => \N__39657\,
            I => \N__39637\
        );

    \I__9100\ : Odrv12
    port map (
            O => \N__39652\,
            I => \c0.n11867\
        );

    \I__9099\ : Odrv4
    port map (
            O => \N__39649\,
            I => \c0.n11867\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__39646\,
            I => \c0.n11867\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__39643\,
            I => \c0.n11867\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__39640\,
            I => \c0.n11867\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__39637\,
            I => \c0.n11867\
        );

    \I__9094\ : InMux
    port map (
            O => \N__39624\,
            I => \N__39619\
        );

    \I__9093\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39616\
        );

    \I__9092\ : CascadeMux
    port map (
            O => \N__39622\,
            I => \N__39613\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__39619\,
            I => \N__39609\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__39616\,
            I => \N__39606\
        );

    \I__9089\ : InMux
    port map (
            O => \N__39613\,
            I => \N__39603\
        );

    \I__9088\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39600\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__39609\,
            I => \N__39593\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__39606\,
            I => \N__39593\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__39603\,
            I => \N__39593\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__39600\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__9083\ : Odrv4
    port map (
            O => \N__39593\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__9082\ : SRMux
    port map (
            O => \N__39588\,
            I => \N__39585\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__9080\ : Span4Mux_h
    port map (
            O => \N__39582\,
            I => \N__39579\
        );

    \I__9079\ : Odrv4
    port map (
            O => \N__39579\,
            I => \c0.n4_adj_2147\
        );

    \I__9078\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39573\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__39573\,
            I => \N__39569\
        );

    \I__9076\ : InMux
    port map (
            O => \N__39572\,
            I => \N__39566\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__39569\,
            I => \N__39563\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__39566\,
            I => \N__39560\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__39563\,
            I => n13116
        );

    \I__9072\ : Odrv12
    port map (
            O => \N__39560\,
            I => n13116
        );

    \I__9071\ : CascadeMux
    port map (
            O => \N__39555\,
            I => \N__39549\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__39554\,
            I => \N__39546\
        );

    \I__9069\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39542\
        );

    \I__9068\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39538\
        );

    \I__9067\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39535\
        );

    \I__9066\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39530\
        );

    \I__9065\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39530\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__39542\,
            I => \N__39527\
        );

    \I__9063\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39524\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__39538\,
            I => \N__39520\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__39535\,
            I => \N__39516\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__39530\,
            I => \N__39511\
        );

    \I__9059\ : Span4Mux_v
    port map (
            O => \N__39527\,
            I => \N__39511\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__39524\,
            I => \N__39508\
        );

    \I__9057\ : CascadeMux
    port map (
            O => \N__39523\,
            I => \N__39505\
        );

    \I__9056\ : Span4Mux_h
    port map (
            O => \N__39520\,
            I => \N__39502\
        );

    \I__9055\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39499\
        );

    \I__9054\ : Span4Mux_v
    port map (
            O => \N__39516\,
            I => \N__39492\
        );

    \I__9053\ : Span4Mux_h
    port map (
            O => \N__39511\,
            I => \N__39492\
        );

    \I__9052\ : Span4Mux_v
    port map (
            O => \N__39508\,
            I => \N__39492\
        );

    \I__9051\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39489\
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__39502\,
            I => rx_data_6
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__39499\,
            I => rx_data_6
        );

    \I__9048\ : Odrv4
    port map (
            O => \N__39492\,
            I => rx_data_6
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__39489\,
            I => rx_data_6
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__39480\,
            I => \N__39473\
        );

    \I__9045\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39470\
        );

    \I__9044\ : CascadeMux
    port map (
            O => \N__39478\,
            I => \N__39466\
        );

    \I__9043\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39463\
        );

    \I__9042\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39459\
        );

    \I__9041\ : InMux
    port map (
            O => \N__39473\,
            I => \N__39456\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__39470\,
            I => \N__39453\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__39469\,
            I => \N__39450\
        );

    \I__9038\ : InMux
    port map (
            O => \N__39466\,
            I => \N__39447\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__39463\,
            I => \N__39443\
        );

    \I__9036\ : CascadeMux
    port map (
            O => \N__39462\,
            I => \N__39440\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__39459\,
            I => \N__39433\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__39456\,
            I => \N__39433\
        );

    \I__9033\ : Span4Mux_h
    port map (
            O => \N__39453\,
            I => \N__39433\
        );

    \I__9032\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39430\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__39447\,
            I => \N__39427\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__39446\,
            I => \N__39424\
        );

    \I__9029\ : Span4Mux_h
    port map (
            O => \N__39443\,
            I => \N__39421\
        );

    \I__9028\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39418\
        );

    \I__9027\ : Span4Mux_h
    port map (
            O => \N__39433\,
            I => \N__39415\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__39430\,
            I => \N__39410\
        );

    \I__9025\ : Span4Mux_v
    port map (
            O => \N__39427\,
            I => \N__39410\
        );

    \I__9024\ : InMux
    port map (
            O => \N__39424\,
            I => \N__39407\
        );

    \I__9023\ : Odrv4
    port map (
            O => \N__39421\,
            I => rx_data_1
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__39418\,
            I => rx_data_1
        );

    \I__9021\ : Odrv4
    port map (
            O => \N__39415\,
            I => rx_data_1
        );

    \I__9020\ : Odrv4
    port map (
            O => \N__39410\,
            I => rx_data_1
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__39407\,
            I => rx_data_1
        );

    \I__9018\ : CascadeMux
    port map (
            O => \N__39396\,
            I => \N__39391\
        );

    \I__9017\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39382\
        );

    \I__9016\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39379\
        );

    \I__9015\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39376\
        );

    \I__9014\ : InMux
    port map (
            O => \N__39390\,
            I => \N__39373\
        );

    \I__9013\ : InMux
    port map (
            O => \N__39389\,
            I => \N__39363\
        );

    \I__9012\ : InMux
    port map (
            O => \N__39388\,
            I => \N__39363\
        );

    \I__9011\ : InMux
    port map (
            O => \N__39387\,
            I => \N__39363\
        );

    \I__9010\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39354\
        );

    \I__9009\ : InMux
    port map (
            O => \N__39385\,
            I => \N__39354\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__39382\,
            I => \N__39351\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__39379\,
            I => \N__39348\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__39376\,
            I => \N__39343\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__39373\,
            I => \N__39343\
        );

    \I__9004\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39336\
        );

    \I__9003\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39336\
        );

    \I__9002\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39336\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__39363\,
            I => \N__39333\
        );

    \I__9000\ : InMux
    port map (
            O => \N__39362\,
            I => \N__39330\
        );

    \I__8999\ : InMux
    port map (
            O => \N__39361\,
            I => \N__39327\
        );

    \I__8998\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39324\
        );

    \I__8997\ : InMux
    port map (
            O => \N__39359\,
            I => \N__39321\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__39354\,
            I => \N__39318\
        );

    \I__8995\ : Span4Mux_h
    port map (
            O => \N__39351\,
            I => \N__39311\
        );

    \I__8994\ : Span4Mux_h
    port map (
            O => \N__39348\,
            I => \N__39311\
        );

    \I__8993\ : Span4Mux_v
    port map (
            O => \N__39343\,
            I => \N__39311\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__39336\,
            I => \N__39306\
        );

    \I__8991\ : Span4Mux_v
    port map (
            O => \N__39333\,
            I => \N__39306\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__39330\,
            I => \N__39303\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__39327\,
            I => \c0.n17072\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__39324\,
            I => \c0.n17072\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__39321\,
            I => \c0.n17072\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__39318\,
            I => \c0.n17072\
        );

    \I__8985\ : Odrv4
    port map (
            O => \N__39311\,
            I => \c0.n17072\
        );

    \I__8984\ : Odrv4
    port map (
            O => \N__39306\,
            I => \c0.n17072\
        );

    \I__8983\ : Odrv4
    port map (
            O => \N__39303\,
            I => \c0.n17072\
        );

    \I__8982\ : CascadeMux
    port map (
            O => \N__39288\,
            I => \N__39285\
        );

    \I__8981\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39282\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__39282\,
            I => \N__39278\
        );

    \I__8979\ : InMux
    port map (
            O => \N__39281\,
            I => \N__39275\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__39278\,
            I => \N__39272\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__39275\,
            I => \c0.data_in_frame_3_1\
        );

    \I__8976\ : Odrv4
    port map (
            O => \N__39272\,
            I => \c0.data_in_frame_3_1\
        );

    \I__8975\ : CascadeMux
    port map (
            O => \N__39267\,
            I => \c0.n17472_cascade_\
        );

    \I__8974\ : InMux
    port map (
            O => \N__39264\,
            I => \N__39260\
        );

    \I__8973\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39255\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__39260\,
            I => \N__39252\
        );

    \I__8971\ : InMux
    port map (
            O => \N__39259\,
            I => \N__39249\
        );

    \I__8970\ : CascadeMux
    port map (
            O => \N__39258\,
            I => \N__39246\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__39255\,
            I => \N__39243\
        );

    \I__8968\ : Span4Mux_v
    port map (
            O => \N__39252\,
            I => \N__39238\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__39249\,
            I => \N__39238\
        );

    \I__8966\ : InMux
    port map (
            O => \N__39246\,
            I => \N__39235\
        );

    \I__8965\ : Span4Mux_v
    port map (
            O => \N__39243\,
            I => \N__39232\
        );

    \I__8964\ : Span4Mux_h
    port map (
            O => \N__39238\,
            I => \N__39229\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__39235\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__39232\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__39229\,
            I => \c0.data_out_frame2_0_6\
        );

    \I__8960\ : InMux
    port map (
            O => \N__39222\,
            I => \N__39201\
        );

    \I__8959\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39195\
        );

    \I__8958\ : InMux
    port map (
            O => \N__39220\,
            I => \N__39195\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__39219\,
            I => \N__39191\
        );

    \I__8956\ : CascadeMux
    port map (
            O => \N__39218\,
            I => \N__39187\
        );

    \I__8955\ : InMux
    port map (
            O => \N__39217\,
            I => \N__39179\
        );

    \I__8954\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39179\
        );

    \I__8953\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39174\
        );

    \I__8952\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39174\
        );

    \I__8951\ : InMux
    port map (
            O => \N__39213\,
            I => \N__39163\
        );

    \I__8950\ : InMux
    port map (
            O => \N__39212\,
            I => \N__39163\
        );

    \I__8949\ : InMux
    port map (
            O => \N__39211\,
            I => \N__39163\
        );

    \I__8948\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39163\
        );

    \I__8947\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39163\
        );

    \I__8946\ : InMux
    port map (
            O => \N__39208\,
            I => \N__39160\
        );

    \I__8945\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39157\
        );

    \I__8944\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39154\
        );

    \I__8943\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39149\
        );

    \I__8942\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39149\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__39201\,
            I => \N__39146\
        );

    \I__8940\ : InMux
    port map (
            O => \N__39200\,
            I => \N__39143\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39139\
        );

    \I__8938\ : InMux
    port map (
            O => \N__39194\,
            I => \N__39136\
        );

    \I__8937\ : InMux
    port map (
            O => \N__39191\,
            I => \N__39133\
        );

    \I__8936\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39126\
        );

    \I__8935\ : InMux
    port map (
            O => \N__39187\,
            I => \N__39119\
        );

    \I__8934\ : InMux
    port map (
            O => \N__39186\,
            I => \N__39119\
        );

    \I__8933\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39119\
        );

    \I__8932\ : InMux
    port map (
            O => \N__39184\,
            I => \N__39116\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__39179\,
            I => \N__39103\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__39174\,
            I => \N__39103\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__39163\,
            I => \N__39103\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39103\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__39157\,
            I => \N__39103\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__39154\,
            I => \N__39103\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__39149\,
            I => \N__39096\
        );

    \I__8924\ : Span4Mux_v
    port map (
            O => \N__39146\,
            I => \N__39096\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__39143\,
            I => \N__39096\
        );

    \I__8922\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39090\
        );

    \I__8921\ : Span4Mux_v
    port map (
            O => \N__39139\,
            I => \N__39087\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__39136\,
            I => \N__39082\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__39133\,
            I => \N__39082\
        );

    \I__8918\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39079\
        );

    \I__8917\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39072\
        );

    \I__8916\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39072\
        );

    \I__8915\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39072\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__39126\,
            I => \N__39067\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__39119\,
            I => \N__39067\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__39116\,
            I => \N__39060\
        );

    \I__8911\ : Span4Mux_v
    port map (
            O => \N__39103\,
            I => \N__39060\
        );

    \I__8910\ : Span4Mux_h
    port map (
            O => \N__39096\,
            I => \N__39060\
        );

    \I__8909\ : InMux
    port map (
            O => \N__39095\,
            I => \N__39056\
        );

    \I__8908\ : InMux
    port map (
            O => \N__39094\,
            I => \N__39051\
        );

    \I__8907\ : InMux
    port map (
            O => \N__39093\,
            I => \N__39051\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__39090\,
            I => \N__39044\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__39087\,
            I => \N__39044\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__39082\,
            I => \N__39044\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N__39037\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__39072\,
            I => \N__39037\
        );

    \I__8901\ : Span4Mux_v
    port map (
            O => \N__39067\,
            I => \N__39037\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__39060\,
            I => \N__39034\
        );

    \I__8899\ : CascadeMux
    port map (
            O => \N__39059\,
            I => \N__39031\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__39056\,
            I => \N__39025\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__39051\,
            I => \N__39025\
        );

    \I__8896\ : Sp12to4
    port map (
            O => \N__39044\,
            I => \N__39022\
        );

    \I__8895\ : Span4Mux_h
    port map (
            O => \N__39037\,
            I => \N__39017\
        );

    \I__8894\ : Span4Mux_v
    port map (
            O => \N__39034\,
            I => \N__39017\
        );

    \I__8893\ : InMux
    port map (
            O => \N__39031\,
            I => \N__39013\
        );

    \I__8892\ : InMux
    port map (
            O => \N__39030\,
            I => \N__39010\
        );

    \I__8891\ : Span12Mux_h
    port map (
            O => \N__39025\,
            I => \N__39007\
        );

    \I__8890\ : Span12Mux_v
    port map (
            O => \N__39022\,
            I => \N__39004\
        );

    \I__8889\ : Span4Mux_v
    port map (
            O => \N__39017\,
            I => \N__39001\
        );

    \I__8888\ : InMux
    port map (
            O => \N__39016\,
            I => \N__38998\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__39013\,
            I => rx_data_ready
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__39010\,
            I => rx_data_ready
        );

    \I__8885\ : Odrv12
    port map (
            O => \N__39007\,
            I => rx_data_ready
        );

    \I__8884\ : Odrv12
    port map (
            O => \N__39004\,
            I => rx_data_ready
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__39001\,
            I => rx_data_ready
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__38998\,
            I => rx_data_ready
        );

    \I__8881\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__38982\,
            I => \N__38979\
        );

    \I__8879\ : Span4Mux_v
    port map (
            O => \N__38979\,
            I => \N__38974\
        );

    \I__8878\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38971\
        );

    \I__8877\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38968\
        );

    \I__8876\ : Span4Mux_h
    port map (
            O => \N__38974\,
            I => \N__38964\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__38971\,
            I => \N__38961\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__38968\,
            I => \N__38958\
        );

    \I__8873\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38955\
        );

    \I__8872\ : Span4Mux_h
    port map (
            O => \N__38964\,
            I => \N__38950\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__38961\,
            I => \N__38950\
        );

    \I__8870\ : Sp12to4
    port map (
            O => \N__38958\,
            I => \N__38947\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__38955\,
            I => data_in_3_2
        );

    \I__8868\ : Odrv4
    port map (
            O => \N__38950\,
            I => data_in_3_2
        );

    \I__8867\ : Odrv12
    port map (
            O => \N__38947\,
            I => data_in_3_2
        );

    \I__8866\ : InMux
    port map (
            O => \N__38940\,
            I => \N__38936\
        );

    \I__8865\ : InMux
    port map (
            O => \N__38939\,
            I => \N__38933\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__38936\,
            I => \N__38929\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__38933\,
            I => \N__38926\
        );

    \I__8862\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38923\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__38929\,
            I => \N__38919\
        );

    \I__8860\ : Span4Mux_v
    port map (
            O => \N__38926\,
            I => \N__38914\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__38923\,
            I => \N__38914\
        );

    \I__8858\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38911\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__38919\,
            I => \N__38906\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__38914\,
            I => \N__38906\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__38911\,
            I => data_in_2_2
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__38906\,
            I => data_in_2_2
        );

    \I__8853\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38896\
        );

    \I__8852\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38893\
        );

    \I__8851\ : CascadeMux
    port map (
            O => \N__38899\,
            I => \N__38889\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__38896\,
            I => \N__38886\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__38893\,
            I => \N__38882\
        );

    \I__8848\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38879\
        );

    \I__8847\ : InMux
    port map (
            O => \N__38889\,
            I => \N__38876\
        );

    \I__8846\ : Span4Mux_v
    port map (
            O => \N__38886\,
            I => \N__38873\
        );

    \I__8845\ : InMux
    port map (
            O => \N__38885\,
            I => \N__38870\
        );

    \I__8844\ : Span4Mux_v
    port map (
            O => \N__38882\,
            I => \N__38867\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__38879\,
            I => \N__38864\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__38876\,
            I => \c0.data_in_frame_1_3\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__38873\,
            I => \c0.data_in_frame_1_3\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__38870\,
            I => \c0.data_in_frame_1_3\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__38867\,
            I => \c0.data_in_frame_1_3\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__38864\,
            I => \c0.data_in_frame_1_3\
        );

    \I__8837\ : CascadeMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__8836\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38846\
        );

    \I__8835\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38843\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__38846\,
            I => \N__38840\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__38843\,
            I => \N__38835\
        );

    \I__8832\ : Span4Mux_v
    port map (
            O => \N__38840\,
            I => \N__38835\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__38835\,
            I => \c0.data_in_frame_5_4\
        );

    \I__8830\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38829\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__38829\,
            I => \N__38824\
        );

    \I__8828\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38819\
        );

    \I__8827\ : InMux
    port map (
            O => \N__38827\,
            I => \N__38816\
        );

    \I__8826\ : Span4Mux_h
    port map (
            O => \N__38824\,
            I => \N__38813\
        );

    \I__8825\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38808\
        );

    \I__8824\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38808\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__38819\,
            I => \N__38803\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__38816\,
            I => \N__38803\
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__38813\,
            I => \c0.data_in_frame_1_2\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__38808\,
            I => \c0.data_in_frame_1_2\
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__38803\,
            I => \c0.data_in_frame_1_2\
        );

    \I__8818\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38793\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__38793\,
            I => \c0.n21_adj_2357\
        );

    \I__8816\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38786\
        );

    \I__8815\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38783\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__38786\,
            I => \c0.delay_counter_12\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__38783\,
            I => \c0.delay_counter_12\
        );

    \I__8812\ : InMux
    port map (
            O => \N__38778\,
            I => \N__38775\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__38775\,
            I => \c0.n16_adj_2212\
        );

    \I__8810\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38766\
        );

    \I__8809\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38766\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__38766\,
            I => \c0.delay_counter_2\
        );

    \I__8807\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38760\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__38760\,
            I => \c0.n26\
        );

    \I__8805\ : InMux
    port map (
            O => \N__38757\,
            I => \N__38753\
        );

    \I__8804\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38750\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__38753\,
            I => \c0.delay_counter_0\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__38750\,
            I => \c0.delay_counter_0\
        );

    \I__8801\ : InMux
    port map (
            O => \N__38745\,
            I => \N__38741\
        );

    \I__8800\ : InMux
    port map (
            O => \N__38744\,
            I => \N__38738\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__38741\,
            I => \c0.delay_counter_6\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__38738\,
            I => \c0.delay_counter_6\
        );

    \I__8797\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__38730\,
            I => \c0.n22_adj_2390\
        );

    \I__8795\ : InMux
    port map (
            O => \N__38727\,
            I => \N__38721\
        );

    \I__8794\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38721\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__38721\,
            I => \c0.delay_counter_10\
        );

    \I__8792\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38715\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__38715\,
            I => \c0.n18_adj_2220\
        );

    \I__8790\ : CascadeMux
    port map (
            O => \N__38712\,
            I => \N__38708\
        );

    \I__8789\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38703\
        );

    \I__8788\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38703\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__38703\,
            I => \c0.delay_counter_13\
        );

    \I__8786\ : InMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__38697\,
            I => \c0.n15_adj_2211\
        );

    \I__8784\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__38691\,
            I => \N__38687\
        );

    \I__8782\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38684\
        );

    \I__8781\ : Span4Mux_h
    port map (
            O => \N__38687\,
            I => \N__38681\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__38684\,
            I => \r_Tx_Data_5\
        );

    \I__8779\ : Odrv4
    port map (
            O => \N__38681\,
            I => \r_Tx_Data_5\
        );

    \I__8778\ : InMux
    port map (
            O => \N__38676\,
            I => \N__38672\
        );

    \I__8777\ : InMux
    port map (
            O => \N__38675\,
            I => \N__38669\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__38672\,
            I => \c0.delay_counter_11\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__38669\,
            I => \c0.delay_counter_11\
        );

    \I__8774\ : InMux
    port map (
            O => \N__38664\,
            I => \N__38657\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__38663\,
            I => \N__38654\
        );

    \I__8772\ : InMux
    port map (
            O => \N__38662\,
            I => \N__38649\
        );

    \I__8771\ : CascadeMux
    port map (
            O => \N__38661\,
            I => \N__38643\
        );

    \I__8770\ : CascadeMux
    port map (
            O => \N__38660\,
            I => \N__38640\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__38657\,
            I => \N__38632\
        );

    \I__8768\ : InMux
    port map (
            O => \N__38654\,
            I => \N__38625\
        );

    \I__8767\ : InMux
    port map (
            O => \N__38653\,
            I => \N__38625\
        );

    \I__8766\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38625\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__38649\,
            I => \N__38622\
        );

    \I__8764\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38615\
        );

    \I__8763\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38615\
        );

    \I__8762\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38615\
        );

    \I__8761\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38608\
        );

    \I__8760\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38608\
        );

    \I__8759\ : InMux
    port map (
            O => \N__38639\,
            I => \N__38608\
        );

    \I__8758\ : InMux
    port map (
            O => \N__38638\,
            I => \N__38605\
        );

    \I__8757\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38598\
        );

    \I__8756\ : InMux
    port map (
            O => \N__38636\,
            I => \N__38598\
        );

    \I__8755\ : InMux
    port map (
            O => \N__38635\,
            I => \N__38598\
        );

    \I__8754\ : Span4Mux_h
    port map (
            O => \N__38632\,
            I => \N__38595\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__38625\,
            I => \c0.n9453\
        );

    \I__8752\ : Odrv4
    port map (
            O => \N__38622\,
            I => \c0.n9453\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__38615\,
            I => \c0.n9453\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__38608\,
            I => \c0.n9453\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__38605\,
            I => \c0.n9453\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__38598\,
            I => \c0.n9453\
        );

    \I__8747\ : Odrv4
    port map (
            O => \N__38595\,
            I => \c0.n9453\
        );

    \I__8746\ : InMux
    port map (
            O => \N__38580\,
            I => \N__38571\
        );

    \I__8745\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38571\
        );

    \I__8744\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38571\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38555\
        );

    \I__8742\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38552\
        );

    \I__8741\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38543\
        );

    \I__8740\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38543\
        );

    \I__8739\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38543\
        );

    \I__8738\ : InMux
    port map (
            O => \N__38566\,
            I => \N__38543\
        );

    \I__8737\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38534\
        );

    \I__8736\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38534\
        );

    \I__8735\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38534\
        );

    \I__8734\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38534\
        );

    \I__8733\ : InMux
    port map (
            O => \N__38561\,
            I => \N__38527\
        );

    \I__8732\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38527\
        );

    \I__8731\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38527\
        );

    \I__8730\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38524\
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__38555\,
            I => \c0.n16267\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__38552\,
            I => \c0.n16267\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__38543\,
            I => \c0.n16267\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__38534\,
            I => \c0.n16267\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__38527\,
            I => \c0.n16267\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__38524\,
            I => \c0.n16267\
        );

    \I__8723\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38508\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__38508\,
            I => \c0.n17_adj_2219\
        );

    \I__8721\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38501\
        );

    \I__8720\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38498\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__38501\,
            I => \c0.delay_counter_8\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__38498\,
            I => \c0.delay_counter_8\
        );

    \I__8717\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38489\
        );

    \I__8716\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38486\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__38489\,
            I => \c0.delay_counter_3\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__38486\,
            I => \c0.delay_counter_3\
        );

    \I__8713\ : InMux
    port map (
            O => \N__38481\,
            I => \N__38478\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__38478\,
            I => \c0.n18_adj_2388\
        );

    \I__8711\ : InMux
    port map (
            O => \N__38475\,
            I => \N__38472\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__38472\,
            I => n17765
        );

    \I__8709\ : CascadeMux
    port map (
            O => \N__38469\,
            I => \n17392_cascade_\
        );

    \I__8708\ : InMux
    port map (
            O => \N__38466\,
            I => \N__38463\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__38463\,
            I => n17416
        );

    \I__8706\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38457\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__38457\,
            I => \c0.n20_adj_2255\
        );

    \I__8704\ : InMux
    port map (
            O => \N__38454\,
            I => \N__38450\
        );

    \I__8703\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38447\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__38450\,
            I => \c0.delay_counter_7\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__38447\,
            I => \c0.delay_counter_7\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__38442\,
            I => \N__38439\
        );

    \I__8699\ : InMux
    port map (
            O => \N__38439\,
            I => \N__38435\
        );

    \I__8698\ : InMux
    port map (
            O => \N__38438\,
            I => \N__38432\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__38435\,
            I => \c0.delay_counter_5\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__38432\,
            I => \c0.delay_counter_5\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__38427\,
            I => \c0.n24_adj_2389_cascade_\
        );

    \I__8694\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__38421\,
            I => \N__38418\
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__38418\,
            I => n17327
        );

    \I__8691\ : CascadeMux
    port map (
            O => \N__38415\,
            I => \N__38411\
        );

    \I__8690\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38408\
        );

    \I__8689\ : InMux
    port map (
            O => \N__38411\,
            I => \N__38405\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__38408\,
            I => \N__38402\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__38405\,
            I => \c0.delay_counter_1\
        );

    \I__8686\ : Odrv4
    port map (
            O => \N__38402\,
            I => \c0.delay_counter_1\
        );

    \I__8685\ : CascadeMux
    port map (
            O => \N__38397\,
            I => \N__38394\
        );

    \I__8684\ : InMux
    port map (
            O => \N__38394\,
            I => \N__38390\
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__38393\,
            I => \N__38387\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__38390\,
            I => \N__38384\
        );

    \I__8681\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38381\
        );

    \I__8680\ : Odrv4
    port map (
            O => \N__38384\,
            I => \c0.delay_counter_9\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__38381\,
            I => \c0.delay_counter_9\
        );

    \I__8678\ : InMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__38373\,
            I => \c0.n26_adj_2391\
        );

    \I__8676\ : CascadeMux
    port map (
            O => \N__38370\,
            I => \N__38366\
        );

    \I__8675\ : InMux
    port map (
            O => \N__38369\,
            I => \N__38361\
        );

    \I__8674\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38361\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__38361\,
            I => \c0.delay_counter_4\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__38358\,
            I => \c0.n9453_cascade_\
        );

    \I__8671\ : InMux
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__38352\,
            I => \c0.n24_adj_2342\
        );

    \I__8669\ : InMux
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__38346\,
            I => \c0.n453\
        );

    \I__8667\ : InMux
    port map (
            O => \N__38343\,
            I => \N__38337\
        );

    \I__8666\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38332\
        );

    \I__8665\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38332\
        );

    \I__8664\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38329\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__38337\,
            I => n4_adj_2414
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__38332\,
            I => n4_adj_2414
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__38329\,
            I => n4_adj_2414
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__38322\,
            I => \N__38319\
        );

    \I__8659\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38316\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38313\
        );

    \I__8657\ : Odrv4
    port map (
            O => \N__38313\,
            I => \c0.n19\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__38310\,
            I => \n9524_cascade_\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__38307\,
            I => \c0.n16267_cascade_\
        );

    \I__8654\ : InMux
    port map (
            O => \N__38304\,
            I => \N__38301\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__38301\,
            I => \c0.n445\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__38298\,
            I => \N__38295\
        );

    \I__8651\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38292\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__38292\,
            I => \c0.n23_adj_2314\
        );

    \I__8649\ : CascadeMux
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__8648\ : InMux
    port map (
            O => \N__38286\,
            I => \N__38283\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__38283\,
            I => \c0.n28\
        );

    \I__8646\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38277\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__38277\,
            I => n5_adj_2407
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__38274\,
            I => \N__38271\
        );

    \I__8643\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__38268\,
            I => \c0.n5_adj_2141\
        );

    \I__8641\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38261\
        );

    \I__8640\ : InMux
    port map (
            O => \N__38264\,
            I => \N__38258\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__38261\,
            I => \r_Tx_Data_2\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__38258\,
            I => \r_Tx_Data_2\
        );

    \I__8637\ : InMux
    port map (
            O => \N__38253\,
            I => \N__38250\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__38250\,
            I => \N__38246\
        );

    \I__8635\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38243\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__38246\,
            I => \N__38240\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__38243\,
            I => \r_Tx_Data_4\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__38240\,
            I => \r_Tx_Data_4\
        );

    \I__8631\ : CascadeMux
    port map (
            O => \N__38235\,
            I => \n18196_cascade_\
        );

    \I__8630\ : InMux
    port map (
            O => \N__38232\,
            I => \N__38229\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__38229\,
            I => n18199
        );

    \I__8628\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__38223\,
            I => \c0.tx.n31\
        );

    \I__8626\ : InMux
    port map (
            O => \N__38220\,
            I => \N__38217\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__38217\,
            I => n17759
        );

    \I__8624\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38211\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__38211\,
            I => \N__38208\
        );

    \I__8622\ : Odrv4
    port map (
            O => \N__38208\,
            I => n17664
        );

    \I__8621\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38202\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__38202\,
            I => \N__38199\
        );

    \I__8619\ : Odrv4
    port map (
            O => \N__38199\,
            I => \c0.n18166\
        );

    \I__8618\ : InMux
    port map (
            O => \N__38196\,
            I => \N__38193\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__38193\,
            I => \N__38190\
        );

    \I__8616\ : Span4Mux_v
    port map (
            O => \N__38190\,
            I => \N__38187\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__38187\,
            I => \c0.n2_adj_2145\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__38184\,
            I => \N__38181\
        );

    \I__8613\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38178\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__38178\,
            I => \N__38175\
        );

    \I__8611\ : Span4Mux_v
    port map (
            O => \N__38175\,
            I => \N__38172\
        );

    \I__8610\ : Span4Mux_h
    port map (
            O => \N__38172\,
            I => \N__38169\
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__38169\,
            I => \c0.n17701\
        );

    \I__8608\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38163\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__38163\,
            I => \N__38160\
        );

    \I__8606\ : Odrv4
    port map (
            O => \N__38160\,
            I => n18169
        );

    \I__8605\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__38154\,
            I => \N__38150\
        );

    \I__8603\ : CascadeMux
    port map (
            O => \N__38153\,
            I => \N__38147\
        );

    \I__8602\ : Span4Mux_v
    port map (
            O => \N__38150\,
            I => \N__38144\
        );

    \I__8601\ : InMux
    port map (
            O => \N__38147\,
            I => \N__38141\
        );

    \I__8600\ : Odrv4
    port map (
            O => \N__38144\,
            I => rand_setpoint_7
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__38141\,
            I => rand_setpoint_7
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__38136\,
            I => \N__38132\
        );

    \I__8597\ : InMux
    port map (
            O => \N__38135\,
            I => \N__38127\
        );

    \I__8596\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38127\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__38127\,
            I => data_out_0_0
        );

    \I__8594\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38121\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__38121\,
            I => \N__38117\
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__38120\,
            I => \N__38114\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__38117\,
            I => \N__38111\
        );

    \I__8590\ : InMux
    port map (
            O => \N__38114\,
            I => \N__38108\
        );

    \I__8589\ : Odrv4
    port map (
            O => \N__38111\,
            I => rand_setpoint_16
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__38108\,
            I => rand_setpoint_16
        );

    \I__8587\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38100\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__38100\,
            I => \N__38096\
        );

    \I__8585\ : CascadeMux
    port map (
            O => \N__38099\,
            I => \N__38093\
        );

    \I__8584\ : Span4Mux_v
    port map (
            O => \N__38096\,
            I => \N__38090\
        );

    \I__8583\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38087\
        );

    \I__8582\ : Odrv4
    port map (
            O => \N__38090\,
            I => rand_setpoint_15
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__38087\,
            I => rand_setpoint_15
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__38082\,
            I => \N__38079\
        );

    \I__8579\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38076\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__38076\,
            I => n10_adj_2450
        );

    \I__8577\ : CascadeMux
    port map (
            O => \N__38073\,
            I => \n10_adj_2411_cascade_\
        );

    \I__8576\ : CascadeMux
    port map (
            O => \N__38070\,
            I => \N__38066\
        );

    \I__8575\ : InMux
    port map (
            O => \N__38069\,
            I => \N__38062\
        );

    \I__8574\ : InMux
    port map (
            O => \N__38066\,
            I => \N__38059\
        );

    \I__8573\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38056\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__38062\,
            I => \N__38053\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__38059\,
            I => \N__38050\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__38056\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__8569\ : Odrv4
    port map (
            O => \N__38053\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__8568\ : Odrv12
    port map (
            O => \N__38050\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__8567\ : SRMux
    port map (
            O => \N__38043\,
            I => \N__38040\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__38040\,
            I => \N__38037\
        );

    \I__8565\ : Span4Mux_h
    port map (
            O => \N__38037\,
            I => \N__38034\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__38034\,
            I => \c0.n16718\
        );

    \I__8563\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__8561\ : Span4Mux_h
    port map (
            O => \N__38025\,
            I => \N__38022\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__38022\,
            I => \N__38019\
        );

    \I__8559\ : Span4Mux_h
    port map (
            O => \N__38019\,
            I => \N__38015\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__38018\,
            I => \N__38012\
        );

    \I__8557\ : Span4Mux_h
    port map (
            O => \N__38015\,
            I => \N__38009\
        );

    \I__8556\ : InMux
    port map (
            O => \N__38012\,
            I => \N__38006\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__38009\,
            I => rand_setpoint_0
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__38006\,
            I => rand_setpoint_0
        );

    \I__8553\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37998\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__37998\,
            I => n2
        );

    \I__8551\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37991\
        );

    \I__8550\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37988\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__37991\,
            I => data_out_2_0
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__37988\,
            I => data_out_2_0
        );

    \I__8547\ : InMux
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__8545\ : Span4Mux_v
    port map (
            O => \N__37977\,
            I => \N__37974\
        );

    \I__8544\ : Span4Mux_v
    port map (
            O => \N__37974\,
            I => \N__37970\
        );

    \I__8543\ : InMux
    port map (
            O => \N__37973\,
            I => \N__37967\
        );

    \I__8542\ : Odrv4
    port map (
            O => \N__37970\,
            I => n4_adj_2427
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__37967\,
            I => n4_adj_2427
        );

    \I__8540\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37956\
        );

    \I__8539\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37956\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37953\
        );

    \I__8537\ : Odrv12
    port map (
            O => \N__37953\,
            I => n4_adj_2416
        );

    \I__8536\ : InMux
    port map (
            O => \N__37950\,
            I => \N__37938\
        );

    \I__8535\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37938\
        );

    \I__8534\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37938\
        );

    \I__8533\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37938\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37935\
        );

    \I__8531\ : Span12Mux_h
    port map (
            O => \N__37935\,
            I => \N__37930\
        );

    \I__8530\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37925\
        );

    \I__8529\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37925\
        );

    \I__8528\ : Odrv12
    port map (
            O => \N__37930\,
            I => \r_Bit_Index_1_adj_2436\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__37925\,
            I => \r_Bit_Index_1_adj_2436\
        );

    \I__8526\ : InMux
    port map (
            O => \N__37920\,
            I => \N__37908\
        );

    \I__8525\ : InMux
    port map (
            O => \N__37919\,
            I => \N__37908\
        );

    \I__8524\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37908\
        );

    \I__8523\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37908\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__37908\,
            I => \N__37904\
        );

    \I__8521\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \N__37899\
        );

    \I__8520\ : Sp12to4
    port map (
            O => \N__37904\,
            I => \N__37896\
        );

    \I__8519\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37891\
        );

    \I__8518\ : InMux
    port map (
            O => \N__37902\,
            I => \N__37891\
        );

    \I__8517\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37888\
        );

    \I__8516\ : Span12Mux_v
    port map (
            O => \N__37896\,
            I => \N__37885\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__37891\,
            I => \N__37882\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__37888\,
            I => \r_Bit_Index_2_adj_2435\
        );

    \I__8513\ : Odrv12
    port map (
            O => \N__37885\,
            I => \r_Bit_Index_2_adj_2435\
        );

    \I__8512\ : Odrv4
    port map (
            O => \N__37882\,
            I => \r_Bit_Index_2_adj_2435\
        );

    \I__8511\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37872\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__37872\,
            I => \N__37869\
        );

    \I__8509\ : Span4Mux_v
    port map (
            O => \N__37869\,
            I => \N__37865\
        );

    \I__8508\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37862\
        );

    \I__8507\ : Span4Mux_h
    port map (
            O => \N__37865\,
            I => \N__37857\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37857\
        );

    \I__8505\ : Span4Mux_v
    port map (
            O => \N__37857\,
            I => \N__37854\
        );

    \I__8504\ : Span4Mux_h
    port map (
            O => \N__37854\,
            I => \N__37848\
        );

    \I__8503\ : InMux
    port map (
            O => \N__37853\,
            I => \N__37841\
        );

    \I__8502\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37841\
        );

    \I__8501\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37841\
        );

    \I__8500\ : Odrv4
    port map (
            O => \N__37848\,
            I => \r_Bit_Index_0\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__37841\,
            I => \r_Bit_Index_0\
        );

    \I__8498\ : InMux
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__37833\,
            I => \N__37830\
        );

    \I__8496\ : Span4Mux_h
    port map (
            O => \N__37830\,
            I => \N__37826\
        );

    \I__8495\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37823\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__37826\,
            I => \N__37818\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37818\
        );

    \I__8492\ : Span4Mux_h
    port map (
            O => \N__37818\,
            I => \N__37815\
        );

    \I__8491\ : Span4Mux_v
    port map (
            O => \N__37815\,
            I => \N__37812\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__37812\,
            I => \c0.rx.n10158\
        );

    \I__8489\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37805\
        );

    \I__8488\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37802\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__37805\,
            I => \N__37797\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__37802\,
            I => \N__37797\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__37797\,
            I => \N__37794\
        );

    \I__8484\ : Span4Mux_h
    port map (
            O => \N__37794\,
            I => \N__37790\
        );

    \I__8483\ : CascadeMux
    port map (
            O => \N__37793\,
            I => \N__37787\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__37790\,
            I => \N__37784\
        );

    \I__8481\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37781\
        );

    \I__8480\ : Span4Mux_h
    port map (
            O => \N__37784\,
            I => \N__37778\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__37781\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__37778\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__8477\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__37770\,
            I => \c0.n48\
        );

    \I__8475\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37758\
        );

    \I__8474\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37758\
        );

    \I__8473\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37758\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__37758\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__8471\ : SRMux
    port map (
            O => \N__37755\,
            I => \N__37752\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__37752\,
            I => \N__37749\
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__37749\,
            I => \c0.n16698\
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__37746\,
            I => \N__37742\
        );

    \I__8467\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37737\
        );

    \I__8466\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37721\
        );

    \I__8465\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37721\
        );

    \I__8464\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37721\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__37737\,
            I => \N__37718\
        );

    \I__8462\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37715\
        );

    \I__8461\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37710\
        );

    \I__8460\ : InMux
    port map (
            O => \N__37734\,
            I => \N__37710\
        );

    \I__8459\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37707\
        );

    \I__8458\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37704\
        );

    \I__8457\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37701\
        );

    \I__8456\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37696\
        );

    \I__8455\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37696\
        );

    \I__8454\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37693\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37687\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__37718\,
            I => \N__37682\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__37715\,
            I => \N__37682\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__37710\,
            I => \N__37671\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__37707\,
            I => \N__37671\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__37704\,
            I => \N__37671\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__37701\,
            I => \N__37671\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__37696\,
            I => \N__37671\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__37693\,
            I => \N__37668\
        );

    \I__8444\ : InMux
    port map (
            O => \N__37692\,
            I => \N__37661\
        );

    \I__8443\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37661\
        );

    \I__8442\ : InMux
    port map (
            O => \N__37690\,
            I => \N__37661\
        );

    \I__8441\ : Span4Mux_v
    port map (
            O => \N__37687\,
            I => \N__37658\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__37682\,
            I => \N__37649\
        );

    \I__8439\ : Span4Mux_v
    port map (
            O => \N__37671\,
            I => \N__37649\
        );

    \I__8438\ : Span4Mux_h
    port map (
            O => \N__37668\,
            I => \N__37649\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__37661\,
            I => \N__37649\
        );

    \I__8436\ : Odrv4
    port map (
            O => \N__37658\,
            I => \c0.n15179\
        );

    \I__8435\ : Odrv4
    port map (
            O => \N__37649\,
            I => \c0.n15179\
        );

    \I__8434\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37641\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__37641\,
            I => \c0.n17686\
        );

    \I__8432\ : InMux
    port map (
            O => \N__37638\,
            I => \N__37633\
        );

    \I__8431\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37630\
        );

    \I__8430\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37627\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37624\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__37630\,
            I => \N__37619\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__37627\,
            I => \N__37616\
        );

    \I__8426\ : Span4Mux_v
    port map (
            O => \N__37624\,
            I => \N__37613\
        );

    \I__8425\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37610\
        );

    \I__8424\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37607\
        );

    \I__8423\ : Span12Mux_s4_h
    port map (
            O => \N__37619\,
            I => \N__37600\
        );

    \I__8422\ : Span12Mux_v
    port map (
            O => \N__37616\,
            I => \N__37600\
        );

    \I__8421\ : Sp12to4
    port map (
            O => \N__37613\,
            I => \N__37600\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__37610\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__37607\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__8418\ : Odrv12
    port map (
            O => \N__37600\,
            I => \c0.data_out_frame2_0_4\
        );

    \I__8417\ : InMux
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__37590\,
            I => \c0.n17688\
        );

    \I__8415\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__37584\,
            I => \N__37577\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__37583\,
            I => \N__37574\
        );

    \I__8412\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37569\
        );

    \I__8411\ : InMux
    port map (
            O => \N__37581\,
            I => \N__37569\
        );

    \I__8410\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37565\
        );

    \I__8409\ : Span4Mux_h
    port map (
            O => \N__37577\,
            I => \N__37562\
        );

    \I__8408\ : InMux
    port map (
            O => \N__37574\,
            I => \N__37559\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__37569\,
            I => \N__37556\
        );

    \I__8406\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37553\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37550\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__37562\,
            I => \N__37547\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__37559\,
            I => \N__37542\
        );

    \I__8402\ : Span12Mux_s11_h
    port map (
            O => \N__37556\,
            I => \N__37542\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__37553\,
            I => \N__37539\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__37550\,
            I => \N__37536\
        );

    \I__8399\ : Span4Mux_h
    port map (
            O => \N__37547\,
            I => \N__37533\
        );

    \I__8398\ : Odrv12
    port map (
            O => \N__37542\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__8397\ : Odrv4
    port map (
            O => \N__37539\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__37536\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__37533\,
            I => \c0.data_out_frame2_0_3\
        );

    \I__8394\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37520\
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__37523\,
            I => \N__37517\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__37520\,
            I => \N__37514\
        );

    \I__8391\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37511\
        );

    \I__8390\ : Span4Mux_h
    port map (
            O => \N__37514\,
            I => \N__37508\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__37511\,
            I => \c0.data_in_frame_3_7\
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__37508\,
            I => \c0.data_in_frame_3_7\
        );

    \I__8387\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37499\
        );

    \I__8386\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37496\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__37499\,
            I => \c0.n2126\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__37496\,
            I => \c0.n2126\
        );

    \I__8383\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__8382\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37484\
        );

    \I__8381\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37481\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__37484\,
            I => \N__37478\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__37481\,
            I => \c0.data_in_frame_3_0\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__37478\,
            I => \c0.data_in_frame_3_0\
        );

    \I__8377\ : InMux
    port map (
            O => \N__37473\,
            I => \N__37468\
        );

    \I__8376\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37465\
        );

    \I__8375\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37461\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__37468\,
            I => \N__37458\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__37465\,
            I => \N__37455\
        );

    \I__8372\ : InMux
    port map (
            O => \N__37464\,
            I => \N__37452\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__37461\,
            I => \c0.n2138\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__37458\,
            I => \c0.n2138\
        );

    \I__8369\ : Odrv4
    port map (
            O => \N__37455\,
            I => \c0.n2138\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__37452\,
            I => \c0.n2138\
        );

    \I__8367\ : InMux
    port map (
            O => \N__37443\,
            I => \N__37440\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__37440\,
            I => \N__37435\
        );

    \I__8365\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37430\
        );

    \I__8364\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37430\
        );

    \I__8363\ : Span4Mux_h
    port map (
            O => \N__37435\,
            I => \N__37427\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__37430\,
            I => \c0.data_in_frame_2_1\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__37427\,
            I => \c0.data_in_frame_2_1\
        );

    \I__8360\ : CascadeMux
    port map (
            O => \N__37422\,
            I => \N__37419\
        );

    \I__8359\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37414\
        );

    \I__8358\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37411\
        );

    \I__8357\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37408\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__37414\,
            I => \c0.data_in_frame_2_2\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__37411\,
            I => \c0.data_in_frame_2_2\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__37408\,
            I => \c0.data_in_frame_2_2\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__37401\,
            I => \c0.n18_adj_2316_cascade_\
        );

    \I__8352\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37393\
        );

    \I__8351\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37390\
        );

    \I__8350\ : InMux
    port map (
            O => \N__37396\,
            I => \N__37386\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__37393\,
            I => \N__37381\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__37390\,
            I => \N__37381\
        );

    \I__8347\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37373\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__37386\,
            I => \N__37370\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__37381\,
            I => \N__37367\
        );

    \I__8344\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37364\
        );

    \I__8343\ : InMux
    port map (
            O => \N__37379\,
            I => \N__37357\
        );

    \I__8342\ : InMux
    port map (
            O => \N__37378\,
            I => \N__37357\
        );

    \I__8341\ : InMux
    port map (
            O => \N__37377\,
            I => \N__37357\
        );

    \I__8340\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37354\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__37373\,
            I => \c0.data_in_frame_0_7\
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__37370\,
            I => \c0.data_in_frame_0_7\
        );

    \I__8337\ : Odrv4
    port map (
            O => \N__37367\,
            I => \c0.data_in_frame_0_7\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__37364\,
            I => \c0.data_in_frame_0_7\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__37357\,
            I => \c0.data_in_frame_0_7\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__37354\,
            I => \c0.data_in_frame_0_7\
        );

    \I__8333\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37338\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__37338\,
            I => \c0.n23_adj_2322\
        );

    \I__8331\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37331\
        );

    \I__8330\ : CascadeMux
    port map (
            O => \N__37334\,
            I => \N__37328\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37324\
        );

    \I__8328\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37321\
        );

    \I__8327\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37318\
        );

    \I__8326\ : Span4Mux_h
    port map (
            O => \N__37324\,
            I => \N__37315\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__37321\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__37318\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__37315\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__8322\ : SRMux
    port map (
            O => \N__37308\,
            I => \N__37305\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__37305\,
            I => \N__37302\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__37302\,
            I => \c0.n13381\
        );

    \I__8319\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37296\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__37296\,
            I => \N__37292\
        );

    \I__8317\ : CascadeMux
    port map (
            O => \N__37295\,
            I => \N__37289\
        );

    \I__8316\ : Span4Mux_v
    port map (
            O => \N__37292\,
            I => \N__37286\
        );

    \I__8315\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37282\
        );

    \I__8314\ : Span4Mux_h
    port map (
            O => \N__37286\,
            I => \N__37279\
        );

    \I__8313\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37276\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__37282\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__8311\ : Odrv4
    port map (
            O => \N__37279\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__37276\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__8309\ : SRMux
    port map (
            O => \N__37269\,
            I => \N__37266\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__37266\,
            I => \N__37263\
        );

    \I__8307\ : Span4Mux_v
    port map (
            O => \N__37263\,
            I => \N__37260\
        );

    \I__8306\ : Span4Mux_h
    port map (
            O => \N__37260\,
            I => \N__37257\
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__37257\,
            I => \c0.n8_adj_2333\
        );

    \I__8304\ : CascadeMux
    port map (
            O => \N__37254\,
            I => \N__37249\
        );

    \I__8303\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37246\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__37252\,
            I => \N__37242\
        );

    \I__8301\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37239\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37246\,
            I => \N__37235\
        );

    \I__8299\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37232\
        );

    \I__8298\ : InMux
    port map (
            O => \N__37242\,
            I => \N__37229\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__37239\,
            I => \N__37226\
        );

    \I__8296\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37223\
        );

    \I__8295\ : Span12Mux_h
    port map (
            O => \N__37235\,
            I => \N__37220\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__37232\,
            I => \N__37215\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__37229\,
            I => \N__37215\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__37226\,
            I => \N__37212\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__37223\,
            I => data_out_frame2_8_2
        );

    \I__8290\ : Odrv12
    port map (
            O => \N__37220\,
            I => data_out_frame2_8_2
        );

    \I__8289\ : Odrv4
    port map (
            O => \N__37215\,
            I => data_out_frame2_8_2
        );

    \I__8288\ : Odrv4
    port map (
            O => \N__37212\,
            I => data_out_frame2_8_2
        );

    \I__8287\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37200\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37197\
        );

    \I__8285\ : Span12Mux_s6_h
    port map (
            O => \N__37197\,
            I => \N__37194\
        );

    \I__8284\ : Odrv12
    port map (
            O => \N__37194\,
            I => \c0.n16\
        );

    \I__8283\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37188\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__37188\,
            I => \N__37182\
        );

    \I__8281\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37179\
        );

    \I__8280\ : InMux
    port map (
            O => \N__37186\,
            I => \N__37176\
        );

    \I__8279\ : InMux
    port map (
            O => \N__37185\,
            I => \N__37171\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__37182\,
            I => \N__37168\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__37179\,
            I => \N__37163\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__37176\,
            I => \N__37163\
        );

    \I__8275\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37160\
        );

    \I__8274\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37157\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__37171\,
            I => \N__37152\
        );

    \I__8272\ : Span4Mux_h
    port map (
            O => \N__37168\,
            I => \N__37143\
        );

    \I__8271\ : Span4Mux_v
    port map (
            O => \N__37163\,
            I => \N__37143\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__37160\,
            I => \N__37143\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37143\
        );

    \I__8268\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37140\
        );

    \I__8267\ : InMux
    port map (
            O => \N__37155\,
            I => \N__37137\
        );

    \I__8266\ : Span4Mux_v
    port map (
            O => \N__37152\,
            I => \N__37132\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__37143\,
            I => \N__37132\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__37140\,
            I => \N__37129\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__37137\,
            I => \N__37126\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__37132\,
            I => \N__37123\
        );

    \I__8261\ : Span4Mux_h
    port map (
            O => \N__37129\,
            I => \N__37120\
        );

    \I__8260\ : Odrv4
    port map (
            O => \N__37126\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__37123\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__8258\ : Odrv4
    port map (
            O => \N__37120\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__8257\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37109\
        );

    \I__8256\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37106\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__37109\,
            I => \N__37102\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37099\
        );

    \I__8253\ : InMux
    port map (
            O => \N__37105\,
            I => \N__37096\
        );

    \I__8252\ : Span4Mux_v
    port map (
            O => \N__37102\,
            I => \N__37089\
        );

    \I__8251\ : Span4Mux_h
    port map (
            O => \N__37099\,
            I => \N__37089\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__37096\,
            I => \N__37089\
        );

    \I__8249\ : Span4Mux_h
    port map (
            O => \N__37089\,
            I => \N__37085\
        );

    \I__8248\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37082\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__37085\,
            I => \N__37074\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__37082\,
            I => \N__37071\
        );

    \I__8245\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37062\
        );

    \I__8244\ : InMux
    port map (
            O => \N__37080\,
            I => \N__37062\
        );

    \I__8243\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37062\
        );

    \I__8242\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37062\
        );

    \I__8241\ : InMux
    port map (
            O => \N__37077\,
            I => \N__37059\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__37074\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__8239\ : Odrv4
    port map (
            O => \N__37071\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__37062\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__37059\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__8236\ : CascadeMux
    port map (
            O => \N__37050\,
            I => \c0.n15171_cascade_\
        );

    \I__8235\ : CascadeMux
    port map (
            O => \N__37047\,
            I => \N__37040\
        );

    \I__8234\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37037\
        );

    \I__8233\ : InMux
    port map (
            O => \N__37045\,
            I => \N__37034\
        );

    \I__8232\ : InMux
    port map (
            O => \N__37044\,
            I => \N__37029\
        );

    \I__8231\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37029\
        );

    \I__8230\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37026\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__37037\,
            I => \c0.data_in_frame_1_6\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__37034\,
            I => \c0.data_in_frame_1_6\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__37029\,
            I => \c0.data_in_frame_1_6\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__37026\,
            I => \c0.data_in_frame_1_6\
        );

    \I__8225\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__37014\,
            I => \N__37011\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__37011\,
            I => \N__37007\
        );

    \I__8222\ : InMux
    port map (
            O => \N__37010\,
            I => \N__37004\
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__37007\,
            I => \c0.n2124\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__37004\,
            I => \c0.n2124\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__8218\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36989\
        );

    \I__8216\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36986\
        );

    \I__8215\ : Span4Mux_v
    port map (
            O => \N__36989\,
            I => \N__36983\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__36986\,
            I => data_in_frame_6_6
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__36983\,
            I => data_in_frame_6_6
        );

    \I__8212\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36975\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__36975\,
            I => \c0.n17214\
        );

    \I__8210\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36969\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__36969\,
            I => \c0.n28_adj_2374\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__36966\,
            I => \c0.n27_adj_2381_cascade_\
        );

    \I__8207\ : InMux
    port map (
            O => \N__36963\,
            I => \N__36960\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__36960\,
            I => \c0.n29\
        );

    \I__8205\ : CascadeMux
    port map (
            O => \N__36957\,
            I => \c0.n12491_cascade_\
        );

    \I__8204\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36950\
        );

    \I__8203\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36944\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__36950\,
            I => \N__36941\
        );

    \I__8201\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36938\
        );

    \I__8200\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36935\
        );

    \I__8199\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36932\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__36944\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8197\ : Odrv4
    port map (
            O => \N__36941\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__36938\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__36935\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__36932\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8193\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36918\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36914\
        );

    \I__8191\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36911\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__36914\,
            I => \c0.n10259\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__36911\,
            I => \c0.n10259\
        );

    \I__8188\ : InMux
    port map (
            O => \N__36906\,
            I => \N__36903\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__36903\,
            I => \N__36899\
        );

    \I__8186\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36895\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__36899\,
            I => \N__36892\
        );

    \I__8184\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36889\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__36895\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8182\ : Odrv4
    port map (
            O => \N__36892\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__36889\,
            I => \c0.data_in_frame_2_7\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__36882\,
            I => \N__36878\
        );

    \I__8179\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36873\
        );

    \I__8178\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36870\
        );

    \I__8177\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36867\
        );

    \I__8176\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36864\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__36873\,
            I => \N__36858\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__36870\,
            I => \N__36853\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__36867\,
            I => \N__36853\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__36864\,
            I => \N__36850\
        );

    \I__8171\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36847\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__36862\,
            I => \N__36844\
        );

    \I__8169\ : CascadeMux
    port map (
            O => \N__36861\,
            I => \N__36841\
        );

    \I__8168\ : Span4Mux_v
    port map (
            O => \N__36858\,
            I => \N__36835\
        );

    \I__8167\ : Span4Mux_v
    port map (
            O => \N__36853\,
            I => \N__36835\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__36850\,
            I => \N__36830\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__36847\,
            I => \N__36830\
        );

    \I__8164\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36827\
        );

    \I__8163\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36824\
        );

    \I__8162\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36821\
        );

    \I__8161\ : Span4Mux_h
    port map (
            O => \N__36835\,
            I => \N__36818\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__36830\,
            I => \N__36815\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__36827\,
            I => rx_data_2
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__36824\,
            I => rx_data_2
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__36821\,
            I => rx_data_2
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__36818\,
            I => rx_data_2
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__36815\,
            I => rx_data_2
        );

    \I__8154\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36795\
        );

    \I__8153\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36790\
        );

    \I__8152\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36790\
        );

    \I__8151\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36787\
        );

    \I__8150\ : InMux
    port map (
            O => \N__36800\,
            I => \N__36782\
        );

    \I__8149\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36782\
        );

    \I__8148\ : InMux
    port map (
            O => \N__36798\,
            I => \N__36779\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__36795\,
            I => \N__36775\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__36790\,
            I => \N__36770\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__36787\,
            I => \N__36770\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__36782\,
            I => \N__36765\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__36779\,
            I => \N__36765\
        );

    \I__8142\ : CascadeMux
    port map (
            O => \N__36778\,
            I => \N__36762\
        );

    \I__8141\ : Span4Mux_h
    port map (
            O => \N__36775\,
            I => \N__36757\
        );

    \I__8140\ : Span4Mux_h
    port map (
            O => \N__36770\,
            I => \N__36757\
        );

    \I__8139\ : Span4Mux_v
    port map (
            O => \N__36765\,
            I => \N__36754\
        );

    \I__8138\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36751\
        );

    \I__8137\ : Span4Mux_h
    port map (
            O => \N__36757\,
            I => \N__36748\
        );

    \I__8136\ : Span4Mux_h
    port map (
            O => \N__36754\,
            I => \N__36745\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__36751\,
            I => rx_data_0
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__36748\,
            I => rx_data_0
        );

    \I__8133\ : Odrv4
    port map (
            O => \N__36745\,
            I => rx_data_0
        );

    \I__8132\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36735\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36732\
        );

    \I__8130\ : Sp12to4
    port map (
            O => \N__36732\,
            I => \N__36729\
        );

    \I__8129\ : Span12Mux_v
    port map (
            O => \N__36729\,
            I => \N__36726\
        );

    \I__8128\ : Span12Mux_h
    port map (
            O => \N__36726\,
            I => \N__36723\
        );

    \I__8127\ : Odrv12
    port map (
            O => \N__36723\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__8126\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36711\
        );

    \I__8125\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36711\
        );

    \I__8124\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36711\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__36711\,
            I => \N__36707\
        );

    \I__8122\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36704\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__36707\,
            I => \N__36699\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__36704\,
            I => \N__36699\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__36699\,
            I => \N__36696\
        );

    \I__8118\ : Span4Mux_v
    port map (
            O => \N__36696\,
            I => \N__36693\
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__36693\,
            I => n10010
        );

    \I__8116\ : CascadeMux
    port map (
            O => \N__36690\,
            I => \N__36684\
        );

    \I__8115\ : CascadeMux
    port map (
            O => \N__36689\,
            I => \N__36681\
        );

    \I__8114\ : CascadeMux
    port map (
            O => \N__36688\,
            I => \N__36676\
        );

    \I__8113\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36670\
        );

    \I__8112\ : InMux
    port map (
            O => \N__36684\,
            I => \N__36670\
        );

    \I__8111\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36665\
        );

    \I__8110\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36665\
        );

    \I__8109\ : InMux
    port map (
            O => \N__36679\,
            I => \N__36662\
        );

    \I__8108\ : InMux
    port map (
            O => \N__36676\,
            I => \N__36659\
        );

    \I__8107\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36656\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__36670\,
            I => \N__36652\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__36665\,
            I => \N__36649\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__36662\,
            I => \N__36646\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__36659\,
            I => \N__36641\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36641\
        );

    \I__8101\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36638\
        );

    \I__8100\ : Span4Mux_h
    port map (
            O => \N__36652\,
            I => \N__36635\
        );

    \I__8099\ : Span4Mux_h
    port map (
            O => \N__36649\,
            I => \N__36632\
        );

    \I__8098\ : Span4Mux_v
    port map (
            O => \N__36646\,
            I => \N__36627\
        );

    \I__8097\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36627\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__36638\,
            I => rx_data_5
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__36635\,
            I => rx_data_5
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__36632\,
            I => rx_data_5
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__36627\,
            I => rx_data_5
        );

    \I__8092\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36615\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__36615\,
            I => \N__36612\
        );

    \I__8090\ : Odrv12
    port map (
            O => \N__36612\,
            I => \c0.n24_adj_2317\
        );

    \I__8089\ : CascadeMux
    port map (
            O => \N__36609\,
            I => \N__36606\
        );

    \I__8088\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36603\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__36603\,
            I => \N__36600\
        );

    \I__8086\ : Odrv4
    port map (
            O => \N__36600\,
            I => \c0.n22_adj_2319\
        );

    \I__8085\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36594\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__36594\,
            I => \c0.n21_adj_2323\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__36591\,
            I => \N__36588\
        );

    \I__8082\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36585\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__36585\,
            I => \c0.n22_adj_2313\
        );

    \I__8080\ : InMux
    port map (
            O => \N__36582\,
            I => \c0.n16071\
        );

    \I__8079\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36576\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__36576\,
            I => \c0.n21_adj_2262\
        );

    \I__8077\ : InMux
    port map (
            O => \N__36573\,
            I => \c0.n16072\
        );

    \I__8076\ : InMux
    port map (
            O => \N__36570\,
            I => \bfn_12_32_0_\
        );

    \I__8075\ : InMux
    port map (
            O => \N__36567\,
            I => \c0.n16074\
        );

    \I__8074\ : InMux
    port map (
            O => \N__36564\,
            I => \c0.n16075\
        );

    \I__8073\ : InMux
    port map (
            O => \N__36561\,
            I => \c0.n16076\
        );

    \I__8072\ : InMux
    port map (
            O => \N__36558\,
            I => \c0.n16077\
        );

    \I__8071\ : InMux
    port map (
            O => \N__36555\,
            I => \c0.n16078\
        );

    \I__8070\ : CEMux
    port map (
            O => \N__36552\,
            I => \N__36548\
        );

    \I__8069\ : CEMux
    port map (
            O => \N__36551\,
            I => \N__36545\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__36548\,
            I => \N__36542\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__36545\,
            I => \N__36539\
        );

    \I__8066\ : Span4Mux_h
    port map (
            O => \N__36542\,
            I => \N__36536\
        );

    \I__8065\ : Span4Mux_s2_v
    port map (
            O => \N__36539\,
            I => \N__36533\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__36536\,
            I => \c0.n10594\
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__36533\,
            I => \c0.n10594\
        );

    \I__8062\ : InMux
    port map (
            O => \N__36528\,
            I => \N__36525\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__36525\,
            I => \c0.n16353\
        );

    \I__8060\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36519\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__36516\,
            I => \c0.n26_adj_2368\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__36513\,
            I => \N__36510\
        );

    \I__8056\ : InMux
    port map (
            O => \N__36510\,
            I => \N__36507\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__36507\,
            I => \N__36504\
        );

    \I__8054\ : Odrv12
    port map (
            O => \N__36504\,
            I => \c0.n16474\
        );

    \I__8053\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36498\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__36498\,
            I => \c0.n18_adj_2360\
        );

    \I__8051\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36492\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__36492\,
            I => \c0.n27\
        );

    \I__8049\ : InMux
    port map (
            O => \N__36489\,
            I => \c0.n16066\
        );

    \I__8048\ : InMux
    port map (
            O => \N__36486\,
            I => \c0.n16067\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__36483\,
            I => \N__36480\
        );

    \I__8046\ : InMux
    port map (
            O => \N__36480\,
            I => \N__36477\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__36477\,
            I => \c0.n25_adj_2386\
        );

    \I__8044\ : InMux
    port map (
            O => \N__36474\,
            I => \c0.n16068\
        );

    \I__8043\ : InMux
    port map (
            O => \N__36471\,
            I => \c0.n16069\
        );

    \I__8042\ : InMux
    port map (
            O => \N__36468\,
            I => \c0.n16070\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__36465\,
            I => \n4_adj_2419_cascade_\
        );

    \I__8040\ : CascadeMux
    port map (
            O => \N__36462\,
            I => \n5_adj_2407_cascade_\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__36459\,
            I => \n10_adj_2444_cascade_\
        );

    \I__8038\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36453\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__36453\,
            I => n8_adj_2447
        );

    \I__8036\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36447\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__36447\,
            I => n4_adj_2419
        );

    \I__8034\ : InMux
    port map (
            O => \N__36444\,
            I => \N__36441\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__36441\,
            I => \N__36438\
        );

    \I__8032\ : Span4Mux_v
    port map (
            O => \N__36438\,
            I => \N__36435\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__36435\,
            I => \c0.n17696\
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__36432\,
            I => \n18073_cascade_\
        );

    \I__8029\ : CascadeMux
    port map (
            O => \N__36429\,
            I => \c0.tx.n10688_cascade_\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__36426\,
            I => \N__36422\
        );

    \I__8027\ : InMux
    port map (
            O => \N__36425\,
            I => \N__36417\
        );

    \I__8026\ : InMux
    port map (
            O => \N__36422\,
            I => \N__36417\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__36417\,
            I => \r_Tx_Data_1\
        );

    \I__8024\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36411\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__36411\,
            I => \N__36407\
        );

    \I__8022\ : CascadeMux
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__8021\ : Span4Mux_v
    port map (
            O => \N__36407\,
            I => \N__36401\
        );

    \I__8020\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36398\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__36401\,
            I => rand_setpoint_1
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__36398\,
            I => rand_setpoint_1
        );

    \I__8017\ : InMux
    port map (
            O => \N__36393\,
            I => \N__36389\
        );

    \I__8016\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__36389\,
            I => \N__36383\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__36386\,
            I => \r_Tx_Data_3\
        );

    \I__8013\ : Odrv4
    port map (
            O => \N__36383\,
            I => \r_Tx_Data_3\
        );

    \I__8012\ : InMux
    port map (
            O => \N__36378\,
            I => \N__36375\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__36375\,
            I => n18070
        );

    \I__8010\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36367\
        );

    \I__8009\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36362\
        );

    \I__8008\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36362\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__36367\,
            I => \c0.tx.n10688\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__36362\,
            I => \c0.tx.n10688\
        );

    \I__8005\ : CascadeMux
    port map (
            O => \N__36357\,
            I => \n10_adj_2409_cascade_\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__36354\,
            I => \c0.n8_adj_2183_cascade_\
        );

    \I__8003\ : InMux
    port map (
            O => \N__36351\,
            I => \N__36348\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__36348\,
            I => \c0.n17671\
        );

    \I__8001\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36342\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__36342\,
            I => \N__36339\
        );

    \I__7999\ : Span4Mux_h
    port map (
            O => \N__36339\,
            I => \N__36335\
        );

    \I__7998\ : CascadeMux
    port map (
            O => \N__36338\,
            I => \N__36332\
        );

    \I__7997\ : Sp12to4
    port map (
            O => \N__36335\,
            I => \N__36329\
        );

    \I__7996\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36326\
        );

    \I__7995\ : Odrv12
    port map (
            O => \N__36329\,
            I => rand_setpoint_4
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__36326\,
            I => rand_setpoint_4
        );

    \I__7993\ : CascadeMux
    port map (
            O => \N__36321\,
            I => \data_out_10__7__N_110_cascade_\
        );

    \I__7992\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36315\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36311\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__36314\,
            I => \N__36308\
        );

    \I__7989\ : Span4Mux_h
    port map (
            O => \N__36311\,
            I => \N__36305\
        );

    \I__7988\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36302\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__36305\,
            I => rand_setpoint_6
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__36302\,
            I => rand_setpoint_6
        );

    \I__7985\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36294\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36290\
        );

    \I__7983\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36287\
        );

    \I__7982\ : Span4Mux_h
    port map (
            O => \N__36290\,
            I => \N__36284\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__36287\,
            I => \c0.data_out_1_2\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__36284\,
            I => \c0.data_out_1_2\
        );

    \I__7979\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__36276\,
            I => \N__36272\
        );

    \I__7977\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36269\
        );

    \I__7976\ : Span4Mux_v
    port map (
            O => \N__36272\,
            I => \N__36266\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__36269\,
            I => \N__36263\
        );

    \I__7974\ : Span4Mux_h
    port map (
            O => \N__36266\,
            I => \N__36258\
        );

    \I__7973\ : Span4Mux_v
    port map (
            O => \N__36263\,
            I => \N__36258\
        );

    \I__7972\ : Span4Mux_v
    port map (
            O => \N__36258\,
            I => \N__36254\
        );

    \I__7971\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36251\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__36254\,
            I => blink_counter_24
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__36251\,
            I => blink_counter_24
        );

    \I__7968\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36242\
        );

    \I__7967\ : InMux
    port map (
            O => \N__36245\,
            I => \N__36239\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36236\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__36239\,
            I => \N__36233\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__36236\,
            I => \N__36230\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__36233\,
            I => \N__36227\
        );

    \I__7962\ : Span4Mux_v
    port map (
            O => \N__36230\,
            I => \N__36223\
        );

    \I__7961\ : Span4Mux_v
    port map (
            O => \N__36227\,
            I => \N__36220\
        );

    \I__7960\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36217\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__36223\,
            I => blink_counter_23
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__36220\,
            I => blink_counter_23
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__36217\,
            I => blink_counter_23
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__36210\,
            I => \N__36207\
        );

    \I__7955\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36204\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__36204\,
            I => \N__36200\
        );

    \I__7953\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36197\
        );

    \I__7952\ : Span4Mux_v
    port map (
            O => \N__36200\,
            I => \N__36194\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__36197\,
            I => \N__36191\
        );

    \I__7950\ : Span4Mux_v
    port map (
            O => \N__36194\,
            I => \N__36187\
        );

    \I__7949\ : Span12Mux_v
    port map (
            O => \N__36191\,
            I => \N__36184\
        );

    \I__7948\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36181\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__36187\,
            I => blink_counter_22
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__36184\,
            I => blink_counter_22
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__36181\,
            I => blink_counter_22
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__36174\,
            I => \N__36171\
        );

    \I__7943\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36167\
        );

    \I__7942\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36164\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__36167\,
            I => \N__36161\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__36164\,
            I => \N__36158\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__36161\,
            I => \N__36155\
        );

    \I__7938\ : Span12Mux_v
    port map (
            O => \N__36158\,
            I => \N__36151\
        );

    \I__7937\ : Span4Mux_v
    port map (
            O => \N__36155\,
            I => \N__36148\
        );

    \I__7936\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36145\
        );

    \I__7935\ : Odrv12
    port map (
            O => \N__36151\,
            I => blink_counter_21
        );

    \I__7934\ : Odrv4
    port map (
            O => \N__36148\,
            I => blink_counter_21
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__36145\,
            I => blink_counter_21
        );

    \I__7932\ : InMux
    port map (
            O => \N__36138\,
            I => \N__36135\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36132\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__36132\,
            I => n10140
        );

    \I__7929\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36126\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__36126\,
            I => n8
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__36123\,
            I => \n4_adj_2417_cascade_\
        );

    \I__7926\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36115\
        );

    \I__7925\ : InMux
    port map (
            O => \N__36119\,
            I => \N__36110\
        );

    \I__7924\ : InMux
    port map (
            O => \N__36118\,
            I => \N__36110\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36104\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__36110\,
            I => \N__36104\
        );

    \I__7921\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36101\
        );

    \I__7920\ : Span4Mux_v
    port map (
            O => \N__36104\,
            I => \N__36096\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__36101\,
            I => \N__36096\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__36096\,
            I => \FRAME_MATCHER_state_31_N_1406_2\
        );

    \I__7917\ : CascadeMux
    port map (
            O => \N__36093\,
            I => \N__36087\
        );

    \I__7916\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36083\
        );

    \I__7915\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36078\
        );

    \I__7914\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36078\
        );

    \I__7913\ : InMux
    port map (
            O => \N__36087\,
            I => \N__36073\
        );

    \I__7912\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36073\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__36083\,
            I => \N__36066\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__36078\,
            I => \N__36063\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__36073\,
            I => \N__36058\
        );

    \I__7908\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36055\
        );

    \I__7907\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36050\
        );

    \I__7906\ : InMux
    port map (
            O => \N__36070\,
            I => \N__36050\
        );

    \I__7905\ : InMux
    port map (
            O => \N__36069\,
            I => \N__36047\
        );

    \I__7904\ : Span12Mux_v
    port map (
            O => \N__36066\,
            I => \N__36044\
        );

    \I__7903\ : Span4Mux_v
    port map (
            O => \N__36063\,
            I => \N__36041\
        );

    \I__7902\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36036\
        );

    \I__7901\ : InMux
    port map (
            O => \N__36061\,
            I => \N__36036\
        );

    \I__7900\ : Span4Mux_h
    port map (
            O => \N__36058\,
            I => \N__36031\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__36055\,
            I => \N__36031\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__36050\,
            I => \N__36028\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__36047\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__7896\ : Odrv12
    port map (
            O => \N__36044\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__7895\ : Odrv4
    port map (
            O => \N__36041\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__36036\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__36031\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__7892\ : Odrv4
    port map (
            O => \N__36028\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__7891\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__36012\,
            I => \N__36009\
        );

    \I__7889\ : Span4Mux_v
    port map (
            O => \N__36009\,
            I => \N__36006\
        );

    \I__7888\ : Span4Mux_v
    port map (
            O => \N__36006\,
            I => \N__36002\
        );

    \I__7887\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35999\
        );

    \I__7886\ : Odrv4
    port map (
            O => \N__36002\,
            I => blink_counter_25
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__35999\,
            I => blink_counter_25
        );

    \I__7884\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35991\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__35991\,
            I => n17428
        );

    \I__7882\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35985\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__35985\,
            I => \N__35982\
        );

    \I__7880\ : Span4Mux_v
    port map (
            O => \N__35982\,
            I => \N__35979\
        );

    \I__7879\ : Odrv4
    port map (
            O => \N__35979\,
            I => n17427
        );

    \I__7878\ : IoInMux
    port map (
            O => \N__35976\,
            I => \N__35973\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__35973\,
            I => \N__35970\
        );

    \I__7876\ : Span4Mux_s3_v
    port map (
            O => \N__35970\,
            I => \N__35967\
        );

    \I__7875\ : Span4Mux_v
    port map (
            O => \N__35967\,
            I => \N__35964\
        );

    \I__7874\ : Sp12to4
    port map (
            O => \N__35964\,
            I => \N__35961\
        );

    \I__7873\ : Odrv12
    port map (
            O => \N__35961\,
            I => \LED_c\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__35958\,
            I => \N__35954\
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__35957\,
            I => \N__35951\
        );

    \I__7870\ : InMux
    port map (
            O => \N__35954\,
            I => \N__35947\
        );

    \I__7869\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35942\
        );

    \I__7868\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35942\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__35947\,
            I => \N__35937\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__35942\,
            I => \N__35934\
        );

    \I__7865\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35929\
        );

    \I__7864\ : InMux
    port map (
            O => \N__35940\,
            I => \N__35929\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__35937\,
            I => \N__35926\
        );

    \I__7862\ : Span4Mux_h
    port map (
            O => \N__35934\,
            I => \N__35923\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__35929\,
            I => \N__35920\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__35926\,
            I => \N__35917\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__35923\,
            I => \N__35914\
        );

    \I__7858\ : Span4Mux_v
    port map (
            O => \N__35920\,
            I => \N__35911\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__35917\,
            I => n3779
        );

    \I__7856\ : Odrv4
    port map (
            O => \N__35914\,
            I => n3779
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__35911\,
            I => n3779
        );

    \I__7854\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35899\
        );

    \I__7853\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35896\
        );

    \I__7852\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35893\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__35899\,
            I => \N__35888\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35883\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__35893\,
            I => \N__35883\
        );

    \I__7848\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35878\
        );

    \I__7847\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35878\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__35888\,
            I => \FRAME_MATCHER_i_31__N_1273\
        );

    \I__7845\ : Odrv4
    port map (
            O => \N__35883\,
            I => \FRAME_MATCHER_i_31__N_1273\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__35878\,
            I => \FRAME_MATCHER_i_31__N_1273\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__7842\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__35865\,
            I => n6_adj_2488
        );

    \I__7840\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35859\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__35859\,
            I => \N__35855\
        );

    \I__7838\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35852\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__35855\,
            I => \N__35849\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__35852\,
            I => data_out_3_0
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__35849\,
            I => data_out_3_0
        );

    \I__7834\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35841\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__35841\,
            I => \N__35838\
        );

    \I__7832\ : Span4Mux_h
    port map (
            O => \N__35838\,
            I => \N__35835\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__35835\,
            I => n18175
        );

    \I__7830\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35829\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__35829\,
            I => \N__35825\
        );

    \I__7828\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35822\
        );

    \I__7827\ : Span12Mux_s11_h
    port map (
            O => \N__35825\,
            I => \N__35814\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35811\
        );

    \I__7825\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35806\
        );

    \I__7824\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35806\
        );

    \I__7823\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35799\
        );

    \I__7822\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35799\
        );

    \I__7821\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35799\
        );

    \I__7820\ : Odrv12
    port map (
            O => \N__35814\,
            I => n5
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__35811\,
            I => n5
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__35806\,
            I => n5
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__35799\,
            I => n5
        );

    \I__7816\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35787\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__35787\,
            I => \N__35783\
        );

    \I__7814\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35780\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__35783\,
            I => n1_adj_2486
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__35780\,
            I => n1_adj_2486
        );

    \I__7811\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35772\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__35772\,
            I => \N__35769\
        );

    \I__7809\ : Odrv4
    port map (
            O => \N__35769\,
            I => n9378
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__35766\,
            I => \N__35762\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__35765\,
            I => \N__35759\
        );

    \I__7806\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35754\
        );

    \I__7805\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35751\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__35758\,
            I => \N__35747\
        );

    \I__7803\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35740\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__35754\,
            I => \N__35737\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35734\
        );

    \I__7800\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35729\
        );

    \I__7799\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35729\
        );

    \I__7798\ : CascadeMux
    port map (
            O => \N__35746\,
            I => \N__35726\
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__35745\,
            I => \N__35720\
        );

    \I__7796\ : CascadeMux
    port map (
            O => \N__35744\,
            I => \N__35716\
        );

    \I__7795\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35713\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__35740\,
            I => \N__35708\
        );

    \I__7793\ : Span4Mux_h
    port map (
            O => \N__35737\,
            I => \N__35705\
        );

    \I__7792\ : Span4Mux_h
    port map (
            O => \N__35734\,
            I => \N__35699\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__35729\,
            I => \N__35696\
        );

    \I__7790\ : InMux
    port map (
            O => \N__35726\,
            I => \N__35693\
        );

    \I__7789\ : InMux
    port map (
            O => \N__35725\,
            I => \N__35690\
        );

    \I__7788\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35683\
        );

    \I__7787\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35683\
        );

    \I__7786\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35683\
        );

    \I__7785\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35679\
        );

    \I__7784\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35676\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35673\
        );

    \I__7782\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35668\
        );

    \I__7781\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35668\
        );

    \I__7780\ : Span4Mux_v
    port map (
            O => \N__35708\,
            I => \N__35663\
        );

    \I__7779\ : Span4Mux_v
    port map (
            O => \N__35705\,
            I => \N__35663\
        );

    \I__7778\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35660\
        );

    \I__7777\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35655\
        );

    \I__7776\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35655\
        );

    \I__7775\ : Span4Mux_v
    port map (
            O => \N__35699\,
            I => \N__35644\
        );

    \I__7774\ : Span4Mux_h
    port map (
            O => \N__35696\,
            I => \N__35644\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__35693\,
            I => \N__35644\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__35690\,
            I => \N__35644\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35644\
        );

    \I__7770\ : InMux
    port map (
            O => \N__35682\,
            I => \N__35641\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__35679\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__35676\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7767\ : Odrv12
    port map (
            O => \N__35673\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__35668\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7765\ : Odrv4
    port map (
            O => \N__35663\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__35660\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__35655\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__35644\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__35641\,
            I => \FRAME_MATCHER_state_1\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__35622\,
            I => \N__35619\
        );

    \I__7759\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35616\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__35616\,
            I => \N__35613\
        );

    \I__7757\ : Odrv12
    port map (
            O => \N__35613\,
            I => \c0.n16261\
        );

    \I__7756\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35607\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__35607\,
            I => \N__35602\
        );

    \I__7754\ : InMux
    port map (
            O => \N__35606\,
            I => \N__35599\
        );

    \I__7753\ : CascadeMux
    port map (
            O => \N__35605\,
            I => \N__35596\
        );

    \I__7752\ : Span4Mux_h
    port map (
            O => \N__35602\,
            I => \N__35590\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35590\
        );

    \I__7750\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35587\
        );

    \I__7749\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35584\
        );

    \I__7748\ : Span4Mux_h
    port map (
            O => \N__35590\,
            I => \N__35579\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__35587\,
            I => \N__35574\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35574\
        );

    \I__7745\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35569\
        );

    \I__7744\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35569\
        );

    \I__7743\ : Span4Mux_v
    port map (
            O => \N__35579\,
            I => \N__35566\
        );

    \I__7742\ : Span12Mux_s11_h
    port map (
            O => \N__35574\,
            I => \N__35563\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__35569\,
            I => \N__35560\
        );

    \I__7740\ : Odrv4
    port map (
            O => \N__35566\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2167\
        );

    \I__7739\ : Odrv12
    port map (
            O => \N__35563\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2167\
        );

    \I__7738\ : Odrv12
    port map (
            O => \N__35560\,
            I => \c0.r_SM_Main_2_N_2034_0_adj_2167\
        );

    \I__7737\ : SRMux
    port map (
            O => \N__35553\,
            I => \N__35546\
        );

    \I__7736\ : InMux
    port map (
            O => \N__35552\,
            I => \N__35541\
        );

    \I__7735\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35541\
        );

    \I__7734\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35536\
        );

    \I__7733\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35536\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__35546\,
            I => \N__35529\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__35541\,
            I => \N__35526\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__35536\,
            I => \N__35523\
        );

    \I__7729\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35518\
        );

    \I__7728\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35518\
        );

    \I__7727\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35515\
        );

    \I__7726\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35512\
        );

    \I__7725\ : Odrv12
    port map (
            O => \N__35529\,
            I => \c0.n10018\
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__35526\,
            I => \c0.n10018\
        );

    \I__7723\ : Odrv4
    port map (
            O => \N__35523\,
            I => \c0.n10018\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__35518\,
            I => \c0.n10018\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__35515\,
            I => \c0.n10018\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__35512\,
            I => \c0.n10018\
        );

    \I__7719\ : InMux
    port map (
            O => \N__35499\,
            I => \N__35496\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__35496\,
            I => n10088
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__35493\,
            I => \N__35489\
        );

    \I__7716\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35486\
        );

    \I__7715\ : InMux
    port map (
            O => \N__35489\,
            I => \N__35483\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__35486\,
            I => \N__35480\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__35483\,
            I => \N__35477\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__35480\,
            I => \N__35474\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__35477\,
            I => \N__35471\
        );

    \I__7710\ : Span4Mux_h
    port map (
            O => \N__35474\,
            I => \N__35468\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__35471\,
            I => n17086
        );

    \I__7708\ : Odrv4
    port map (
            O => \N__35468\,
            I => n17086
        );

    \I__7707\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35457\
        );

    \I__7706\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35457\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__35457\,
            I => n17063
        );

    \I__7704\ : InMux
    port map (
            O => \N__35454\,
            I => \N__35448\
        );

    \I__7703\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35448\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__35448\,
            I => n17089
        );

    \I__7701\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35442\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__35442\,
            I => n17090
        );

    \I__7699\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35433\
        );

    \I__7698\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35433\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__35433\,
            I => n3_adj_2485
        );

    \I__7696\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__35427\,
            I => \N__35424\
        );

    \I__7694\ : Odrv4
    port map (
            O => \N__35424\,
            I => n6
        );

    \I__7693\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35415\
        );

    \I__7692\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35415\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__35415\,
            I => n17349
        );

    \I__7690\ : CascadeMux
    port map (
            O => \N__35412\,
            I => \n3_adj_2485_cascade_\
        );

    \I__7689\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35406\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__35406\,
            I => \N__35402\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__35405\,
            I => \N__35398\
        );

    \I__7686\ : Span4Mux_h
    port map (
            O => \N__35402\,
            I => \N__35395\
        );

    \I__7685\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35390\
        );

    \I__7684\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35390\
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__35395\,
            I => data_in_2_1
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__35390\,
            I => data_in_2_1
        );

    \I__7681\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35381\
        );

    \I__7680\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35378\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__35381\,
            I => \N__35374\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__35378\,
            I => \N__35371\
        );

    \I__7677\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35367\
        );

    \I__7676\ : Span4Mux_v
    port map (
            O => \N__35374\,
            I => \N__35364\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__35371\,
            I => \N__35361\
        );

    \I__7674\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35358\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__35367\,
            I => \N__35353\
        );

    \I__7672\ : Span4Mux_v
    port map (
            O => \N__35364\,
            I => \N__35353\
        );

    \I__7671\ : Odrv4
    port map (
            O => \N__35361\,
            I => data_in_1_1
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__35358\,
            I => data_in_1_1
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__35353\,
            I => data_in_1_1
        );

    \I__7668\ : CascadeMux
    port map (
            O => \N__35346\,
            I => \N__35342\
        );

    \I__7667\ : CascadeMux
    port map (
            O => \N__35345\,
            I => \N__35339\
        );

    \I__7666\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35336\
        );

    \I__7665\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35333\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__35336\,
            I => \N__35330\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__35333\,
            I => \c0.data_in_frame_3_5\
        );

    \I__7662\ : Odrv12
    port map (
            O => \N__35330\,
            I => \c0.data_in_frame_3_5\
        );

    \I__7661\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35321\
        );

    \I__7660\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35318\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35314\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__35318\,
            I => \N__35311\
        );

    \I__7657\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35308\
        );

    \I__7656\ : Sp12to4
    port map (
            O => \N__35314\,
            I => \N__35303\
        );

    \I__7655\ : Sp12to4
    port map (
            O => \N__35311\,
            I => \N__35303\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__35308\,
            I => \c0.data_in_frame_2_3\
        );

    \I__7653\ : Odrv12
    port map (
            O => \N__35303\,
            I => \c0.data_in_frame_2_3\
        );

    \I__7652\ : CascadeMux
    port map (
            O => \N__35298\,
            I => \N__35294\
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__35297\,
            I => \N__35289\
        );

    \I__7650\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35284\
        );

    \I__7649\ : InMux
    port map (
            O => \N__35293\,
            I => \N__35281\
        );

    \I__7648\ : CascadeMux
    port map (
            O => \N__35292\,
            I => \N__35278\
        );

    \I__7647\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35269\
        );

    \I__7646\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35269\
        );

    \I__7645\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35269\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__35284\,
            I => \N__35264\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__35281\,
            I => \N__35264\
        );

    \I__7642\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35261\
        );

    \I__7641\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35258\
        );

    \I__7640\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35255\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__35269\,
            I => \N__35250\
        );

    \I__7638\ : Span4Mux_v
    port map (
            O => \N__35264\,
            I => \N__35250\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__35261\,
            I => rx_data_3
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__35258\,
            I => rx_data_3
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__35255\,
            I => rx_data_3
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__35250\,
            I => rx_data_3
        );

    \I__7633\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35238\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__35238\,
            I => \N__35234\
        );

    \I__7631\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35230\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__35234\,
            I => \N__35227\
        );

    \I__7629\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35224\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__35230\,
            I => \N__35221\
        );

    \I__7627\ : Odrv4
    port map (
            O => \N__35227\,
            I => data_in_3_3
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__35224\,
            I => data_in_3_3
        );

    \I__7625\ : Odrv12
    port map (
            O => \N__35221\,
            I => data_in_3_3
        );

    \I__7624\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35207\
        );

    \I__7622\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35204\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__35207\,
            I => \N__35201\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__35204\,
            I => \N__35197\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__35201\,
            I => \N__35194\
        );

    \I__7618\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35191\
        );

    \I__7617\ : Span12Mux_h
    port map (
            O => \N__35197\,
            I => \N__35188\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__35194\,
            I => \N__35185\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__35191\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__7614\ : Odrv12
    port map (
            O => \N__35188\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__35185\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__7612\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35175\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__35175\,
            I => \N__35172\
        );

    \I__7610\ : Span4Mux_h
    port map (
            O => \N__35172\,
            I => \N__35169\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__35169\,
            I => \c0.n50\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__35166\,
            I => \c0.n47_cascade_\
        );

    \I__7607\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35160\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__35160\,
            I => \c0.n49\
        );

    \I__7605\ : InMux
    port map (
            O => \N__35157\,
            I => \N__35154\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__35154\,
            I => \N__35151\
        );

    \I__7603\ : Span12Mux_h
    port map (
            O => \N__35151\,
            I => \N__35148\
        );

    \I__7602\ : Odrv12
    port map (
            O => \N__35148\,
            I => \c0.n51\
        );

    \I__7601\ : CascadeMux
    port map (
            O => \N__35145\,
            I => \c0.n56_cascade_\
        );

    \I__7600\ : InMux
    port map (
            O => \N__35142\,
            I => \N__35139\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35136\
        );

    \I__7598\ : Span4Mux_h
    port map (
            O => \N__35136\,
            I => \N__35133\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__35133\,
            I => \c0.n45\
        );

    \I__7596\ : CascadeMux
    port map (
            O => \N__35130\,
            I => \c0.n10018_cascade_\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__35127\,
            I => \N__35124\
        );

    \I__7594\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35121\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35116\
        );

    \I__7592\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35113\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__35119\,
            I => \N__35110\
        );

    \I__7590\ : Span4Mux_v
    port map (
            O => \N__35116\,
            I => \N__35105\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__35113\,
            I => \N__35105\
        );

    \I__7588\ : InMux
    port map (
            O => \N__35110\,
            I => \N__35102\
        );

    \I__7587\ : Span4Mux_h
    port map (
            O => \N__35105\,
            I => \N__35099\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__35102\,
            I => \c0.data_in_frame_2_0\
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__35099\,
            I => \c0.data_in_frame_2_0\
        );

    \I__7584\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35089\
        );

    \I__7583\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35084\
        );

    \I__7582\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35084\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__35089\,
            I => \N__35081\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__35084\,
            I => \N__35078\
        );

    \I__7579\ : Span4Mux_h
    port map (
            O => \N__35081\,
            I => \N__35075\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__35078\,
            I => \N__35071\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__35075\,
            I => \N__35068\
        );

    \I__7576\ : InMux
    port map (
            O => \N__35074\,
            I => \N__35065\
        );

    \I__7575\ : Span4Mux_v
    port map (
            O => \N__35071\,
            I => \N__35062\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__35068\,
            I => data_in_3_6
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__35065\,
            I => data_in_3_6
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__35062\,
            I => data_in_3_6
        );

    \I__7571\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35052\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__35052\,
            I => \N__35047\
        );

    \I__7569\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35044\
        );

    \I__7568\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35041\
        );

    \I__7567\ : Odrv12
    port map (
            O => \N__35047\,
            I => data_in_1_0
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__35044\,
            I => data_in_1_0
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__35041\,
            I => data_in_1_0
        );

    \I__7564\ : InMux
    port map (
            O => \N__35034\,
            I => \N__35031\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35027\
        );

    \I__7562\ : InMux
    port map (
            O => \N__35030\,
            I => \N__35023\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__35027\,
            I => \N__35020\
        );

    \I__7560\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35017\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__35023\,
            I => data_in_0_0
        );

    \I__7558\ : Odrv4
    port map (
            O => \N__35020\,
            I => data_in_0_0
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__35017\,
            I => data_in_0_0
        );

    \I__7556\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35006\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__35009\,
            I => \N__35003\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__35006\,
            I => \N__35000\
        );

    \I__7553\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34996\
        );

    \I__7552\ : Span4Mux_h
    port map (
            O => \N__35000\,
            I => \N__34993\
        );

    \I__7551\ : InMux
    port map (
            O => \N__34999\,
            I => \N__34990\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34987\
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__34993\,
            I => data_in_3_1
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__34990\,
            I => data_in_3_1
        );

    \I__7547\ : Odrv12
    port map (
            O => \N__34987\,
            I => data_in_3_1
        );

    \I__7546\ : InMux
    port map (
            O => \N__34980\,
            I => \N__34977\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__34977\,
            I => \c0.n2128\
        );

    \I__7544\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34970\
        );

    \I__7543\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34967\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__34970\,
            I => \N__34962\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34962\
        );

    \I__7540\ : Odrv4
    port map (
            O => \N__34962\,
            I => data_in_frame_6_7
        );

    \I__7539\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34955\
        );

    \I__7538\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34952\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__34955\,
            I => \c0.data_in_frame_5_0\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__34952\,
            I => \c0.data_in_frame_5_0\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__34947\,
            I => \c0.n2128_cascade_\
        );

    \I__7534\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34941\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__34941\,
            I => \N__34938\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__34938\,
            I => \c0.n19_adj_2324\
        );

    \I__7531\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34930\
        );

    \I__7530\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34927\
        );

    \I__7529\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34924\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34920\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34917\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__34924\,
            I => \N__34914\
        );

    \I__7525\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34911\
        );

    \I__7524\ : Span12Mux_s11_h
    port map (
            O => \N__34920\,
            I => \N__34908\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__34917\,
            I => \N__34903\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__34914\,
            I => \N__34903\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__34911\,
            I => data_in_3_0
        );

    \I__7520\ : Odrv12
    port map (
            O => \N__34908\,
            I => data_in_3_0
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__34903\,
            I => data_in_3_0
        );

    \I__7518\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34891\
        );

    \I__7517\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34887\
        );

    \I__7516\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34884\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__34891\,
            I => \N__34881\
        );

    \I__7514\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34878\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__34887\,
            I => \c0.data_in_frame_0_3\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__34884\,
            I => \c0.data_in_frame_0_3\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__34881\,
            I => \c0.data_in_frame_0_3\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__34878\,
            I => \c0.data_in_frame_0_3\
        );

    \I__7509\ : CascadeMux
    port map (
            O => \N__34869\,
            I => \N__34866\
        );

    \I__7508\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34862\
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__34865\,
            I => \N__34859\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__34862\,
            I => \N__34856\
        );

    \I__7505\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34851\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__34856\,
            I => \N__34848\
        );

    \I__7503\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34845\
        );

    \I__7502\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34842\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__34851\,
            I => \c0.data_in_frame_0_2\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__34848\,
            I => \c0.data_in_frame_0_2\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__34845\,
            I => \c0.data_in_frame_0_2\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__34842\,
            I => \c0.data_in_frame_0_2\
        );

    \I__7497\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34829\
        );

    \I__7496\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34826\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__34829\,
            I => \N__34821\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34821\
        );

    \I__7493\ : Span4Mux_v
    port map (
            O => \N__34821\,
            I => \N__34817\
        );

    \I__7492\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34814\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__34817\,
            I => \c0.n2120\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__34814\,
            I => \c0.n2120\
        );

    \I__7489\ : CascadeMux
    port map (
            O => \N__34809\,
            I => \c0.n22_adj_2201_cascade_\
        );

    \I__7488\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34803\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__34803\,
            I => \c0.n27_adj_2202\
        );

    \I__7486\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34793\
        );

    \I__7485\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34790\
        );

    \I__7484\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34785\
        );

    \I__7483\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34785\
        );

    \I__7482\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34782\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__34793\,
            I => \c0.data_in_frame_0_5\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__34790\,
            I => \c0.data_in_frame_0_5\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__34785\,
            I => \c0.data_in_frame_0_5\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__34782\,
            I => \c0.data_in_frame_0_5\
        );

    \I__7477\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34768\
        );

    \I__7476\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34760\
        );

    \I__7475\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34757\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34754\
        );

    \I__7473\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34751\
        );

    \I__7472\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34744\
        );

    \I__7471\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34744\
        );

    \I__7470\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34744\
        );

    \I__7469\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34741\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__34760\,
            I => \c0.data_in_frame_0_6\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__34757\,
            I => \c0.data_in_frame_0_6\
        );

    \I__7466\ : Odrv12
    port map (
            O => \N__34754\,
            I => \c0.data_in_frame_0_6\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__34751\,
            I => \c0.data_in_frame_0_6\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__34744\,
            I => \c0.data_in_frame_0_6\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__34741\,
            I => \c0.data_in_frame_0_6\
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__34728\,
            I => \c0.n17469_cascade_\
        );

    \I__7461\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34721\
        );

    \I__7460\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34718\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34715\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__34718\,
            I => \N__34711\
        );

    \I__7457\ : Span4Mux_h
    port map (
            O => \N__34715\,
            I => \N__34707\
        );

    \I__7456\ : CascadeMux
    port map (
            O => \N__34714\,
            I => \N__34704\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__34711\,
            I => \N__34701\
        );

    \I__7454\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34698\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__34707\,
            I => \N__34695\
        );

    \I__7452\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34692\
        );

    \I__7451\ : Sp12to4
    port map (
            O => \N__34701\,
            I => \N__34687\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__34698\,
            I => \N__34687\
        );

    \I__7449\ : Odrv4
    port map (
            O => \N__34695\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__34692\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__7447\ : Odrv12
    port map (
            O => \N__34687\,
            I => \c0.data_out_frame2_0_7\
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__7445\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34674\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34670\
        );

    \I__7443\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34667\
        );

    \I__7442\ : Span4Mux_h
    port map (
            O => \N__34670\,
            I => \N__34664\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__34667\,
            I => data_in_frame_6_1
        );

    \I__7440\ : Odrv4
    port map (
            O => \N__34664\,
            I => data_in_frame_6_1
        );

    \I__7439\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34656\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__34656\,
            I => \N__34652\
        );

    \I__7437\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34649\
        );

    \I__7436\ : Span4Mux_h
    port map (
            O => \N__34652\,
            I => \N__34646\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__34649\,
            I => \c0.data_in_frame_5_1\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__34646\,
            I => \c0.data_in_frame_5_1\
        );

    \I__7433\ : CascadeMux
    port map (
            O => \N__34641\,
            I => \c0.n17114_cascade_\
        );

    \I__7432\ : CascadeMux
    port map (
            O => \N__34638\,
            I => \N__34635\
        );

    \I__7431\ : InMux
    port map (
            O => \N__34635\,
            I => \N__34632\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__34632\,
            I => \N__34629\
        );

    \I__7429\ : Span4Mux_h
    port map (
            O => \N__34629\,
            I => \N__34625\
        );

    \I__7428\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34622\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__34625\,
            I => \N__34619\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__34622\,
            I => \c0.data_in_frame_5_7\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__34619\,
            I => \c0.data_in_frame_5_7\
        );

    \I__7424\ : CascadeMux
    port map (
            O => \N__34614\,
            I => \N__34610\
        );

    \I__7423\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34604\
        );

    \I__7422\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34601\
        );

    \I__7421\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34596\
        );

    \I__7420\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34596\
        );

    \I__7419\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34593\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34590\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__34601\,
            I => \c0.data_in_frame_1_4\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__34596\,
            I => \c0.data_in_frame_1_4\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__34593\,
            I => \c0.data_in_frame_1_4\
        );

    \I__7414\ : Odrv4
    port map (
            O => \N__34590\,
            I => \c0.data_in_frame_1_4\
        );

    \I__7413\ : CascadeMux
    port map (
            O => \N__34581\,
            I => \c0.n17101_cascade_\
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__34578\,
            I => \c0.n10_adj_2299_cascade_\
        );

    \I__7411\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34571\
        );

    \I__7410\ : InMux
    port map (
            O => \N__34574\,
            I => \N__34568\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__34571\,
            I => \c0.n17206\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__34568\,
            I => \c0.n17206\
        );

    \I__7407\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34557\
        );

    \I__7406\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34557\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__34557\,
            I => \c0.n10407\
        );

    \I__7404\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34551\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__34551\,
            I => \N__34547\
        );

    \I__7402\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34544\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__34547\,
            I => \N__34541\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34536\
        );

    \I__7399\ : Span4Mux_h
    port map (
            O => \N__34541\,
            I => \N__34536\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__34536\,
            I => data_in_frame_6_0
        );

    \I__7397\ : CascadeMux
    port map (
            O => \N__34533\,
            I => \c0.n10407_cascade_\
        );

    \I__7396\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34523\
        );

    \I__7395\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34523\
        );

    \I__7394\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34518\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__34523\,
            I => \N__34515\
        );

    \I__7392\ : CascadeMux
    port map (
            O => \N__34522\,
            I => \N__34512\
        );

    \I__7391\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34509\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34506\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__34515\,
            I => \N__34503\
        );

    \I__7388\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34500\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__34509\,
            I => \c0.data_in_frame_1_5\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__34506\,
            I => \c0.data_in_frame_1_5\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__34503\,
            I => \c0.data_in_frame_1_5\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__34500\,
            I => \c0.data_in_frame_1_5\
        );

    \I__7383\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34488\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__34488\,
            I => \c0.n17215\
        );

    \I__7381\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34481\
        );

    \I__7380\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34478\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__34481\,
            I => \N__34471\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__34478\,
            I => \N__34471\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__34477\,
            I => \N__34468\
        );

    \I__7376\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34465\
        );

    \I__7375\ : Span4Mux_h
    port map (
            O => \N__34471\,
            I => \N__34462\
        );

    \I__7374\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34459\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__34465\,
            I => \N__34456\
        );

    \I__7372\ : Span4Mux_h
    port map (
            O => \N__34462\,
            I => \N__34453\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__34459\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__7370\ : Odrv12
    port map (
            O => \N__34456\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__7369\ : Odrv4
    port map (
            O => \N__34453\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__7368\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__34443\,
            I => \N__34438\
        );

    \I__7366\ : InMux
    port map (
            O => \N__34442\,
            I => \N__34434\
        );

    \I__7365\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34431\
        );

    \I__7364\ : Span4Mux_h
    port map (
            O => \N__34438\,
            I => \N__34428\
        );

    \I__7363\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34425\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__34434\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__34431\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__34428\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__34425\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__7358\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34413\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__34413\,
            I => \c0.n13284\
        );

    \I__7356\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34404\
        );

    \I__7355\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34404\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__34404\,
            I => \c0.n13628\
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__34401\,
            I => \c0.n13628_cascade_\
        );

    \I__7352\ : InMux
    port map (
            O => \N__34398\,
            I => \N__34392\
        );

    \I__7351\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34387\
        );

    \I__7350\ : InMux
    port map (
            O => \N__34396\,
            I => \N__34387\
        );

    \I__7349\ : CascadeMux
    port map (
            O => \N__34395\,
            I => \N__34384\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34379\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34379\
        );

    \I__7346\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34376\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__34379\,
            I => \N__34373\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__34376\,
            I => tx2_active
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__34373\,
            I => tx2_active
        );

    \I__7342\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34365\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__34365\,
            I => \N__34361\
        );

    \I__7340\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34358\
        );

    \I__7339\ : Span4Mux_h
    port map (
            O => \N__34361\,
            I => \N__34355\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__34358\,
            I => \c0.data_in_frame_3_2\
        );

    \I__7337\ : Odrv4
    port map (
            O => \N__34355\,
            I => \c0.data_in_frame_3_2\
        );

    \I__7336\ : CascadeMux
    port map (
            O => \N__34350\,
            I => \N__34347\
        );

    \I__7335\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34344\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__34344\,
            I => \N__34340\
        );

    \I__7333\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34337\
        );

    \I__7332\ : Span4Mux_v
    port map (
            O => \N__34340\,
            I => \N__34334\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__34337\,
            I => data_in_frame_6_2
        );

    \I__7330\ : Odrv4
    port map (
            O => \N__34334\,
            I => data_in_frame_6_2
        );

    \I__7329\ : CascadeMux
    port map (
            O => \N__34329\,
            I => \c0.n17475_cascade_\
        );

    \I__7328\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34322\
        );

    \I__7327\ : CascadeMux
    port map (
            O => \N__34325\,
            I => \N__34319\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34315\
        );

    \I__7325\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34309\
        );

    \I__7324\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34309\
        );

    \I__7323\ : Span4Mux_h
    port map (
            O => \N__34315\,
            I => \N__34306\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__34314\,
            I => \N__34303\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__34309\,
            I => \N__34300\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__34306\,
            I => \N__34297\
        );

    \I__7319\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34294\
        );

    \I__7318\ : Span12Mux_s4_h
    port map (
            O => \N__34300\,
            I => \N__34291\
        );

    \I__7317\ : Span4Mux_h
    port map (
            O => \N__34297\,
            I => \N__34288\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__34294\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__7315\ : Odrv12
    port map (
            O => \N__34291\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__7314\ : Odrv4
    port map (
            O => \N__34288\,
            I => \c0.data_out_frame2_0_5\
        );

    \I__7313\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34278\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__34278\,
            I => \N__34275\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__34275\,
            I => \N__34272\
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__34272\,
            I => \c0.n16352\
        );

    \I__7309\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34266\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__34266\,
            I => \c0.n24_adj_2340\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__34263\,
            I => \N__34260\
        );

    \I__7306\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34257\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__34257\,
            I => \N__34254\
        );

    \I__7304\ : Span4Mux_h
    port map (
            O => \N__34254\,
            I => \N__34250\
        );

    \I__7303\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34247\
        );

    \I__7302\ : Sp12to4
    port map (
            O => \N__34250\,
            I => \N__34244\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__34247\,
            I => data_in_frame_6_5
        );

    \I__7300\ : Odrv12
    port map (
            O => \N__34244\,
            I => data_in_frame_6_5
        );

    \I__7299\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34233\
        );

    \I__7298\ : InMux
    port map (
            O => \N__34238\,
            I => \N__34233\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__34233\,
            I => \N__34230\
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__34230\,
            I => \c0.n2122\
        );

    \I__7295\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34223\
        );

    \I__7294\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34220\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__34223\,
            I => data_out_0_5
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__34220\,
            I => data_out_0_5
        );

    \I__7291\ : InMux
    port map (
            O => \N__34215\,
            I => \N__34211\
        );

    \I__7290\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34208\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__34211\,
            I => data_out_2_2
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__34208\,
            I => data_out_2_2
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__34203\,
            I => \n2699_cascade_\
        );

    \I__7286\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34196\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34193\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__34196\,
            I => \N__34190\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__34193\,
            I => data_out_3_4
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__34190\,
            I => data_out_3_4
        );

    \I__7281\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34176\
        );

    \I__7280\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34176\
        );

    \I__7279\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34176\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__34176\,
            I => n2699
        );

    \I__7277\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34169\
        );

    \I__7276\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34166\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__34169\,
            I => data_out_3_2
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__34166\,
            I => data_out_3_2
        );

    \I__7273\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34157\
        );

    \I__7272\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34154\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__34157\,
            I => \N__34150\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__34154\,
            I => \N__34147\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34144\
        );

    \I__7268\ : Span4Mux_v
    port map (
            O => \N__34150\,
            I => \N__34141\
        );

    \I__7267\ : Span4Mux_h
    port map (
            O => \N__34147\,
            I => \N__34138\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__34144\,
            I => \c0.data_in_frame_2_6\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__34141\,
            I => \c0.data_in_frame_2_6\
        );

    \I__7264\ : Odrv4
    port map (
            O => \N__34138\,
            I => \c0.data_in_frame_2_6\
        );

    \I__7263\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__34128\,
            I => \N__34125\
        );

    \I__7261\ : Span4Mux_h
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__34122\,
            I => \c0.n17713\
        );

    \I__7259\ : SRMux
    port map (
            O => \N__34119\,
            I => \N__34116\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__34116\,
            I => \c0.n4_adj_2325\
        );

    \I__7257\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34099\
        );

    \I__7256\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34099\
        );

    \I__7255\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34099\
        );

    \I__7254\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34088\
        );

    \I__7253\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34088\
        );

    \I__7252\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34088\
        );

    \I__7251\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34088\
        );

    \I__7250\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34088\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34083\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__34088\,
            I => \N__34083\
        );

    \I__7247\ : Odrv12
    port map (
            O => \N__34083\,
            I => \c0.tx2_transmit_N_1996\
        );

    \I__7246\ : InMux
    port map (
            O => \N__34080\,
            I => \N__34077\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__34077\,
            I => \c0.n17676\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__34074\,
            I => \N__34071\
        );

    \I__7243\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34068\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__34068\,
            I => \N__34064\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__34067\,
            I => \N__34061\
        );

    \I__7240\ : Span4Mux_v
    port map (
            O => \N__34064\,
            I => \N__34058\
        );

    \I__7239\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34055\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__34058\,
            I => rand_setpoint_14
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__34055\,
            I => rand_setpoint_14
        );

    \I__7236\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34047\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__34047\,
            I => \c0.n17703\
        );

    \I__7234\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34038\
        );

    \I__7233\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34038\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__34038\,
            I => \c0.data_out_1_4\
        );

    \I__7231\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34032\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__34032\,
            I => \c0.n17675\
        );

    \I__7229\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34026\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__34026\,
            I => \N__34023\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__34023\,
            I => \c0.n17697\
        );

    \I__7226\ : InMux
    port map (
            O => \N__34020\,
            I => \N__34017\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__34017\,
            I => \N__34014\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__34014\,
            I => n18271
        );

    \I__7223\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \n10_adj_2408_cascade_\
        );

    \I__7222\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34002\
        );

    \I__7221\ : InMux
    port map (
            O => \N__34007\,
            I => \N__34002\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__34002\,
            I => \c0.data_out_2_3\
        );

    \I__7219\ : CascadeMux
    port map (
            O => \N__33999\,
            I => \c0.n18268_cascade_\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__33996\,
            I => \c0.tx.n55_cascade_\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__33993\,
            I => \N__33990\
        );

    \I__7216\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33987\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__33987\,
            I => \c0.n5_adj_2136\
        );

    \I__7214\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33980\
        );

    \I__7213\ : CascadeMux
    port map (
            O => \N__33983\,
            I => \N__33977\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__33980\,
            I => \N__33974\
        );

    \I__7211\ : InMux
    port map (
            O => \N__33977\,
            I => \N__33971\
        );

    \I__7210\ : Odrv4
    port map (
            O => \N__33974\,
            I => rand_setpoint_12
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__33971\,
            I => rand_setpoint_12
        );

    \I__7208\ : CascadeMux
    port map (
            O => \N__33966\,
            I => \N__33963\
        );

    \I__7207\ : InMux
    port map (
            O => \N__33963\,
            I => \N__33960\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__33960\,
            I => \c0.n5\
        );

    \I__7205\ : CascadeMux
    port map (
            O => \N__33957\,
            I => \c0.n18172_cascade_\
        );

    \I__7204\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33951\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__33951\,
            I => \c0.n17764\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__33948\,
            I => \c0.n17639_cascade_\
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__33945\,
            I => \N__33941\
        );

    \I__7200\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33938\
        );

    \I__7199\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33935\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__33938\,
            I => rand_setpoint_20
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__33935\,
            I => rand_setpoint_20
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__33930\,
            I => \N__33926\
        );

    \I__7195\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33923\
        );

    \I__7194\ : InMux
    port map (
            O => \N__33926\,
            I => \N__33920\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__33923\,
            I => rand_setpoint_22
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__33920\,
            I => rand_setpoint_22
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__7190\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33909\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__33909\,
            I => \N__33906\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__33903\,
            I => \c0.n17647\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__33900\,
            I => \N__33896\
        );

    \I__7185\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33893\
        );

    \I__7184\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33890\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__33893\,
            I => rand_setpoint_19
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__33890\,
            I => rand_setpoint_19
        );

    \I__7181\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \c0.n17631_cascade_\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__33882\,
            I => \N__33878\
        );

    \I__7179\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33875\
        );

    \I__7178\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33872\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__33875\,
            I => rand_setpoint_18
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__33872\,
            I => rand_setpoint_18
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__33867\,
            I => \c0.n17627_cascade_\
        );

    \I__7174\ : CascadeMux
    port map (
            O => \N__33864\,
            I => \N__33860\
        );

    \I__7173\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33857\
        );

    \I__7172\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33854\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__33857\,
            I => rand_setpoint_21
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__33854\,
            I => rand_setpoint_21
        );

    \I__7169\ : CascadeMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__7168\ : InMux
    port map (
            O => \N__33846\,
            I => \N__33843\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__33843\,
            I => \N__33840\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__7165\ : Span4Mux_h
    port map (
            O => \N__33837\,
            I => \N__33834\
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__33834\,
            I => \c0.n17643\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__33831\,
            I => \N__33827\
        );

    \I__7162\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33824\
        );

    \I__7161\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33821\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__33824\,
            I => rand_setpoint_2
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__33821\,
            I => rand_setpoint_2
        );

    \I__7158\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33812\
        );

    \I__7157\ : CascadeMux
    port map (
            O => \N__33815\,
            I => \N__33809\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__33812\,
            I => \N__33806\
        );

    \I__7155\ : InMux
    port map (
            O => \N__33809\,
            I => \N__33803\
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__33806\,
            I => rand_setpoint_3
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__33803\,
            I => rand_setpoint_3
        );

    \I__7152\ : CascadeMux
    port map (
            O => \N__33798\,
            I => \N__33795\
        );

    \I__7151\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33790\
        );

    \I__7150\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33787\
        );

    \I__7149\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33784\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__33790\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__33787\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__33784\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__7145\ : SRMux
    port map (
            O => \N__33777\,
            I => \N__33774\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33771\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__33771\,
            I => \N__33768\
        );

    \I__7142\ : Odrv4
    port map (
            O => \N__33768\,
            I => \c0.n16141\
        );

    \I__7141\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33761\
        );

    \I__7140\ : CascadeMux
    port map (
            O => \N__33764\,
            I => \N__33758\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__33761\,
            I => \N__33755\
        );

    \I__7138\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33752\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__33755\,
            I => rand_setpoint_23
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__33752\,
            I => rand_setpoint_23
        );

    \I__7135\ : CascadeMux
    port map (
            O => \N__33747\,
            I => \n21_adj_2487_cascade_\
        );

    \I__7134\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33736\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__33740\,
            I => \N__33733\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__33739\,
            I => \N__33729\
        );

    \I__7130\ : Span4Mux_v
    port map (
            O => \N__33736\,
            I => \N__33725\
        );

    \I__7129\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33720\
        );

    \I__7128\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33720\
        );

    \I__7127\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33715\
        );

    \I__7126\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33715\
        );

    \I__7125\ : Odrv4
    port map (
            O => \N__33725\,
            I => n63_adj_2418
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__33720\,
            I => n63_adj_2418
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__33715\,
            I => n63_adj_2418
        );

    \I__7122\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33705\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__33705\,
            I => n6_adj_2410
        );

    \I__7120\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33699\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__33699\,
            I => \N__33695\
        );

    \I__7118\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33692\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__33695\,
            I => n2061
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__33692\,
            I => n2061
        );

    \I__7115\ : CascadeMux
    port map (
            O => \N__33687\,
            I => \N__33684\
        );

    \I__7114\ : InMux
    port map (
            O => \N__33684\,
            I => \N__33681\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__33681\,
            I => \N__33678\
        );

    \I__7112\ : Span4Mux_h
    port map (
            O => \N__33678\,
            I => \N__33675\
        );

    \I__7111\ : Span4Mux_h
    port map (
            O => \N__33675\,
            I => \N__33672\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__33672\,
            I => \c0.n51_adj_2173\
        );

    \I__7109\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33663\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__33663\,
            I => \N__33660\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__33660\,
            I => \c0.n10166\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__33657\,
            I => \N__33652\
        );

    \I__7104\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33648\
        );

    \I__7103\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33643\
        );

    \I__7102\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33643\
        );

    \I__7101\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33640\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__33648\,
            I => \N__33637\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__33643\,
            I => \N__33634\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__33640\,
            I => \N__33631\
        );

    \I__7097\ : Span12Mux_v
    port map (
            O => \N__33637\,
            I => \N__33628\
        );

    \I__7096\ : Span4Mux_v
    port map (
            O => \N__33634\,
            I => \N__33625\
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__33631\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__7094\ : Odrv12
    port map (
            O => \N__33628\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__7093\ : Odrv4
    port map (
            O => \N__33625\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__7092\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__7090\ : Span4Mux_v
    port map (
            O => \N__33612\,
            I => \N__33609\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__7088\ : Span4Mux_h
    port map (
            O => \N__33606\,
            I => \N__33603\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__33603\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_30\
        );

    \I__7086\ : SRMux
    port map (
            O => \N__33600\,
            I => \N__33597\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33594\
        );

    \I__7084\ : Span4Mux_h
    port map (
            O => \N__33594\,
            I => \N__33591\
        );

    \I__7083\ : Span4Mux_h
    port map (
            O => \N__33591\,
            I => \N__33588\
        );

    \I__7082\ : Odrv4
    port map (
            O => \N__33588\,
            I => \c0.n16696\
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__33585\,
            I => \c0.n8_adj_2385_cascade_\
        );

    \I__7080\ : SRMux
    port map (
            O => \N__33582\,
            I => \N__33579\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__33579\,
            I => \N__33576\
        );

    \I__7078\ : Span4Mux_s2_v
    port map (
            O => \N__33576\,
            I => \N__33573\
        );

    \I__7077\ : Span4Mux_h
    port map (
            O => \N__33573\,
            I => \N__33570\
        );

    \I__7076\ : Span4Mux_h
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__33567\,
            I => \N__33564\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__33564\,
            I => \c0.n16670\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__33561\,
            I => \c0.n17367_cascade_\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__33558\,
            I => \n9_cascade_\
        );

    \I__7071\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33550\
        );

    \I__7070\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33547\
        );

    \I__7069\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33544\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__33550\,
            I => \c0.n10139\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__33547\,
            I => \c0.n10139\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__33544\,
            I => \c0.n10139\
        );

    \I__7065\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33531\
        );

    \I__7064\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33528\
        );

    \I__7063\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33523\
        );

    \I__7062\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33523\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__33531\,
            I => \N__33516\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33511\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33511\
        );

    \I__7058\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33502\
        );

    \I__7057\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33502\
        );

    \I__7056\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33502\
        );

    \I__7055\ : InMux
    port map (
            O => \N__33519\,
            I => \N__33502\
        );

    \I__7054\ : Span4Mux_h
    port map (
            O => \N__33516\,
            I => \N__33499\
        );

    \I__7053\ : Sp12to4
    port map (
            O => \N__33511\,
            I => \N__33494\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33494\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__33499\,
            I => \c0.n11833\
        );

    \I__7050\ : Odrv12
    port map (
            O => \N__33494\,
            I => \c0.n11833\
        );

    \I__7049\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33484\
        );

    \I__7048\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33479\
        );

    \I__7047\ : InMux
    port map (
            O => \N__33487\,
            I => \N__33479\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__33484\,
            I => \N__33476\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__33479\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__7044\ : Odrv4
    port map (
            O => \N__33476\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__7043\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33466\
        );

    \I__7042\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33463\
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__33469\,
            I => \N__33460\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33455\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33455\
        );

    \I__7038\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33452\
        );

    \I__7037\ : Span4Mux_h
    port map (
            O => \N__33455\,
            I => \N__33449\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__33452\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__7035\ : Odrv4
    port map (
            O => \N__33449\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__7034\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33441\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__33441\,
            I => \N__33438\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__33438\,
            I => \N__33433\
        );

    \I__7031\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33430\
        );

    \I__7030\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33427\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__33433\,
            I => \N__33422\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__33430\,
            I => \N__33422\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__33427\,
            I => n9
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__33422\,
            I => n9
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__33417\,
            I => \N__33413\
        );

    \I__7024\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33409\
        );

    \I__7023\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33406\
        );

    \I__7022\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33403\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__33409\,
            I => \N__33400\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__33406\,
            I => \N__33397\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__33403\,
            I => \c0.data_in_frame_2_4\
        );

    \I__7018\ : Odrv12
    port map (
            O => \N__33400\,
            I => \c0.data_in_frame_2_4\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__33397\,
            I => \c0.data_in_frame_2_4\
        );

    \I__7016\ : CascadeMux
    port map (
            O => \N__33390\,
            I => \FRAME_MATCHER_i_31__N_1273_cascade_\
        );

    \I__7015\ : CascadeMux
    port map (
            O => \N__33387\,
            I => \n17086_cascade_\
        );

    \I__7014\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33375\
        );

    \I__7013\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33375\
        );

    \I__7012\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33372\
        );

    \I__7011\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33367\
        );

    \I__7010\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33367\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__33375\,
            I => n63_adj_2428
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__33372\,
            I => n63_adj_2428
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__33367\,
            I => n63_adj_2428
        );

    \I__7006\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33356\
        );

    \I__7005\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33351\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33348\
        );

    \I__7003\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33343\
        );

    \I__7002\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33343\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__33351\,
            I => n63
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__33348\,
            I => n63
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__33343\,
            I => n63
        );

    \I__6998\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33333\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33329\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__33332\,
            I => \N__33326\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__33329\,
            I => \N__33323\
        );

    \I__6994\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33319\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__33323\,
            I => \N__33316\
        );

    \I__6992\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33313\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__33319\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__33316\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__33313\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__6988\ : SRMux
    port map (
            O => \N__33306\,
            I => \N__33303\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__6985\ : Span4Mux_h
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__33294\,
            I => \c0.n16666\
        );

    \I__6983\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33287\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__33290\,
            I => \N__33284\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__33287\,
            I => \N__33281\
        );

    \I__6980\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33277\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__33281\,
            I => \N__33274\
        );

    \I__6978\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33271\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__33277\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__33274\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__33271\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__6974\ : SRMux
    port map (
            O => \N__33264\,
            I => \N__33261\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__33261\,
            I => \N__33258\
        );

    \I__6972\ : Span4Mux_h
    port map (
            O => \N__33258\,
            I => \N__33255\
        );

    \I__6971\ : Odrv4
    port map (
            O => \N__33255\,
            I => \c0.n16674\
        );

    \I__6970\ : InMux
    port map (
            O => \N__33252\,
            I => \N__33243\
        );

    \I__6969\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33240\
        );

    \I__6968\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33237\
        );

    \I__6967\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33229\
        );

    \I__6966\ : InMux
    port map (
            O => \N__33248\,
            I => \N__33226\
        );

    \I__6965\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33215\
        );

    \I__6964\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33212\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33207\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__33240\,
            I => \N__33207\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__33237\,
            I => \N__33204\
        );

    \I__6960\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33201\
        );

    \I__6959\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33198\
        );

    \I__6958\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33194\
        );

    \I__6957\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33191\
        );

    \I__6956\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33188\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__33229\,
            I => \N__33179\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__33226\,
            I => \N__33179\
        );

    \I__6953\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33176\
        );

    \I__6952\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33173\
        );

    \I__6951\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33170\
        );

    \I__6950\ : InMux
    port map (
            O => \N__33222\,
            I => \N__33167\
        );

    \I__6949\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33164\
        );

    \I__6948\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33161\
        );

    \I__6947\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33156\
        );

    \I__6946\ : InMux
    port map (
            O => \N__33218\,
            I => \N__33153\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__33215\,
            I => \N__33143\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__33212\,
            I => \N__33143\
        );

    \I__6943\ : Span4Mux_h
    port map (
            O => \N__33207\,
            I => \N__33134\
        );

    \I__6942\ : Span4Mux_s2_v
    port map (
            O => \N__33204\,
            I => \N__33134\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33134\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__33198\,
            I => \N__33134\
        );

    \I__6939\ : InMux
    port map (
            O => \N__33197\,
            I => \N__33131\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33124\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33124\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__33188\,
            I => \N__33124\
        );

    \I__6935\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33121\
        );

    \I__6934\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33118\
        );

    \I__6933\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33115\
        );

    \I__6932\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33112\
        );

    \I__6931\ : Span4Mux_s3_v
    port map (
            O => \N__33179\,
            I => \N__33099\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__33176\,
            I => \N__33099\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__33173\,
            I => \N__33099\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__33170\,
            I => \N__33099\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__33167\,
            I => \N__33099\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__33164\,
            I => \N__33099\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__33161\,
            I => \N__33096\
        );

    \I__6924\ : InMux
    port map (
            O => \N__33160\,
            I => \N__33093\
        );

    \I__6923\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33090\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33085\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__33153\,
            I => \N__33085\
        );

    \I__6920\ : InMux
    port map (
            O => \N__33152\,
            I => \N__33082\
        );

    \I__6919\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33079\
        );

    \I__6918\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33076\
        );

    \I__6917\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33073\
        );

    \I__6916\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33070\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__33143\,
            I => \N__33063\
        );

    \I__6914\ : Span4Mux_v
    port map (
            O => \N__33134\,
            I => \N__33063\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__33131\,
            I => \N__33063\
        );

    \I__6912\ : Span4Mux_s3_v
    port map (
            O => \N__33124\,
            I => \N__33052\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33052\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33052\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__33115\,
            I => \N__33052\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33052\
        );

    \I__6907\ : Span4Mux_v
    port map (
            O => \N__33099\,
            I => \N__33045\
        );

    \I__6906\ : Span4Mux_s2_h
    port map (
            O => \N__33096\,
            I => \N__33045\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__33093\,
            I => \N__33045\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__33090\,
            I => \N__33040\
        );

    \I__6903\ : Span4Mux_h
    port map (
            O => \N__33085\,
            I => \N__33040\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__33082\,
            I => \N__33028\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__33079\,
            I => \N__33028\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33028\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__33073\,
            I => \N__33028\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33028\
        );

    \I__6897\ : Span4Mux_v
    port map (
            O => \N__33063\,
            I => \N__33025\
        );

    \I__6896\ : Span4Mux_v
    port map (
            O => \N__33052\,
            I => \N__33020\
        );

    \I__6895\ : Span4Mux_h
    port map (
            O => \N__33045\,
            I => \N__33020\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__33040\,
            I => \N__33017\
        );

    \I__6893\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33014\
        );

    \I__6892\ : Span12Mux_s10_v
    port map (
            O => \N__33028\,
            I => \N__33008\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__33025\,
            I => \N__33005\
        );

    \I__6890\ : Span4Mux_h
    port map (
            O => \N__33020\,
            I => \N__33002\
        );

    \I__6889\ : Span4Mux_v
    port map (
            O => \N__33017\,
            I => \N__32999\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__33014\,
            I => \N__32996\
        );

    \I__6887\ : InMux
    port map (
            O => \N__33013\,
            I => \N__32993\
        );

    \I__6886\ : InMux
    port map (
            O => \N__33012\,
            I => \N__32990\
        );

    \I__6885\ : InMux
    port map (
            O => \N__33011\,
            I => \N__32987\
        );

    \I__6884\ : Odrv12
    port map (
            O => \N__33008\,
            I => \c0.n1034\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__33005\,
            I => \c0.n1034\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__33002\,
            I => \c0.n1034\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__32999\,
            I => \c0.n1034\
        );

    \I__6880\ : Odrv12
    port map (
            O => \N__32996\,
            I => \c0.n1034\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__32993\,
            I => \c0.n1034\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__32990\,
            I => \c0.n1034\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__32987\,
            I => \c0.n1034\
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__32970\,
            I => \n10140_cascade_\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \c0.n23_cascade_\
        );

    \I__6874\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32961\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__32961\,
            I => \c0.n26_adj_2210\
        );

    \I__6872\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32955\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__32955\,
            I => \c0.n18\
        );

    \I__6870\ : CascadeMux
    port map (
            O => \N__32952\,
            I => \c0.n30_adj_2213_cascade_\
        );

    \I__6869\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32946\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__32946\,
            I => \N__32943\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__32943\,
            I => \c0.n17_adj_2214\
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__32940\,
            I => \n31_adj_2415_cascade_\
        );

    \I__6865\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32933\
        );

    \I__6864\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32930\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__32933\,
            I => \N__32927\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__32930\,
            I => data_in_frame_6_3
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__32927\,
            I => data_in_frame_6_3
        );

    \I__6860\ : InMux
    port map (
            O => \N__32922\,
            I => \N__32917\
        );

    \I__6859\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32911\
        );

    \I__6858\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32911\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32908\
        );

    \I__6856\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32905\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__32911\,
            I => data_in_3_7
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__32908\,
            I => data_in_3_7
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__32905\,
            I => data_in_3_7
        );

    \I__6852\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32895\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__32895\,
            I => \c0.n6_adj_2358\
        );

    \I__6850\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32889\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32885\
        );

    \I__6848\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32881\
        );

    \I__6847\ : Span4Mux_v
    port map (
            O => \N__32885\,
            I => \N__32877\
        );

    \I__6846\ : CascadeMux
    port map (
            O => \N__32884\,
            I => \N__32874\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32869\
        );

    \I__6844\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32866\
        );

    \I__6843\ : Span4Mux_v
    port map (
            O => \N__32877\,
            I => \N__32862\
        );

    \I__6842\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32857\
        );

    \I__6841\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32857\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__32872\,
            I => \N__32854\
        );

    \I__6839\ : Span4Mux_h
    port map (
            O => \N__32869\,
            I => \N__32849\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__32866\,
            I => \N__32849\
        );

    \I__6837\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32846\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__32862\,
            I => \N__32841\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32841\
        );

    \I__6834\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32838\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__32849\,
            I => \N__32833\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__32846\,
            I => \N__32833\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__32841\,
            I => \N__32830\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__32838\,
            I => \N__32827\
        );

    \I__6829\ : Span4Mux_h
    port map (
            O => \N__32833\,
            I => \N__32824\
        );

    \I__6828\ : Span4Mux_h
    port map (
            O => \N__32830\,
            I => \N__32819\
        );

    \I__6827\ : Span4Mux_v
    port map (
            O => \N__32827\,
            I => \N__32819\
        );

    \I__6826\ : Span4Mux_h
    port map (
            O => \N__32824\,
            I => \N__32816\
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__32819\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__32816\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__32811\,
            I => \N__32807\
        );

    \I__6822\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32804\
        );

    \I__6821\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32801\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32798\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32795\
        );

    \I__6818\ : Span4Mux_v
    port map (
            O => \N__32798\,
            I => \N__32792\
        );

    \I__6817\ : Span4Mux_h
    port map (
            O => \N__32795\,
            I => \N__32788\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__32792\,
            I => \N__32785\
        );

    \I__6815\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32782\
        );

    \I__6814\ : Span4Mux_h
    port map (
            O => \N__32788\,
            I => \N__32779\
        );

    \I__6813\ : Span4Mux_h
    port map (
            O => \N__32785\,
            I => \N__32774\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__32782\,
            I => \N__32774\
        );

    \I__6811\ : Odrv4
    port map (
            O => \N__32779\,
            I => \c0.n15164\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__32774\,
            I => \c0.n15164\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__32769\,
            I => \c0.n17072_cascade_\
        );

    \I__6808\ : InMux
    port map (
            O => \N__32766\,
            I => \N__32762\
        );

    \I__6807\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32759\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__32762\,
            I => \N__32756\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__32759\,
            I => \c0.n10215\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__32756\,
            I => \c0.n10215\
        );

    \I__6803\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32746\
        );

    \I__6802\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32742\
        );

    \I__6801\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32739\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__32746\,
            I => \N__32736\
        );

    \I__6799\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32733\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__32742\,
            I => \c0.data_in_frame_0_4\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__32739\,
            I => \c0.data_in_frame_0_4\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__32736\,
            I => \c0.data_in_frame_0_4\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__32733\,
            I => \c0.data_in_frame_0_4\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__32724\,
            I => \c0.n10215_cascade_\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__32721\,
            I => \c0.n17206_cascade_\
        );

    \I__6792\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32715\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__32712\,
            I => \c0.n20_adj_2195\
        );

    \I__6789\ : CascadeMux
    port map (
            O => \N__32709\,
            I => \N__32703\
        );

    \I__6788\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32697\
        );

    \I__6787\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32697\
        );

    \I__6786\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32692\
        );

    \I__6785\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32687\
        );

    \I__6784\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32687\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__32697\,
            I => \N__32684\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__32696\,
            I => \N__32681\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__32695\,
            I => \N__32677\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__32692\,
            I => \N__32674\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__32687\,
            I => \N__32671\
        );

    \I__6778\ : Span4Mux_h
    port map (
            O => \N__32684\,
            I => \N__32668\
        );

    \I__6777\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32665\
        );

    \I__6776\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32660\
        );

    \I__6775\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32660\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__32674\,
            I => \N__32655\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__32671\,
            I => \N__32655\
        );

    \I__6772\ : Span4Mux_h
    port map (
            O => \N__32668\,
            I => \N__32652\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__32665\,
            I => \N__32647\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32647\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__32655\,
            I => \N__32644\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__32652\,
            I => \N__32641\
        );

    \I__6767\ : Span12Mux_h
    port map (
            O => \N__32647\,
            I => \N__32637\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__32644\,
            I => \N__32634\
        );

    \I__6765\ : Span4Mux_v
    port map (
            O => \N__32641\,
            I => \N__32631\
        );

    \I__6764\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32628\
        );

    \I__6763\ : Odrv12
    port map (
            O => \N__32637\,
            I => \c0.n39\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__32634\,
            I => \c0.n39\
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__32631\,
            I => \c0.n39\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__32628\,
            I => \c0.n39\
        );

    \I__6759\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32615\
        );

    \I__6758\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32612\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__32615\,
            I => \c0.n2137\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__32612\,
            I => \c0.n2137\
        );

    \I__6755\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32604\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__32604\,
            I => \c0.n16475\
        );

    \I__6753\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32597\
        );

    \I__6752\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32594\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__32597\,
            I => \c0.data_in_frame_5_5\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__32594\,
            I => \c0.data_in_frame_5_5\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__32589\,
            I => \N__32586\
        );

    \I__6748\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32583\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__32583\,
            I => \N__32580\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__32580\,
            I => \N__32577\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__32577\,
            I => \c0.n17373\
        );

    \I__6744\ : InMux
    port map (
            O => \N__32574\,
            I => \N__32571\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__32571\,
            I => \c0.n19_adj_2303\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \c0.n17076_cascade_\
        );

    \I__6741\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32556\
        );

    \I__6740\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32553\
        );

    \I__6739\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32546\
        );

    \I__6738\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32546\
        );

    \I__6737\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32546\
        );

    \I__6736\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32541\
        );

    \I__6735\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32541\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__32556\,
            I => n17075
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__32553\,
            I => n17075
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__32546\,
            I => n17075
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__32541\,
            I => n17075
        );

    \I__6730\ : CascadeMux
    port map (
            O => \N__32532\,
            I => \N__32528\
        );

    \I__6729\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32525\
        );

    \I__6728\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32522\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__32525\,
            I => data_in_frame_6_4
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__32522\,
            I => data_in_frame_6_4
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__32517\,
            I => \c0.n2122_cascade_\
        );

    \I__6724\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32511\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__32511\,
            I => \N__32508\
        );

    \I__6722\ : Span4Mux_h
    port map (
            O => \N__32508\,
            I => \N__32503\
        );

    \I__6721\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32498\
        );

    \I__6720\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32498\
        );

    \I__6719\ : Odrv4
    port map (
            O => \N__32503\,
            I => \c0.data_in_frame_2_5\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__32498\,
            I => \c0.data_in_frame_2_5\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__32493\,
            I => \N__32489\
        );

    \I__6716\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32486\
        );

    \I__6715\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32483\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__32486\,
            I => \c0.data_in_frame_5_6\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__32483\,
            I => \c0.data_in_frame_5_6\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__32478\,
            I => \c0.n2124_cascade_\
        );

    \I__6711\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32471\
        );

    \I__6710\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32468\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__32471\,
            I => \c0.data_in_frame_5_3\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__32468\,
            I => \c0.data_in_frame_5_3\
        );

    \I__6707\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32455\
        );

    \I__6706\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32448\
        );

    \I__6705\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32448\
        );

    \I__6704\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32448\
        );

    \I__6703\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32436\
        );

    \I__6702\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32436\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__32455\,
            I => \N__32433\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32430\
        );

    \I__6699\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32425\
        );

    \I__6698\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32425\
        );

    \I__6697\ : InMux
    port map (
            O => \N__32445\,
            I => \N__32418\
        );

    \I__6696\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32418\
        );

    \I__6695\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32405\
        );

    \I__6694\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32405\
        );

    \I__6693\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32405\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32402\
        );

    \I__6691\ : Span4Mux_s1_h
    port map (
            O => \N__32433\,
            I => \N__32395\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__32430\,
            I => \N__32395\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__32425\,
            I => \N__32395\
        );

    \I__6688\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32392\
        );

    \I__6687\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32389\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32385\
        );

    \I__6685\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32378\
        );

    \I__6684\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32378\
        );

    \I__6683\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32378\
        );

    \I__6682\ : InMux
    port map (
            O => \N__32414\,
            I => \N__32371\
        );

    \I__6681\ : InMux
    port map (
            O => \N__32413\,
            I => \N__32371\
        );

    \I__6680\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32371\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32364\
        );

    \I__6678\ : Span4Mux_s1_h
    port map (
            O => \N__32402\,
            I => \N__32364\
        );

    \I__6677\ : Span4Mux_h
    port map (
            O => \N__32395\,
            I => \N__32359\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__32392\,
            I => \N__32354\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__32389\,
            I => \N__32354\
        );

    \I__6674\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32351\
        );

    \I__6673\ : Span4Mux_v
    port map (
            O => \N__32385\,
            I => \N__32348\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32343\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__32371\,
            I => \N__32343\
        );

    \I__6670\ : InMux
    port map (
            O => \N__32370\,
            I => \N__32338\
        );

    \I__6669\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32338\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__32364\,
            I => \N__32335\
        );

    \I__6667\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32330\
        );

    \I__6666\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32327\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__32359\,
            I => \N__32324\
        );

    \I__6664\ : Span12Mux_s5_h
    port map (
            O => \N__32354\,
            I => \N__32313\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32313\
        );

    \I__6662\ : Sp12to4
    port map (
            O => \N__32348\,
            I => \N__32313\
        );

    \I__6661\ : Span12Mux_v
    port map (
            O => \N__32343\,
            I => \N__32313\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__32338\,
            I => \N__32313\
        );

    \I__6659\ : Span4Mux_h
    port map (
            O => \N__32335\,
            I => \N__32310\
        );

    \I__6658\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32307\
        );

    \I__6657\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32304\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__32330\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__32327\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6654\ : Odrv4
    port map (
            O => \N__32324\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6653\ : Odrv12
    port map (
            O => \N__32313\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__32310\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__32307\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__32304\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__6649\ : InMux
    port map (
            O => \N__32289\,
            I => \N__32284\
        );

    \I__6648\ : InMux
    port map (
            O => \N__32288\,
            I => \N__32281\
        );

    \I__6647\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32278\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__32284\,
            I => \N__32268\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__32281\,
            I => \N__32268\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__32278\,
            I => \N__32268\
        );

    \I__6643\ : InMux
    port map (
            O => \N__32277\,
            I => \N__32265\
        );

    \I__6642\ : CascadeMux
    port map (
            O => \N__32276\,
            I => \N__32262\
        );

    \I__6641\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32257\
        );

    \I__6640\ : Span4Mux_v
    port map (
            O => \N__32268\,
            I => \N__32254\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32251\
        );

    \I__6638\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32248\
        );

    \I__6637\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32244\
        );

    \I__6636\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32241\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__32257\,
            I => \N__32236\
        );

    \I__6634\ : IoSpan4Mux
    port map (
            O => \N__32254\,
            I => \N__32236\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__32251\,
            I => \N__32229\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__32248\,
            I => \N__32229\
        );

    \I__6631\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32226\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32218\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__32241\,
            I => \N__32218\
        );

    \I__6628\ : Span4Mux_s3_h
    port map (
            O => \N__32236\,
            I => \N__32218\
        );

    \I__6627\ : InMux
    port map (
            O => \N__32235\,
            I => \N__32215\
        );

    \I__6626\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32212\
        );

    \I__6625\ : Span4Mux_h
    port map (
            O => \N__32229\,
            I => \N__32209\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__32226\,
            I => \N__32206\
        );

    \I__6623\ : InMux
    port map (
            O => \N__32225\,
            I => \N__32203\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__32218\,
            I => \N__32198\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__32215\,
            I => \N__32198\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__32212\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__32209\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__6618\ : Odrv12
    port map (
            O => \N__32206\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__32203\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__32198\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__6615\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32184\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__32184\,
            I => \N__32181\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__6612\ : Odrv4
    port map (
            O => \N__32178\,
            I => \c0.n17710\
        );

    \I__6611\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32162\
        );

    \I__6610\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32162\
        );

    \I__6609\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32157\
        );

    \I__6608\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32157\
        );

    \I__6607\ : InMux
    port map (
            O => \N__32171\,
            I => \N__32154\
        );

    \I__6606\ : CascadeMux
    port map (
            O => \N__32170\,
            I => \N__32150\
        );

    \I__6605\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32143\
        );

    \I__6604\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32136\
        );

    \I__6603\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32136\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__32162\,
            I => \N__32133\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__32157\,
            I => \N__32128\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32128\
        );

    \I__6599\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32123\
        );

    \I__6598\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32123\
        );

    \I__6597\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32120\
        );

    \I__6596\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32113\
        );

    \I__6595\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32113\
        );

    \I__6594\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32113\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32110\
        );

    \I__6592\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32104\
        );

    \I__6591\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32104\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__32101\
        );

    \I__6589\ : Span4Mux_v
    port map (
            O => \N__32133\,
            I => \N__32096\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__32128\,
            I => \N__32096\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__32087\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32087\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32087\
        );

    \I__6584\ : Span4Mux_v
    port map (
            O => \N__32110\,
            I => \N__32087\
        );

    \I__6583\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32084\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__32104\,
            I => \N__32077\
        );

    \I__6581\ : Span4Mux_v
    port map (
            O => \N__32101\,
            I => \N__32077\
        );

    \I__6580\ : Span4Mux_h
    port map (
            O => \N__32096\,
            I => \N__32077\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__32087\,
            I => \N__32072\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__32084\,
            I => \N__32072\
        );

    \I__6577\ : Span4Mux_h
    port map (
            O => \N__32077\,
            I => \N__32066\
        );

    \I__6576\ : Span4Mux_h
    port map (
            O => \N__32072\,
            I => \N__32063\
        );

    \I__6575\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32056\
        );

    \I__6574\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32056\
        );

    \I__6573\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32056\
        );

    \I__6572\ : Odrv4
    port map (
            O => \N__32066\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__6571\ : Odrv4
    port map (
            O => \N__32063\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__32056\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__6569\ : SRMux
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__32046\,
            I => \c0.n4_adj_2154\
        );

    \I__6567\ : SRMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32037\
        );

    \I__6565\ : Span4Mux_h
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__32034\,
            I => \c0.n4_adj_2345\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__32031\,
            I => \N__32027\
        );

    \I__6562\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32024\
        );

    \I__6561\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32021\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__32024\,
            I => rand_setpoint_28
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__32021\,
            I => rand_setpoint_28
        );

    \I__6558\ : InMux
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__32013\,
            I => \N__32009\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__32012\,
            I => \N__32006\
        );

    \I__6555\ : Span12Mux_s3_v
    port map (
            O => \N__32009\,
            I => \N__32003\
        );

    \I__6554\ : InMux
    port map (
            O => \N__32006\,
            I => \N__32000\
        );

    \I__6553\ : Odrv12
    port map (
            O => \N__32003\,
            I => rand_setpoint_11
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__32000\,
            I => rand_setpoint_11
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__31995\,
            I => \N__31992\
        );

    \I__6550\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31989\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31986\
        );

    \I__6548\ : Span4Mux_s2_v
    port map (
            O => \N__31986\,
            I => \N__31983\
        );

    \I__6547\ : Span4Mux_h
    port map (
            O => \N__31983\,
            I => \N__31980\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__31980\,
            I => \c0.n17585\
        );

    \I__6545\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31974\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__31974\,
            I => \N__31970\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__31973\,
            I => \N__31967\
        );

    \I__6542\ : Span4Mux_s3_v
    port map (
            O => \N__31970\,
            I => \N__31964\
        );

    \I__6541\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31961\
        );

    \I__6540\ : Odrv4
    port map (
            O => \N__31964\,
            I => rand_setpoint_10
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__31961\,
            I => rand_setpoint_10
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__31956\,
            I => \c0.n17583_cascade_\
        );

    \I__6537\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31949\
        );

    \I__6536\ : CascadeMux
    port map (
            O => \N__31952\,
            I => \N__31946\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31943\
        );

    \I__6534\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31940\
        );

    \I__6533\ : Span4Mux_h
    port map (
            O => \N__31943\,
            I => \N__31934\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31930\
        );

    \I__6531\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31927\
        );

    \I__6530\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31922\
        );

    \I__6529\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31922\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__31934\,
            I => \N__31919\
        );

    \I__6527\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31916\
        );

    \I__6526\ : Span4Mux_h
    port map (
            O => \N__31930\,
            I => \N__31913\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__31927\,
            I => \N__31908\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__31922\,
            I => \N__31908\
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__31919\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__31916\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__31913\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6520\ : Odrv12
    port map (
            O => \N__31908\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__6519\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__31896\,
            I => \N__31892\
        );

    \I__6517\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31887\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__31892\,
            I => \N__31884\
        );

    \I__6515\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31879\
        );

    \I__6514\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31879\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31876\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__31884\,
            I => \c0.rx.n17022\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__31879\,
            I => \c0.rx.n17022\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__31876\,
            I => \c0.rx.n17022\
        );

    \I__6509\ : CascadeMux
    port map (
            O => \N__31869\,
            I => \N__31863\
        );

    \I__6508\ : InMux
    port map (
            O => \N__31868\,
            I => \N__31854\
        );

    \I__6507\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31854\
        );

    \I__6506\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31854\
        );

    \I__6505\ : InMux
    port map (
            O => \N__31863\,
            I => \N__31854\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__31854\,
            I => \N__31845\
        );

    \I__6503\ : InMux
    port map (
            O => \N__31853\,
            I => \N__31842\
        );

    \I__6502\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31839\
        );

    \I__6501\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31836\
        );

    \I__6500\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31829\
        );

    \I__6499\ : InMux
    port map (
            O => \N__31849\,
            I => \N__31829\
        );

    \I__6498\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31829\
        );

    \I__6497\ : Span4Mux_s1_v
    port map (
            O => \N__31845\,
            I => \N__31826\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__31842\,
            I => \N__31823\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__31839\,
            I => \N__31818\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31818\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31815\
        );

    \I__6492\ : Sp12to4
    port map (
            O => \N__31826\,
            I => \N__31810\
        );

    \I__6491\ : Span12Mux_s1_v
    port map (
            O => \N__31823\,
            I => \N__31810\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__31818\,
            I => \N__31805\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__31815\,
            I => \N__31805\
        );

    \I__6488\ : Odrv12
    port map (
            O => \N__31810\,
            I => \r_SM_Main_2\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__31805\,
            I => \r_SM_Main_2\
        );

    \I__6486\ : SRMux
    port map (
            O => \N__31800\,
            I => \N__31797\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__6483\ : Span4Mux_h
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__6482\ : Odrv4
    port map (
            O => \N__31788\,
            I => \c0.rx.n17058\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \N__31782\
        );

    \I__6480\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31776\
        );

    \I__6479\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31776\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__31776\,
            I => \N__31771\
        );

    \I__6477\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31768\
        );

    \I__6476\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31764\
        );

    \I__6475\ : Span4Mux_h
    port map (
            O => \N__31771\,
            I => \N__31761\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31758\
        );

    \I__6473\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31755\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__31764\,
            I => \N__31752\
        );

    \I__6471\ : Span4Mux_h
    port map (
            O => \N__31761\,
            I => \N__31749\
        );

    \I__6470\ : Span4Mux_h
    port map (
            O => \N__31758\,
            I => \N__31746\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__31755\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6468\ : Odrv12
    port map (
            O => \N__31752\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__31749\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__31746\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__6465\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31730\
        );

    \I__6464\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31730\
        );

    \I__6463\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31727\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__31730\,
            I => \N__31723\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__31727\,
            I => \N__31720\
        );

    \I__6460\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31716\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__31723\,
            I => \N__31713\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__31720\,
            I => \N__31710\
        );

    \I__6457\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31707\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__31716\,
            I => \N__31698\
        );

    \I__6455\ : Span4Mux_h
    port map (
            O => \N__31713\,
            I => \N__31698\
        );

    \I__6454\ : Span4Mux_s0_v
    port map (
            O => \N__31710\,
            I => \N__31698\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__31707\,
            I => \N__31698\
        );

    \I__6452\ : Odrv4
    port map (
            O => \N__31698\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__6450\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31686\
        );

    \I__6449\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31686\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__31686\,
            I => \N__31683\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__31680\,
            I => \c0.rx.n17080\
        );

    \I__6445\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31671\
        );

    \I__6444\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31668\
        );

    \I__6443\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31665\
        );

    \I__6442\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31662\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__31671\,
            I => \N__31659\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31656\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__31665\,
            I => \N__31652\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__31662\,
            I => \N__31649\
        );

    \I__6437\ : Span4Mux_v
    port map (
            O => \N__31659\,
            I => \N__31646\
        );

    \I__6436\ : Span4Mux_v
    port map (
            O => \N__31656\,
            I => \N__31643\
        );

    \I__6435\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31640\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__31652\,
            I => \N__31633\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__31649\,
            I => \N__31633\
        );

    \I__6432\ : Span4Mux_h
    port map (
            O => \N__31646\,
            I => \N__31633\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__31643\,
            I => rand_data_26
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__31640\,
            I => rand_data_26
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__31633\,
            I => rand_data_26
        );

    \I__6428\ : InMux
    port map (
            O => \N__31626\,
            I => n16035
        );

    \I__6427\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31619\
        );

    \I__6426\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31615\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__31619\,
            I => \N__31611\
        );

    \I__6424\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31608\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31605\
        );

    \I__6422\ : InMux
    port map (
            O => \N__31614\,
            I => \N__31602\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__31611\,
            I => \N__31597\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__31608\,
            I => \N__31597\
        );

    \I__6419\ : Span4Mux_v
    port map (
            O => \N__31605\,
            I => \N__31593\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__31602\,
            I => \N__31590\
        );

    \I__6417\ : Span4Mux_h
    port map (
            O => \N__31597\,
            I => \N__31587\
        );

    \I__6416\ : InMux
    port map (
            O => \N__31596\,
            I => \N__31584\
        );

    \I__6415\ : Span4Mux_v
    port map (
            O => \N__31593\,
            I => \N__31581\
        );

    \I__6414\ : Span12Mux_s6_v
    port map (
            O => \N__31590\,
            I => \N__31578\
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__31587\,
            I => rand_data_27
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__31584\,
            I => rand_data_27
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__31581\,
            I => rand_data_27
        );

    \I__6410\ : Odrv12
    port map (
            O => \N__31578\,
            I => rand_data_27
        );

    \I__6409\ : InMux
    port map (
            O => \N__31569\,
            I => n16036
        );

    \I__6408\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31560\
        );

    \I__6407\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31557\
        );

    \I__6406\ : InMux
    port map (
            O => \N__31564\,
            I => \N__31554\
        );

    \I__6405\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31551\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31548\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__31557\,
            I => \N__31545\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31539\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31539\
        );

    \I__6400\ : Span4Mux_h
    port map (
            O => \N__31548\,
            I => \N__31536\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__31545\,
            I => \N__31533\
        );

    \I__6398\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31530\
        );

    \I__6397\ : Span4Mux_v
    port map (
            O => \N__31539\,
            I => \N__31525\
        );

    \I__6396\ : Span4Mux_h
    port map (
            O => \N__31536\,
            I => \N__31525\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__31533\,
            I => rand_data_28
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__31530\,
            I => rand_data_28
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__31525\,
            I => rand_data_28
        );

    \I__6392\ : InMux
    port map (
            O => \N__31518\,
            I => n16037
        );

    \I__6391\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31510\
        );

    \I__6390\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31507\
        );

    \I__6389\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31503\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31500\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__31507\,
            I => \N__31497\
        );

    \I__6386\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31494\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__31503\,
            I => \N__31491\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__31500\,
            I => \N__31488\
        );

    \I__6383\ : Span4Mux_v
    port map (
            O => \N__31497\,
            I => \N__31483\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__31494\,
            I => \N__31483\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__31491\,
            I => \N__31479\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__31488\,
            I => \N__31474\
        );

    \I__6379\ : Span4Mux_h
    port map (
            O => \N__31483\,
            I => \N__31474\
        );

    \I__6378\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31471\
        );

    \I__6377\ : Span4Mux_h
    port map (
            O => \N__31479\,
            I => \N__31468\
        );

    \I__6376\ : Odrv4
    port map (
            O => \N__31474\,
            I => rand_data_29
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__31471\,
            I => rand_data_29
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__31468\,
            I => rand_data_29
        );

    \I__6373\ : InMux
    port map (
            O => \N__31461\,
            I => n16038
        );

    \I__6372\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31455\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__31455\,
            I => \N__31450\
        );

    \I__6370\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31446\
        );

    \I__6369\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31443\
        );

    \I__6368\ : Span4Mux_s1_h
    port map (
            O => \N__31450\,
            I => \N__31440\
        );

    \I__6367\ : InMux
    port map (
            O => \N__31449\,
            I => \N__31437\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__31446\,
            I => \N__31434\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__31443\,
            I => \N__31431\
        );

    \I__6364\ : Span4Mux_v
    port map (
            O => \N__31440\,
            I => \N__31425\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31425\
        );

    \I__6362\ : Span4Mux_v
    port map (
            O => \N__31434\,
            I => \N__31422\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__31431\,
            I => \N__31419\
        );

    \I__6360\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31416\
        );

    \I__6359\ : Span4Mux_h
    port map (
            O => \N__31425\,
            I => \N__31411\
        );

    \I__6358\ : Span4Mux_h
    port map (
            O => \N__31422\,
            I => \N__31411\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__31419\,
            I => rand_data_30
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__31416\,
            I => rand_data_30
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__31411\,
            I => rand_data_30
        );

    \I__6354\ : InMux
    port map (
            O => \N__31404\,
            I => n16039
        );

    \I__6353\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31396\
        );

    \I__6352\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31393\
        );

    \I__6351\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31389\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__31396\,
            I => \N__31386\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__31393\,
            I => \N__31383\
        );

    \I__6348\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31380\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__31389\,
            I => \N__31377\
        );

    \I__6346\ : Span4Mux_h
    port map (
            O => \N__31386\,
            I => \N__31373\
        );

    \I__6345\ : Span4Mux_v
    port map (
            O => \N__31383\,
            I => \N__31368\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31368\
        );

    \I__6343\ : Span4Mux_v
    port map (
            O => \N__31377\,
            I => \N__31365\
        );

    \I__6342\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31362\
        );

    \I__6341\ : Span4Mux_h
    port map (
            O => \N__31373\,
            I => \N__31357\
        );

    \I__6340\ : Span4Mux_h
    port map (
            O => \N__31368\,
            I => \N__31357\
        );

    \I__6339\ : Sp12to4
    port map (
            O => \N__31365\,
            I => \N__31354\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__31362\,
            I => rand_data_31
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__31357\,
            I => rand_data_31
        );

    \I__6336\ : Odrv12
    port map (
            O => \N__31354\,
            I => rand_data_31
        );

    \I__6335\ : InMux
    port map (
            O => \N__31347\,
            I => n16040
        );

    \I__6334\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31341\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__6332\ : Span4Mux_s2_v
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__6331\ : Span4Mux_h
    port map (
            O => \N__31335\,
            I => \N__31331\
        );

    \I__6330\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31328\
        );

    \I__6329\ : Span4Mux_h
    port map (
            O => \N__31331\,
            I => \N__31325\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__31328\,
            I => rand_setpoint_31
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__31325\,
            I => rand_setpoint_31
        );

    \I__6326\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31316\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__31319\,
            I => \N__31313\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__31316\,
            I => \N__31310\
        );

    \I__6323\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31307\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__31310\,
            I => rand_setpoint_26
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__31307\,
            I => rand_setpoint_26
        );

    \I__6320\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31298\
        );

    \I__6319\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31295\
        );

    \I__6318\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31292\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__31295\,
            I => rand_setpoint_29
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__31292\,
            I => rand_setpoint_29
        );

    \I__6315\ : CascadeMux
    port map (
            O => \N__31287\,
            I => \N__31283\
        );

    \I__6314\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31280\
        );

    \I__6313\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31277\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__31280\,
            I => rand_setpoint_27
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__31277\,
            I => rand_setpoint_27
        );

    \I__6310\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31265\
        );

    \I__6308\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31260\
        );

    \I__6307\ : Span4Mux_v
    port map (
            O => \N__31265\,
            I => \N__31257\
        );

    \I__6306\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31254\
        );

    \I__6305\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31251\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__31260\,
            I => \N__31248\
        );

    \I__6303\ : Span4Mux_v
    port map (
            O => \N__31257\,
            I => \N__31245\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31242\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31239\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__31248\,
            I => \N__31235\
        );

    \I__6299\ : Span4Mux_s3_h
    port map (
            O => \N__31245\,
            I => \N__31232\
        );

    \I__6298\ : Span4Mux_v
    port map (
            O => \N__31242\,
            I => \N__31227\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__31239\,
            I => \N__31227\
        );

    \I__6296\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31224\
        );

    \I__6295\ : Span4Mux_h
    port map (
            O => \N__31235\,
            I => \N__31221\
        );

    \I__6294\ : Odrv4
    port map (
            O => \N__31232\,
            I => rand_data_18
        );

    \I__6293\ : Odrv4
    port map (
            O => \N__31227\,
            I => rand_data_18
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__31224\,
            I => rand_data_18
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__31221\,
            I => rand_data_18
        );

    \I__6290\ : InMux
    port map (
            O => \N__31212\,
            I => n16027
        );

    \I__6289\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31205\
        );

    \I__6288\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31202\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__31205\,
            I => \N__31198\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__31202\,
            I => \N__31195\
        );

    \I__6285\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31191\
        );

    \I__6284\ : Span4Mux_h
    port map (
            O => \N__31198\,
            I => \N__31188\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__31195\,
            I => \N__31185\
        );

    \I__6282\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31182\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31178\
        );

    \I__6280\ : Sp12to4
    port map (
            O => \N__31188\,
            I => \N__31171\
        );

    \I__6279\ : Sp12to4
    port map (
            O => \N__31185\,
            I => \N__31171\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31171\
        );

    \I__6277\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31168\
        );

    \I__6276\ : Span12Mux_s7_v
    port map (
            O => \N__31178\,
            I => \N__31165\
        );

    \I__6275\ : Odrv12
    port map (
            O => \N__31171\,
            I => rand_data_19
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__31168\,
            I => rand_data_19
        );

    \I__6273\ : Odrv12
    port map (
            O => \N__31165\,
            I => rand_data_19
        );

    \I__6272\ : InMux
    port map (
            O => \N__31158\,
            I => n16028
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__31155\,
            I => \N__31151\
        );

    \I__6270\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31146\
        );

    \I__6269\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31143\
        );

    \I__6268\ : InMux
    port map (
            O => \N__31150\,
            I => \N__31140\
        );

    \I__6267\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31137\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__31146\,
            I => \N__31134\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__31143\,
            I => \N__31131\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__31140\,
            I => \N__31128\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31124\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__31134\,
            I => \N__31121\
        );

    \I__6261\ : Span4Mux_h
    port map (
            O => \N__31131\,
            I => \N__31118\
        );

    \I__6260\ : Span4Mux_v
    port map (
            O => \N__31128\,
            I => \N__31115\
        );

    \I__6259\ : InMux
    port map (
            O => \N__31127\,
            I => \N__31112\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__31124\,
            I => \N__31107\
        );

    \I__6257\ : Span4Mux_h
    port map (
            O => \N__31121\,
            I => \N__31107\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__31118\,
            I => rand_data_20
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__31115\,
            I => rand_data_20
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__31112\,
            I => rand_data_20
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__31107\,
            I => rand_data_20
        );

    \I__6252\ : InMux
    port map (
            O => \N__31098\,
            I => n16029
        );

    \I__6251\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31091\
        );

    \I__6250\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31086\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__31091\,
            I => \N__31083\
        );

    \I__6248\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31080\
        );

    \I__6247\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31077\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__31086\,
            I => \N__31074\
        );

    \I__6245\ : Span4Mux_h
    port map (
            O => \N__31083\,
            I => \N__31071\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__31080\,
            I => \N__31068\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__31077\,
            I => \N__31065\
        );

    \I__6242\ : Span4Mux_h
    port map (
            O => \N__31074\,
            I => \N__31061\
        );

    \I__6241\ : Span4Mux_v
    port map (
            O => \N__31071\,
            I => \N__31058\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__31068\,
            I => \N__31055\
        );

    \I__6239\ : Span4Mux_h
    port map (
            O => \N__31065\,
            I => \N__31052\
        );

    \I__6238\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31049\
        );

    \I__6237\ : Span4Mux_h
    port map (
            O => \N__31061\,
            I => \N__31046\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__31058\,
            I => rand_data_21
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__31055\,
            I => rand_data_21
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__31052\,
            I => rand_data_21
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__31049\,
            I => rand_data_21
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__31046\,
            I => rand_data_21
        );

    \I__6231\ : InMux
    port map (
            O => \N__31035\,
            I => n16030
        );

    \I__6230\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31027\
        );

    \I__6229\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31023\
        );

    \I__6228\ : InMux
    port map (
            O => \N__31030\,
            I => \N__31020\
        );

    \I__6227\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31017\
        );

    \I__6226\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31014\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__31023\,
            I => \N__31011\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__31020\,
            I => \N__31008\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__31003\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__31014\,
            I => \N__31003\
        );

    \I__6221\ : Span4Mux_h
    port map (
            O => \N__31011\,
            I => \N__30999\
        );

    \I__6220\ : Span4Mux_v
    port map (
            O => \N__31008\,
            I => \N__30996\
        );

    \I__6219\ : Span4Mux_v
    port map (
            O => \N__31003\,
            I => \N__30993\
        );

    \I__6218\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30990\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__30999\,
            I => \N__30987\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__30996\,
            I => rand_data_22
        );

    \I__6215\ : Odrv4
    port map (
            O => \N__30993\,
            I => rand_data_22
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__30990\,
            I => rand_data_22
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__30987\,
            I => rand_data_22
        );

    \I__6212\ : InMux
    port map (
            O => \N__30978\,
            I => n16031
        );

    \I__6211\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30971\
        );

    \I__6210\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30967\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__30971\,
            I => \N__30964\
        );

    \I__6208\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30961\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__30967\,
            I => \N__30957\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__30964\,
            I => \N__30952\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30952\
        );

    \I__6204\ : InMux
    port map (
            O => \N__30960\,
            I => \N__30949\
        );

    \I__6203\ : Span4Mux_h
    port map (
            O => \N__30957\,
            I => \N__30945\
        );

    \I__6202\ : Span4Mux_v
    port map (
            O => \N__30952\,
            I => \N__30942\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__30949\,
            I => \N__30939\
        );

    \I__6200\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30936\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__30945\,
            I => \N__30933\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__30942\,
            I => rand_data_23
        );

    \I__6197\ : Odrv12
    port map (
            O => \N__30939\,
            I => rand_data_23
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__30936\,
            I => rand_data_23
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__30933\,
            I => rand_data_23
        );

    \I__6194\ : InMux
    port map (
            O => \N__30924\,
            I => n16032
        );

    \I__6193\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30916\
        );

    \I__6192\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30912\
        );

    \I__6191\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30909\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30906\
        );

    \I__6189\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30903\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30900\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__30909\,
            I => \N__30896\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__30906\,
            I => \N__30891\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__30903\,
            I => \N__30891\
        );

    \I__6184\ : Span4Mux_h
    port map (
            O => \N__30900\,
            I => \N__30888\
        );

    \I__6183\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30885\
        );

    \I__6182\ : Span4Mux_v
    port map (
            O => \N__30896\,
            I => \N__30878\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__30891\,
            I => \N__30878\
        );

    \I__6180\ : Span4Mux_h
    port map (
            O => \N__30888\,
            I => \N__30878\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__30885\,
            I => rand_data_24
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__30878\,
            I => rand_data_24
        );

    \I__6177\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30867\
        );

    \I__6175\ : Span4Mux_s2_v
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__30864\,
            I => \N__30860\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__30863\,
            I => \N__30857\
        );

    \I__6172\ : Span4Mux_h
    port map (
            O => \N__30860\,
            I => \N__30854\
        );

    \I__6171\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30851\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__30854\,
            I => rand_setpoint_24
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__30851\,
            I => rand_setpoint_24
        );

    \I__6168\ : InMux
    port map (
            O => \N__30846\,
            I => \bfn_10_28_0_\
        );

    \I__6167\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30839\
        );

    \I__6166\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30835\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__30839\,
            I => \N__30831\
        );

    \I__6164\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30828\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30825\
        );

    \I__6162\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30822\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__30831\,
            I => \N__30819\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30816\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__30825\,
            I => \N__30811\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__30822\,
            I => \N__30811\
        );

    \I__6157\ : Span4Mux_s0_h
    port map (
            O => \N__30819\,
            I => \N__30807\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__30816\,
            I => \N__30804\
        );

    \I__6155\ : Span4Mux_v
    port map (
            O => \N__30811\,
            I => \N__30801\
        );

    \I__6154\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30798\
        );

    \I__6153\ : Span4Mux_h
    port map (
            O => \N__30807\,
            I => \N__30793\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__30804\,
            I => \N__30793\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__30801\,
            I => rand_data_25
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__30798\,
            I => rand_data_25
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__30793\,
            I => rand_data_25
        );

    \I__6148\ : InMux
    port map (
            O => \N__30786\,
            I => n16034
        );

    \I__6147\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30776\
        );

    \I__6146\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30773\
        );

    \I__6145\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30770\
        );

    \I__6144\ : InMux
    port map (
            O => \N__30780\,
            I => \N__30767\
        );

    \I__6143\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30764\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__30776\,
            I => \N__30761\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__30773\,
            I => \N__30758\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__30770\,
            I => \N__30755\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__30767\,
            I => \N__30752\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__30764\,
            I => \N__30748\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__30761\,
            I => \N__30743\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__30758\,
            I => \N__30743\
        );

    \I__6135\ : Span12Mux_h
    port map (
            O => \N__30755\,
            I => \N__30740\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__30752\,
            I => \N__30737\
        );

    \I__6133\ : InMux
    port map (
            O => \N__30751\,
            I => \N__30734\
        );

    \I__6132\ : Span12Mux_h
    port map (
            O => \N__30748\,
            I => \N__30731\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__30743\,
            I => rand_data_10
        );

    \I__6130\ : Odrv12
    port map (
            O => \N__30740\,
            I => rand_data_10
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__30737\,
            I => rand_data_10
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__30734\,
            I => rand_data_10
        );

    \I__6127\ : Odrv12
    port map (
            O => \N__30731\,
            I => rand_data_10
        );

    \I__6126\ : InMux
    port map (
            O => \N__30720\,
            I => n16019
        );

    \I__6125\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30713\
        );

    \I__6124\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30710\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__30713\,
            I => \N__30704\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__30710\,
            I => \N__30701\
        );

    \I__6121\ : InMux
    port map (
            O => \N__30709\,
            I => \N__30698\
        );

    \I__6120\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30695\
        );

    \I__6119\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30692\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__30704\,
            I => \N__30689\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__30701\,
            I => \N__30682\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__30698\,
            I => \N__30682\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30682\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__30692\,
            I => \N__30678\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__30689\,
            I => \N__30673\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__30682\,
            I => \N__30673\
        );

    \I__6111\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30670\
        );

    \I__6110\ : Span12Mux_s8_v
    port map (
            O => \N__30678\,
            I => \N__30667\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__30673\,
            I => rand_data_11
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__30670\,
            I => rand_data_11
        );

    \I__6107\ : Odrv12
    port map (
            O => \N__30667\,
            I => rand_data_11
        );

    \I__6106\ : InMux
    port map (
            O => \N__30660\,
            I => n16020
        );

    \I__6105\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30650\
        );

    \I__6104\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30650\
        );

    \I__6103\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30647\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__30650\,
            I => \N__30642\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__30647\,
            I => \N__30639\
        );

    \I__6100\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30636\
        );

    \I__6099\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30633\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__30642\,
            I => \N__30630\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__30639\,
            I => \N__30626\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30621\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30621\
        );

    \I__6094\ : Sp12to4
    port map (
            O => \N__30630\,
            I => \N__30618\
        );

    \I__6093\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30615\
        );

    \I__6092\ : Span4Mux_h
    port map (
            O => \N__30626\,
            I => \N__30612\
        );

    \I__6091\ : Odrv12
    port map (
            O => \N__30621\,
            I => rand_data_12
        );

    \I__6090\ : Odrv12
    port map (
            O => \N__30618\,
            I => rand_data_12
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__30615\,
            I => rand_data_12
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__30612\,
            I => rand_data_12
        );

    \I__6087\ : InMux
    port map (
            O => \N__30603\,
            I => n16021
        );

    \I__6086\ : InMux
    port map (
            O => \N__30600\,
            I => \N__30595\
        );

    \I__6085\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30591\
        );

    \I__6084\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30588\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__30595\,
            I => \N__30585\
        );

    \I__6082\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30581\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__30591\,
            I => \N__30578\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__30588\,
            I => \N__30575\
        );

    \I__6079\ : Span4Mux_h
    port map (
            O => \N__30585\,
            I => \N__30571\
        );

    \I__6078\ : InMux
    port map (
            O => \N__30584\,
            I => \N__30568\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__30581\,
            I => \N__30565\
        );

    \I__6076\ : Span4Mux_h
    port map (
            O => \N__30578\,
            I => \N__30562\
        );

    \I__6075\ : Span4Mux_v
    port map (
            O => \N__30575\,
            I => \N__30559\
        );

    \I__6074\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30556\
        );

    \I__6073\ : Span4Mux_h
    port map (
            O => \N__30571\,
            I => \N__30553\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__30568\,
            I => rand_data_13
        );

    \I__6071\ : Odrv12
    port map (
            O => \N__30565\,
            I => rand_data_13
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__30562\,
            I => rand_data_13
        );

    \I__6069\ : Odrv4
    port map (
            O => \N__30559\,
            I => rand_data_13
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__30556\,
            I => rand_data_13
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__30553\,
            I => rand_data_13
        );

    \I__6066\ : InMux
    port map (
            O => \N__30540\,
            I => n16022
        );

    \I__6065\ : CascadeMux
    port map (
            O => \N__30537\,
            I => \N__30530\
        );

    \I__6064\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30527\
        );

    \I__6063\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30524\
        );

    \I__6062\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30521\
        );

    \I__6061\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30518\
        );

    \I__6060\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30515\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__30527\,
            I => \N__30512\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30509\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30506\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__30518\,
            I => \N__30503\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__30515\,
            I => \N__30497\
        );

    \I__6054\ : Span4Mux_h
    port map (
            O => \N__30512\,
            I => \N__30497\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__30509\,
            I => \N__30494\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__30506\,
            I => \N__30491\
        );

    \I__6051\ : Sp12to4
    port map (
            O => \N__30503\,
            I => \N__30488\
        );

    \I__6050\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30485\
        );

    \I__6049\ : Span4Mux_v
    port map (
            O => \N__30497\,
            I => \N__30480\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__30494\,
            I => \N__30480\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__30491\,
            I => rand_data_14
        );

    \I__6046\ : Odrv12
    port map (
            O => \N__30488\,
            I => rand_data_14
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__30485\,
            I => rand_data_14
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__30480\,
            I => rand_data_14
        );

    \I__6043\ : InMux
    port map (
            O => \N__30471\,
            I => n16023
        );

    \I__6042\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30462\
        );

    \I__6041\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30459\
        );

    \I__6040\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30454\
        );

    \I__6039\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30454\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30451\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30448\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__30454\,
            I => \N__30443\
        );

    \I__6035\ : Span4Mux_v
    port map (
            O => \N__30451\,
            I => \N__30440\
        );

    \I__6034\ : Span4Mux_v
    port map (
            O => \N__30448\,
            I => \N__30437\
        );

    \I__6033\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30434\
        );

    \I__6032\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30431\
        );

    \I__6031\ : Span4Mux_s2_h
    port map (
            O => \N__30443\,
            I => \N__30426\
        );

    \I__6030\ : Span4Mux_h
    port map (
            O => \N__30440\,
            I => \N__30426\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__30437\,
            I => rand_data_15
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__30434\,
            I => rand_data_15
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__30431\,
            I => rand_data_15
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__30426\,
            I => rand_data_15
        );

    \I__6025\ : InMux
    port map (
            O => \N__30417\,
            I => n16024
        );

    \I__6024\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30410\
        );

    \I__6023\ : InMux
    port map (
            O => \N__30413\,
            I => \N__30407\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__30410\,
            I => \N__30402\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30399\
        );

    \I__6020\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30396\
        );

    \I__6019\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30393\
        );

    \I__6018\ : Span4Mux_h
    port map (
            O => \N__30402\,
            I => \N__30389\
        );

    \I__6017\ : Span12Mux_s4_h
    port map (
            O => \N__30399\,
            I => \N__30384\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__30396\,
            I => \N__30384\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__30393\,
            I => \N__30381\
        );

    \I__6014\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30378\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__30389\,
            I => \N__30375\
        );

    \I__6012\ : Odrv12
    port map (
            O => \N__30384\,
            I => rand_data_16
        );

    \I__6011\ : Odrv12
    port map (
            O => \N__30381\,
            I => rand_data_16
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__30378\,
            I => rand_data_16
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__30375\,
            I => rand_data_16
        );

    \I__6008\ : InMux
    port map (
            O => \N__30366\,
            I => \bfn_10_27_0_\
        );

    \I__6007\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__30360\,
            I => \N__30356\
        );

    \I__6005\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30352\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__30356\,
            I => \N__30348\
        );

    \I__6003\ : InMux
    port map (
            O => \N__30355\,
            I => \N__30345\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__30352\,
            I => \N__30342\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__30351\,
            I => \N__30339\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__30348\,
            I => \N__30336\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__30345\,
            I => \N__30333\
        );

    \I__5998\ : Span4Mux_h
    port map (
            O => \N__30342\,
            I => \N__30330\
        );

    \I__5997\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30326\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__30336\,
            I => \N__30321\
        );

    \I__5995\ : Span4Mux_h
    port map (
            O => \N__30333\,
            I => \N__30321\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__30330\,
            I => \N__30318\
        );

    \I__5993\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30315\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30310\
        );

    \I__5991\ : Span4Mux_h
    port map (
            O => \N__30321\,
            I => \N__30310\
        );

    \I__5990\ : Odrv4
    port map (
            O => \N__30318\,
            I => rand_data_17
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__30315\,
            I => rand_data_17
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__30310\,
            I => rand_data_17
        );

    \I__5987\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30300\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__30300\,
            I => \N__30296\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__30299\,
            I => \N__30293\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__30296\,
            I => \N__30290\
        );

    \I__5983\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30287\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__30290\,
            I => rand_setpoint_17
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__30287\,
            I => rand_setpoint_17
        );

    \I__5980\ : InMux
    port map (
            O => \N__30282\,
            I => n16026
        );

    \I__5979\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30275\
        );

    \I__5978\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30271\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30268\
        );

    \I__5976\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30265\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__30271\,
            I => \N__30261\
        );

    \I__5974\ : Span4Mux_v
    port map (
            O => \N__30268\,
            I => \N__30258\
        );

    \I__5973\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30254\
        );

    \I__5972\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30251\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__30261\,
            I => \N__30247\
        );

    \I__5970\ : Span4Mux_h
    port map (
            O => \N__30258\,
            I => \N__30244\
        );

    \I__5969\ : InMux
    port map (
            O => \N__30257\,
            I => \N__30241\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__30254\,
            I => \N__30236\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__30251\,
            I => \N__30236\
        );

    \I__5966\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30233\
        );

    \I__5965\ : Span4Mux_s2_h
    port map (
            O => \N__30247\,
            I => \N__30228\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__30244\,
            I => \N__30228\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__30241\,
            I => rand_data_1
        );

    \I__5962\ : Odrv12
    port map (
            O => \N__30236\,
            I => rand_data_1
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__30233\,
            I => rand_data_1
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__30228\,
            I => rand_data_1
        );

    \I__5959\ : InMux
    port map (
            O => \N__30219\,
            I => n16010
        );

    \I__5958\ : InMux
    port map (
            O => \N__30216\,
            I => \N__30212\
        );

    \I__5957\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30206\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__30212\,
            I => \N__30202\
        );

    \I__5955\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30197\
        );

    \I__5954\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30197\
        );

    \I__5953\ : InMux
    port map (
            O => \N__30209\,
            I => \N__30194\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__30206\,
            I => \N__30191\
        );

    \I__5951\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30188\
        );

    \I__5950\ : Span12Mux_h
    port map (
            O => \N__30202\,
            I => \N__30185\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__30197\,
            I => rand_data_2
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__30194\,
            I => rand_data_2
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__30191\,
            I => rand_data_2
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__30188\,
            I => rand_data_2
        );

    \I__5945\ : Odrv12
    port map (
            O => \N__30185\,
            I => rand_data_2
        );

    \I__5944\ : InMux
    port map (
            O => \N__30174\,
            I => n16011
        );

    \I__5943\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30166\
        );

    \I__5942\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30163\
        );

    \I__5941\ : InMux
    port map (
            O => \N__30169\,
            I => \N__30159\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__30166\,
            I => \N__30153\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__30163\,
            I => \N__30153\
        );

    \I__5938\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30150\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__30159\,
            I => \N__30147\
        );

    \I__5936\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30144\
        );

    \I__5935\ : Span4Mux_v
    port map (
            O => \N__30153\,
            I => \N__30140\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30137\
        );

    \I__5933\ : Span4Mux_h
    port map (
            O => \N__30147\,
            I => \N__30134\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__30144\,
            I => \N__30131\
        );

    \I__5931\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30128\
        );

    \I__5930\ : Sp12to4
    port map (
            O => \N__30140\,
            I => \N__30123\
        );

    \I__5929\ : Span12Mux_s9_v
    port map (
            O => \N__30137\,
            I => \N__30123\
        );

    \I__5928\ : Odrv4
    port map (
            O => \N__30134\,
            I => rand_data_3
        );

    \I__5927\ : Odrv12
    port map (
            O => \N__30131\,
            I => rand_data_3
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__30128\,
            I => rand_data_3
        );

    \I__5925\ : Odrv12
    port map (
            O => \N__30123\,
            I => rand_data_3
        );

    \I__5924\ : InMux
    port map (
            O => \N__30114\,
            I => n16012
        );

    \I__5923\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30106\
        );

    \I__5922\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30101\
        );

    \I__5921\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30098\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__30106\,
            I => \N__30095\
        );

    \I__5919\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30092\
        );

    \I__5918\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30089\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__30101\,
            I => \N__30083\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30083\
        );

    \I__5915\ : Span4Mux_h
    port map (
            O => \N__30095\,
            I => \N__30080\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__30092\,
            I => \N__30077\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__30089\,
            I => \N__30074\
        );

    \I__5912\ : InMux
    port map (
            O => \N__30088\,
            I => \N__30071\
        );

    \I__5911\ : Span4Mux_h
    port map (
            O => \N__30083\,
            I => \N__30066\
        );

    \I__5910\ : Span4Mux_h
    port map (
            O => \N__30080\,
            I => \N__30066\
        );

    \I__5909\ : Odrv12
    port map (
            O => \N__30077\,
            I => rand_data_4
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__30074\,
            I => rand_data_4
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__30071\,
            I => rand_data_4
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__30066\,
            I => rand_data_4
        );

    \I__5905\ : InMux
    port map (
            O => \N__30057\,
            I => n16013
        );

    \I__5904\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30050\
        );

    \I__5903\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30046\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__30043\
        );

    \I__5901\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30040\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__30046\,
            I => \N__30036\
        );

    \I__5899\ : Span4Mux_h
    port map (
            O => \N__30043\,
            I => \N__30033\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__30040\,
            I => \N__30028\
        );

    \I__5897\ : InMux
    port map (
            O => \N__30039\,
            I => \N__30025\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__30036\,
            I => \N__30022\
        );

    \I__5895\ : Span4Mux_h
    port map (
            O => \N__30033\,
            I => \N__30019\
        );

    \I__5894\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30016\
        );

    \I__5893\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30013\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__30028\,
            I => \N__30006\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__30025\,
            I => \N__30006\
        );

    \I__5890\ : Span4Mux_h
    port map (
            O => \N__30022\,
            I => \N__30006\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__30019\,
            I => rand_data_5
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__30016\,
            I => rand_data_5
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__30013\,
            I => rand_data_5
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__30006\,
            I => rand_data_5
        );

    \I__5885\ : InMux
    port map (
            O => \N__29997\,
            I => n16014
        );

    \I__5884\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29988\
        );

    \I__5883\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29985\
        );

    \I__5882\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29982\
        );

    \I__5881\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29979\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__29988\,
            I => \N__29976\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29973\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__29982\,
            I => \N__29970\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29967\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__29976\,
            I => \N__29962\
        );

    \I__5875\ : Span4Mux_h
    port map (
            O => \N__29973\,
            I => \N__29959\
        );

    \I__5874\ : Span4Mux_v
    port map (
            O => \N__29970\,
            I => \N__29954\
        );

    \I__5873\ : Span4Mux_h
    port map (
            O => \N__29967\,
            I => \N__29954\
        );

    \I__5872\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29951\
        );

    \I__5871\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29948\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__29962\,
            I => \N__29945\
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__29959\,
            I => rand_data_6
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__29954\,
            I => rand_data_6
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__29951\,
            I => rand_data_6
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__29948\,
            I => rand_data_6
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__29945\,
            I => rand_data_6
        );

    \I__5864\ : InMux
    port map (
            O => \N__29934\,
            I => n16015
        );

    \I__5863\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29926\
        );

    \I__5862\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29923\
        );

    \I__5861\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29920\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__29926\,
            I => \N__29917\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__29923\,
            I => \N__29913\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__29920\,
            I => \N__29907\
        );

    \I__5857\ : Span4Mux_v
    port map (
            O => \N__29917\,
            I => \N__29907\
        );

    \I__5856\ : InMux
    port map (
            O => \N__29916\,
            I => \N__29904\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__29913\,
            I => \N__29900\
        );

    \I__5854\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29897\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__29907\,
            I => \N__29892\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__29904\,
            I => \N__29892\
        );

    \I__5851\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29889\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__29900\,
            I => \N__29886\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__29897\,
            I => rand_data_7
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__29892\,
            I => rand_data_7
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__29889\,
            I => rand_data_7
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__29886\,
            I => rand_data_7
        );

    \I__5845\ : InMux
    port map (
            O => \N__29877\,
            I => n16016
        );

    \I__5844\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29869\
        );

    \I__5843\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29866\
        );

    \I__5842\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29863\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29858\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29855\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29852\
        );

    \I__5838\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29847\
        );

    \I__5837\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29847\
        );

    \I__5836\ : Span4Mux_h
    port map (
            O => \N__29858\,
            I => \N__29843\
        );

    \I__5835\ : Span4Mux_h
    port map (
            O => \N__29855\,
            I => \N__29840\
        );

    \I__5834\ : Span4Mux_h
    port map (
            O => \N__29852\,
            I => \N__29835\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__29847\,
            I => \N__29835\
        );

    \I__5832\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29832\
        );

    \I__5831\ : Span4Mux_h
    port map (
            O => \N__29843\,
            I => \N__29827\
        );

    \I__5830\ : Span4Mux_h
    port map (
            O => \N__29840\,
            I => \N__29827\
        );

    \I__5829\ : Odrv4
    port map (
            O => \N__29835\,
            I => rand_data_8
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__29832\,
            I => rand_data_8
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__29827\,
            I => rand_data_8
        );

    \I__5826\ : InMux
    port map (
            O => \N__29820\,
            I => \bfn_10_26_0_\
        );

    \I__5825\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29813\
        );

    \I__5824\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29807\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__29813\,
            I => \N__29804\
        );

    \I__5822\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29799\
        );

    \I__5821\ : InMux
    port map (
            O => \N__29811\,
            I => \N__29799\
        );

    \I__5820\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29796\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__29807\,
            I => \N__29793\
        );

    \I__5818\ : Span4Mux_v
    port map (
            O => \N__29804\,
            I => \N__29790\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__29799\,
            I => \N__29787\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29784\
        );

    \I__5815\ : Span4Mux_v
    port map (
            O => \N__29793\,
            I => \N__29780\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__29790\,
            I => \N__29775\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29775\
        );

    \I__5812\ : Sp12to4
    port map (
            O => \N__29784\,
            I => \N__29772\
        );

    \I__5811\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29769\
        );

    \I__5810\ : Span4Mux_h
    port map (
            O => \N__29780\,
            I => \N__29766\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__29775\,
            I => rand_data_9
        );

    \I__5808\ : Odrv12
    port map (
            O => \N__29772\,
            I => rand_data_9
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__29769\,
            I => rand_data_9
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__29766\,
            I => rand_data_9
        );

    \I__5805\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29754\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__29754\,
            I => \N__29750\
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__29753\,
            I => \N__29747\
        );

    \I__5802\ : Span4Mux_v
    port map (
            O => \N__29750\,
            I => \N__29744\
        );

    \I__5801\ : InMux
    port map (
            O => \N__29747\,
            I => \N__29741\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__29744\,
            I => rand_setpoint_9
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__29741\,
            I => rand_setpoint_9
        );

    \I__5798\ : InMux
    port map (
            O => \N__29736\,
            I => n16018
        );

    \I__5797\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29727\
        );

    \I__5796\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29724\
        );

    \I__5795\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29719\
        );

    \I__5794\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29719\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__29727\,
            I => data_in_3_4
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__29724\,
            I => data_in_3_4
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__29719\,
            I => data_in_3_4
        );

    \I__5790\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29707\
        );

    \I__5789\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29704\
        );

    \I__5788\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29701\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29698\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29695\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29692\
        );

    \I__5784\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29689\
        );

    \I__5783\ : Span4Mux_v
    port map (
            O => \N__29695\,
            I => \N__29686\
        );

    \I__5782\ : Span4Mux_h
    port map (
            O => \N__29692\,
            I => \N__29683\
        );

    \I__5781\ : Span4Mux_v
    port map (
            O => \N__29689\,
            I => \N__29680\
        );

    \I__5780\ : Span4Mux_v
    port map (
            O => \N__29686\,
            I => \N__29676\
        );

    \I__5779\ : Span4Mux_v
    port map (
            O => \N__29683\,
            I => \N__29673\
        );

    \I__5778\ : Span4Mux_v
    port map (
            O => \N__29680\,
            I => \N__29670\
        );

    \I__5777\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29667\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__29676\,
            I => \N__29662\
        );

    \I__5775\ : Span4Mux_v
    port map (
            O => \N__29673\,
            I => \N__29662\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__29670\,
            I => data_in_1_6
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__29667\,
            I => data_in_1_6
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__29662\,
            I => data_in_1_6
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__29655\,
            I => \N__29652\
        );

    \I__5770\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29648\
        );

    \I__5769\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29643\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__29648\,
            I => \N__29640\
        );

    \I__5767\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29637\
        );

    \I__5766\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29634\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__29643\,
            I => \N__29627\
        );

    \I__5764\ : Span4Mux_v
    port map (
            O => \N__29640\,
            I => \N__29627\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29627\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__29634\,
            I => data_in_3_5
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__29627\,
            I => data_in_3_5
        );

    \I__5760\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29619\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__29619\,
            I => \c0.n17402\
        );

    \I__5758\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29613\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__29610\,
            I => \N__29605\
        );

    \I__5755\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29602\
        );

    \I__5754\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29599\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__29605\,
            I => \N__29596\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__29602\,
            I => \N__29593\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__29599\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__29596\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__5749\ : Odrv12
    port map (
            O => \N__29593\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__5748\ : SRMux
    port map (
            O => \N__29586\,
            I => \N__29583\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__29583\,
            I => \N__29580\
        );

    \I__5746\ : Span4Mux_v
    port map (
            O => \N__29580\,
            I => \N__29577\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__29577\,
            I => \N__29574\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__29574\,
            I => \c0.n8_adj_2327\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__5742\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__29565\,
            I => \N__29561\
        );

    \I__5740\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29555\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__29561\,
            I => \N__29552\
        );

    \I__5738\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29549\
        );

    \I__5737\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29546\
        );

    \I__5736\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29543\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__29555\,
            I => \N__29539\
        );

    \I__5734\ : Span4Mux_h
    port map (
            O => \N__29552\,
            I => \N__29534\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__29549\,
            I => \N__29534\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__29546\,
            I => \N__29529\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__29543\,
            I => \N__29529\
        );

    \I__5730\ : InMux
    port map (
            O => \N__29542\,
            I => \N__29526\
        );

    \I__5729\ : Span4Mux_v
    port map (
            O => \N__29539\,
            I => \N__29523\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__29534\,
            I => \N__29520\
        );

    \I__5727\ : Span4Mux_h
    port map (
            O => \N__29529\,
            I => \N__29517\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__29526\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__29523\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__29520\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__29517\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__5722\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__29502\,
            I => \N__29499\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__29499\,
            I => \c0.n10161\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__29496\,
            I => \n2061_cascade_\
        );

    \I__5717\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__29490\,
            I => \c0.n47_adj_2347\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__29487\,
            I => \c0.n9334_cascade_\
        );

    \I__5714\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__29481\,
            I => \c0.n4\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__29478\,
            I => \c0.n15821_cascade_\
        );

    \I__5711\ : SRMux
    port map (
            O => \N__29475\,
            I => \N__29472\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__29472\,
            I => \N__29469\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__29463\,
            I => \c0.n8_adj_2335\
        );

    \I__5706\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29455\
        );

    \I__5705\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29450\
        );

    \I__5704\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29447\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__29455\,
            I => \N__29444\
        );

    \I__5702\ : InMux
    port map (
            O => \N__29454\,
            I => \N__29441\
        );

    \I__5701\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29438\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29435\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29432\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__29444\,
            I => \N__29428\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29425\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__29438\,
            I => \N__29420\
        );

    \I__5695\ : Span4Mux_v
    port map (
            O => \N__29435\,
            I => \N__29420\
        );

    \I__5694\ : Span12Mux_h
    port map (
            O => \N__29432\,
            I => \N__29417\
        );

    \I__5693\ : InMux
    port map (
            O => \N__29431\,
            I => \N__29414\
        );

    \I__5692\ : Span4Mux_h
    port map (
            O => \N__29428\,
            I => \N__29411\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__29425\,
            I => rand_data_0
        );

    \I__5690\ : Odrv4
    port map (
            O => \N__29420\,
            I => rand_data_0
        );

    \I__5689\ : Odrv12
    port map (
            O => \N__29417\,
            I => rand_data_0
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__29414\,
            I => rand_data_0
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__29411\,
            I => rand_data_0
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__29400\,
            I => \n63_cascade_\
        );

    \I__5685\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__29394\,
            I => \N__29388\
        );

    \I__5683\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29381\
        );

    \I__5682\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29381\
        );

    \I__5681\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29381\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__29388\,
            I => data_in_2_7
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__29381\,
            I => data_in_2_7
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__29376\,
            I => \N__29372\
        );

    \I__5677\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29369\
        );

    \I__5676\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29366\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__29369\,
            I => \N__29361\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29361\
        );

    \I__5673\ : Span4Mux_v
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__29358\,
            I => \c0.n10141\
        );

    \I__5671\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29352\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__29352\,
            I => \c0.n10027\
        );

    \I__5669\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__29343\,
            I => \N__29340\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__29340\,
            I => \c0.n17_adj_2370\
        );

    \I__5665\ : CascadeMux
    port map (
            O => \N__29337\,
            I => \c0.n16_adj_2366_cascade_\
        );

    \I__5664\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29330\
        );

    \I__5663\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29325\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__29330\,
            I => \N__29322\
        );

    \I__5661\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29317\
        );

    \I__5660\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29317\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__29325\,
            I => data_in_1_7
        );

    \I__5658\ : Odrv12
    port map (
            O => \N__29322\,
            I => data_in_1_7
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__29317\,
            I => data_in_1_7
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__29310\,
            I => \n9378_cascade_\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__29307\,
            I => \c0.n47_adj_2347_cascade_\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__29304\,
            I => \c0.n13146_cascade_\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__29301\,
            I => \N__29297\
        );

    \I__5652\ : CascadeMux
    port map (
            O => \N__29300\,
            I => \N__29294\
        );

    \I__5651\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29291\
        );

    \I__5650\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29288\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__29291\,
            I => \N__29285\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__29288\,
            I => \c0.data_in_frame_3_4\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__29285\,
            I => \c0.data_in_frame_3_4\
        );

    \I__5646\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29275\
        );

    \I__5645\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29270\
        );

    \I__5644\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29270\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__29275\,
            I => data_in_0_1
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__29270\,
            I => data_in_0_1
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__29265\,
            I => \c0.n7_adj_2384_cascade_\
        );

    \I__5640\ : SRMux
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__29256\,
            I => \c0.n6_adj_2336\
        );

    \I__5637\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29249\
        );

    \I__5636\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29246\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__29249\,
            I => \c0.n10136\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__29246\,
            I => \c0.n10136\
        );

    \I__5633\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29237\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__29240\,
            I => \N__29234\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__29237\,
            I => \N__29229\
        );

    \I__5630\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29226\
        );

    \I__5629\ : InMux
    port map (
            O => \N__29233\,
            I => \N__29221\
        );

    \I__5628\ : InMux
    port map (
            O => \N__29232\,
            I => \N__29221\
        );

    \I__5627\ : Odrv12
    port map (
            O => \N__29229\,
            I => data_in_1_4
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__29226\,
            I => data_in_1_4
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__29221\,
            I => data_in_1_4
        );

    \I__5624\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29206\
        );

    \I__5623\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29206\
        );

    \I__5622\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29203\
        );

    \I__5621\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29200\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__29206\,
            I => data_in_2_3
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__29203\,
            I => data_in_2_3
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__29200\,
            I => data_in_2_3
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__29193\,
            I => \c0.n16_adj_2361_cascade_\
        );

    \I__5616\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29187\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__29187\,
            I => \c0.n17_adj_2362\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__29184\,
            I => \n17075_cascade_\
        );

    \I__5613\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29177\
        );

    \I__5612\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29172\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29169\
        );

    \I__5610\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29166\
        );

    \I__5609\ : InMux
    port map (
            O => \N__29175\,
            I => \N__29163\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__29172\,
            I => data_in_2_5
        );

    \I__5607\ : Odrv12
    port map (
            O => \N__29169\,
            I => data_in_2_5
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__29166\,
            I => data_in_2_5
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__29163\,
            I => data_in_2_5
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__29154\,
            I => \N__29150\
        );

    \I__5603\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29144\
        );

    \I__5602\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29144\
        );

    \I__5601\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29141\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__29144\,
            I => \N__29135\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29135\
        );

    \I__5598\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29132\
        );

    \I__5597\ : Span4Mux_v
    port map (
            O => \N__29135\,
            I => \N__29129\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__29132\,
            I => data_in_2_0
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__29129\,
            I => data_in_2_0
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__29124\,
            I => \c0.n17400_cascade_\
        );

    \I__5593\ : CascadeMux
    port map (
            O => \N__29121\,
            I => \c0.n8_adj_2359_cascade_\
        );

    \I__5592\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__29115\,
            I => \c0.n13450\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__29112\,
            I => \c0.n15_adj_2310_cascade_\
        );

    \I__5589\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29105\
        );

    \I__5588\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29102\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__29105\,
            I => \c0.data_in_frame_3_3\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__29102\,
            I => \c0.data_in_frame_3_3\
        );

    \I__5585\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29094\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__29094\,
            I => \c0.n17659\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__29091\,
            I => \c0.n11867_cascade_\
        );

    \I__5582\ : SRMux
    port map (
            O => \N__29088\,
            I => \N__29085\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__29085\,
            I => \N__29082\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__29082\,
            I => \c0.n4_adj_2187\
        );

    \I__5579\ : SRMux
    port map (
            O => \N__29079\,
            I => \N__29076\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__29076\,
            I => \c0.n4_adj_2152\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__5576\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29067\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__29067\,
            I => \N__29063\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__29066\,
            I => \N__29060\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__29063\,
            I => \N__29044\
        );

    \I__5572\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29041\
        );

    \I__5571\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29036\
        );

    \I__5570\ : InMux
    port map (
            O => \N__29058\,
            I => \N__29036\
        );

    \I__5569\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29033\
        );

    \I__5568\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29028\
        );

    \I__5567\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29028\
        );

    \I__5566\ : InMux
    port map (
            O => \N__29054\,
            I => \N__29025\
        );

    \I__5565\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29019\
        );

    \I__5564\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29014\
        );

    \I__5563\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29014\
        );

    \I__5562\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29009\
        );

    \I__5561\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29009\
        );

    \I__5560\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29000\
        );

    \I__5559\ : InMux
    port map (
            O => \N__29047\,
            I => \N__28994\
        );

    \I__5558\ : Span4Mux_h
    port map (
            O => \N__29044\,
            I => \N__28989\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__29041\,
            I => \N__28989\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__28986\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__29033\,
            I => \N__28981\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__29028\,
            I => \N__28981\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__29025\,
            I => \N__28978\
        );

    \I__5552\ : InMux
    port map (
            O => \N__29024\,
            I => \N__28973\
        );

    \I__5551\ : InMux
    port map (
            O => \N__29023\,
            I => \N__28973\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__29022\,
            I => \N__28963\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__29019\,
            I => \N__28954\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__28954\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__28951\
        );

    \I__5546\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28944\
        );

    \I__5545\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28944\
        );

    \I__5544\ : InMux
    port map (
            O => \N__29006\,
            I => \N__28944\
        );

    \I__5543\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28939\
        );

    \I__5542\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28939\
        );

    \I__5541\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28935\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__29000\,
            I => \N__28929\
        );

    \I__5539\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28926\
        );

    \I__5538\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28920\
        );

    \I__5537\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28917\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__28994\,
            I => \N__28914\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__28989\,
            I => \N__28911\
        );

    \I__5534\ : Span4Mux_s2_h
    port map (
            O => \N__28986\,
            I => \N__28902\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__28981\,
            I => \N__28902\
        );

    \I__5532\ : Span4Mux_v
    port map (
            O => \N__28978\,
            I => \N__28902\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__28973\,
            I => \N__28902\
        );

    \I__5530\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28896\
        );

    \I__5529\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28896\
        );

    \I__5528\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28893\
        );

    \I__5527\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28888\
        );

    \I__5526\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28881\
        );

    \I__5525\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28881\
        );

    \I__5524\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28881\
        );

    \I__5523\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28878\
        );

    \I__5522\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28873\
        );

    \I__5521\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28873\
        );

    \I__5520\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28870\
        );

    \I__5519\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28867\
        );

    \I__5518\ : Span4Mux_v
    port map (
            O => \N__28954\,
            I => \N__28862\
        );

    \I__5517\ : Span4Mux_h
    port map (
            O => \N__28951\,
            I => \N__28862\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28857\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__28939\,
            I => \N__28857\
        );

    \I__5514\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28854\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__28935\,
            I => \N__28851\
        );

    \I__5512\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28846\
        );

    \I__5511\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28846\
        );

    \I__5510\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28843\
        );

    \I__5509\ : Span4Mux_s2_h
    port map (
            O => \N__28929\,
            I => \N__28838\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__28926\,
            I => \N__28838\
        );

    \I__5507\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28831\
        );

    \I__5506\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28831\
        );

    \I__5505\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28831\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__28920\,
            I => \N__28826\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__28917\,
            I => \N__28826\
        );

    \I__5502\ : Span4Mux_v
    port map (
            O => \N__28914\,
            I => \N__28819\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__28911\,
            I => \N__28819\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__28902\,
            I => \N__28819\
        );

    \I__5499\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28813\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__28896\,
            I => \N__28808\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28808\
        );

    \I__5496\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28803\
        );

    \I__5495\ : InMux
    port map (
            O => \N__28891\,
            I => \N__28803\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__28888\,
            I => \N__28794\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28794\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28794\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28794\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28791\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28784\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__28862\,
            I => \N__28784\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__28857\,
            I => \N__28784\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__28854\,
            I => \N__28776\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__28851\,
            I => \N__28776\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__28846\,
            I => \N__28776\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__28843\,
            I => \N__28773\
        );

    \I__5482\ : Span4Mux_h
    port map (
            O => \N__28838\,
            I => \N__28764\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__28831\,
            I => \N__28764\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__28826\,
            I => \N__28764\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__28819\,
            I => \N__28764\
        );

    \I__5478\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28757\
        );

    \I__5477\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28757\
        );

    \I__5476\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28757\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__28813\,
            I => \N__28748\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__28808\,
            I => \N__28748\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28748\
        );

    \I__5472\ : Span4Mux_h
    port map (
            O => \N__28794\,
            I => \N__28748\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__28791\,
            I => \N__28743\
        );

    \I__5470\ : Span4Mux_h
    port map (
            O => \N__28784\,
            I => \N__28743\
        );

    \I__5469\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28740\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__28776\,
            I => \N__28735\
        );

    \I__5467\ : Span4Mux_h
    port map (
            O => \N__28773\,
            I => \N__28735\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__28764\,
            I => \N__28732\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28725\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__28748\,
            I => \N__28725\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__28743\,
            I => \N__28725\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__28740\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__28735\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__28732\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__28725\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__5458\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__5456\ : Span4Mux_h
    port map (
            O => \N__28710\,
            I => \N__28707\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__28707\,
            I => \N__28704\
        );

    \I__5454\ : Odrv4
    port map (
            O => \N__28704\,
            I => \c0.n17761\
        );

    \I__5453\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28696\
        );

    \I__5452\ : InMux
    port map (
            O => \N__28700\,
            I => \N__28689\
        );

    \I__5451\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28689\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__28696\,
            I => \N__28686\
        );

    \I__5449\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28680\
        );

    \I__5448\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28677\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__28689\,
            I => \N__28672\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__28686\,
            I => \N__28669\
        );

    \I__5445\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28664\
        );

    \I__5444\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28664\
        );

    \I__5443\ : CascadeMux
    port map (
            O => \N__28683\,
            I => \N__28656\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28642\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__28677\,
            I => \N__28642\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__28676\,
            I => \N__28633\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__28675\,
            I => \N__28628\
        );

    \I__5438\ : Span4Mux_v
    port map (
            O => \N__28672\,
            I => \N__28621\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__28669\,
            I => \N__28621\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__28664\,
            I => \N__28621\
        );

    \I__5435\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28616\
        );

    \I__5434\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28616\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__28661\,
            I => \N__28607\
        );

    \I__5432\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28602\
        );

    \I__5431\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28602\
        );

    \I__5430\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28591\
        );

    \I__5429\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28591\
        );

    \I__5428\ : CascadeMux
    port map (
            O => \N__28654\,
            I => \N__28586\
        );

    \I__5427\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28580\
        );

    \I__5426\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28580\
        );

    \I__5425\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28577\
        );

    \I__5424\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28572\
        );

    \I__5423\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28572\
        );

    \I__5422\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28567\
        );

    \I__5421\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28567\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__28642\,
            I => \N__28564\
        );

    \I__5419\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28561\
        );

    \I__5418\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28556\
        );

    \I__5417\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28556\
        );

    \I__5416\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28551\
        );

    \I__5415\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28551\
        );

    \I__5414\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28539\
        );

    \I__5413\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28539\
        );

    \I__5412\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28539\
        );

    \I__5411\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28534\
        );

    \I__5410\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28534\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__28621\,
            I => \N__28531\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__28616\,
            I => \N__28528\
        );

    \I__5407\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28523\
        );

    \I__5406\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28523\
        );

    \I__5405\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28520\
        );

    \I__5404\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28517\
        );

    \I__5403\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28510\
        );

    \I__5402\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28510\
        );

    \I__5401\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28510\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__28602\,
            I => \N__28507\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__28601\,
            I => \N__28500\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__28600\,
            I => \N__28494\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__28599\,
            I => \N__28490\
        );

    \I__5396\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28487\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \N__28484\
        );

    \I__5394\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28480\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__28591\,
            I => \N__28477\
        );

    \I__5392\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28474\
        );

    \I__5391\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28469\
        );

    \I__5390\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28469\
        );

    \I__5389\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28466\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28462\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__28577\,
            I => \N__28455\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28455\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__28567\,
            I => \N__28455\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__28564\,
            I => \N__28450\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__28561\,
            I => \N__28450\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__28556\,
            I => \N__28442\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28442\
        );

    \I__5380\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28431\
        );

    \I__5379\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28431\
        );

    \I__5378\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28431\
        );

    \I__5377\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28431\
        );

    \I__5376\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28431\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28426\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28426\
        );

    \I__5373\ : IoSpan4Mux
    port map (
            O => \N__28531\,
            I => \N__28423\
        );

    \I__5372\ : Span4Mux_v
    port map (
            O => \N__28528\,
            I => \N__28420\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__28523\,
            I => \N__28411\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__28520\,
            I => \N__28411\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__28517\,
            I => \N__28411\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__28510\,
            I => \N__28411\
        );

    \I__5367\ : Span4Mux_v
    port map (
            O => \N__28507\,
            I => \N__28408\
        );

    \I__5366\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28401\
        );

    \I__5365\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28401\
        );

    \I__5364\ : InMux
    port map (
            O => \N__28504\,
            I => \N__28401\
        );

    \I__5363\ : InMux
    port map (
            O => \N__28503\,
            I => \N__28394\
        );

    \I__5362\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28394\
        );

    \I__5361\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28394\
        );

    \I__5360\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28387\
        );

    \I__5359\ : InMux
    port map (
            O => \N__28497\,
            I => \N__28387\
        );

    \I__5358\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28387\
        );

    \I__5357\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28384\
        );

    \I__5356\ : InMux
    port map (
            O => \N__28490\,
            I => \N__28381\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__28487\,
            I => \N__28378\
        );

    \I__5354\ : InMux
    port map (
            O => \N__28484\,
            I => \N__28373\
        );

    \I__5353\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28373\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__28480\,
            I => \N__28368\
        );

    \I__5351\ : Span4Mux_s3_h
    port map (
            O => \N__28477\,
            I => \N__28368\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28363\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28363\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__28466\,
            I => \N__28357\
        );

    \I__5347\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28354\
        );

    \I__5346\ : Span4Mux_h
    port map (
            O => \N__28462\,
            I => \N__28347\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__28455\,
            I => \N__28347\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__28450\,
            I => \N__28347\
        );

    \I__5343\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28340\
        );

    \I__5342\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28340\
        );

    \I__5341\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28340\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__28442\,
            I => \N__28329\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__28431\,
            I => \N__28329\
        );

    \I__5338\ : Span4Mux_v
    port map (
            O => \N__28426\,
            I => \N__28329\
        );

    \I__5337\ : Span4Mux_s2_h
    port map (
            O => \N__28423\,
            I => \N__28329\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__28420\,
            I => \N__28329\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__28411\,
            I => \N__28314\
        );

    \I__5334\ : Span4Mux_h
    port map (
            O => \N__28408\,
            I => \N__28314\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__28401\,
            I => \N__28314\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__28394\,
            I => \N__28314\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__28387\,
            I => \N__28314\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__28384\,
            I => \N__28314\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__28381\,
            I => \N__28314\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__28378\,
            I => \N__28305\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28305\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__28368\,
            I => \N__28305\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__28363\,
            I => \N__28305\
        );

    \I__5324\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28302\
        );

    \I__5323\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28299\
        );

    \I__5322\ : InMux
    port map (
            O => \N__28360\,
            I => \N__28296\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__28357\,
            I => \N__28293\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__28354\,
            I => \N__28288\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__28347\,
            I => \N__28288\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28281\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__28329\,
            I => \N__28281\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__28314\,
            I => \N__28281\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__28305\,
            I => \N__28278\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__28302\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__28299\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__28296\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__28293\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__28288\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__28281\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__28278\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__5307\ : SRMux
    port map (
            O => \N__28263\,
            I => \N__28260\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__28260\,
            I => \c0.n4_adj_2155\
        );

    \I__5305\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28251\
        );

    \I__5304\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28251\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__28251\,
            I => \c0.data_in_frame_3_6\
        );

    \I__5302\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__28245\,
            I => n7
        );

    \I__5300\ : InMux
    port map (
            O => \N__28242\,
            I => n16059
        );

    \I__5299\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28236\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__28236\,
            I => n6_adj_2429
        );

    \I__5297\ : InMux
    port map (
            O => \N__28233\,
            I => n16060
        );

    \I__5296\ : InMux
    port map (
            O => \N__28230\,
            I => n16061
        );

    \I__5295\ : InMux
    port map (
            O => \N__28227\,
            I => n16062
        );

    \I__5294\ : InMux
    port map (
            O => \N__28224\,
            I => n16063
        );

    \I__5293\ : InMux
    port map (
            O => \N__28221\,
            I => \bfn_9_32_0_\
        );

    \I__5292\ : InMux
    port map (
            O => \N__28218\,
            I => n16065
        );

    \I__5291\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__28212\,
            I => \c0.n17711\
        );

    \I__5289\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28206\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__28206\,
            I => n15
        );

    \I__5287\ : InMux
    port map (
            O => \N__28203\,
            I => n16051
        );

    \I__5286\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__28197\,
            I => n14
        );

    \I__5284\ : InMux
    port map (
            O => \N__28194\,
            I => n16052
        );

    \I__5283\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28188\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__28188\,
            I => n13
        );

    \I__5281\ : InMux
    port map (
            O => \N__28185\,
            I => n16053
        );

    \I__5280\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28179\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__28179\,
            I => n12
        );

    \I__5278\ : InMux
    port map (
            O => \N__28176\,
            I => n16054
        );

    \I__5277\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__28170\,
            I => n11
        );

    \I__5275\ : InMux
    port map (
            O => \N__28167\,
            I => n16055
        );

    \I__5274\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28161\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__28161\,
            I => n10_adj_2420
        );

    \I__5272\ : InMux
    port map (
            O => \N__28158\,
            I => \bfn_9_31_0_\
        );

    \I__5271\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__28152\,
            I => n9_adj_2421
        );

    \I__5269\ : InMux
    port map (
            O => \N__28149\,
            I => n16057
        );

    \I__5268\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28143\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__28143\,
            I => n8_adj_2412
        );

    \I__5266\ : InMux
    port map (
            O => \N__28140\,
            I => n16058
        );

    \I__5265\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__28134\,
            I => n24
        );

    \I__5263\ : InMux
    port map (
            O => \N__28131\,
            I => n16042
        );

    \I__5262\ : InMux
    port map (
            O => \N__28128\,
            I => \N__28125\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__28125\,
            I => n23_adj_2425
        );

    \I__5260\ : InMux
    port map (
            O => \N__28122\,
            I => n16043
        );

    \I__5259\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__28116\,
            I => n22_adj_2426
        );

    \I__5257\ : InMux
    port map (
            O => \N__28113\,
            I => n16044
        );

    \I__5256\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__28107\,
            I => n21
        );

    \I__5254\ : InMux
    port map (
            O => \N__28104\,
            I => n16045
        );

    \I__5253\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28098\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__28098\,
            I => n20
        );

    \I__5251\ : InMux
    port map (
            O => \N__28095\,
            I => n16046
        );

    \I__5250\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28089\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__28089\,
            I => n19
        );

    \I__5248\ : InMux
    port map (
            O => \N__28086\,
            I => n16047
        );

    \I__5247\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__28080\,
            I => n18
        );

    \I__5245\ : InMux
    port map (
            O => \N__28077\,
            I => \bfn_9_30_0_\
        );

    \I__5244\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28071\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__28071\,
            I => n17
        );

    \I__5242\ : InMux
    port map (
            O => \N__28068\,
            I => n16049
        );

    \I__5241\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28062\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__28062\,
            I => n16
        );

    \I__5239\ : InMux
    port map (
            O => \N__28059\,
            I => n16050
        );

    \I__5238\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28049\
        );

    \I__5237\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28049\
        );

    \I__5236\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28045\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__28049\,
            I => \N__28042\
        );

    \I__5234\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28039\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__28045\,
            I => \N__28034\
        );

    \I__5232\ : Span12Mux_s5_v
    port map (
            O => \N__28042\,
            I => \N__28034\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__28039\,
            I => data_in_1_2
        );

    \I__5230\ : Odrv12
    port map (
            O => \N__28034\,
            I => data_in_1_2
        );

    \I__5229\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28026\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28023\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__28020\,
            I => \c0.n17388\
        );

    \I__5225\ : SRMux
    port map (
            O => \N__28017\,
            I => \N__28014\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__28014\,
            I => \N__28011\
        );

    \I__5223\ : Span4Mux_h
    port map (
            O => \N__28011\,
            I => \N__28008\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__28008\,
            I => \c0.n3_adj_2272\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__5220\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27997\
        );

    \I__5219\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27993\
        );

    \I__5218\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27990\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27987\
        );

    \I__5216\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27984\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27979\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27979\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__27987\,
            I => \N__27974\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27974\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__27979\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__27974\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__5209\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27966\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N__27963\
        );

    \I__5207\ : Span4Mux_h
    port map (
            O => \N__27963\,
            I => \N__27960\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__27960\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_10\
        );

    \I__5205\ : SRMux
    port map (
            O => \N__27957\,
            I => \N__27954\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__27954\,
            I => \N__27951\
        );

    \I__5203\ : Span4Mux_s1_h
    port map (
            O => \N__27951\,
            I => \N__27948\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__27948\,
            I => \N__27945\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__27945\,
            I => \c0.n3_adj_2264\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__27942\,
            I => \N__27938\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__27941\,
            I => \N__27934\
        );

    \I__5198\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27929\
        );

    \I__5197\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27929\
        );

    \I__5196\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27925\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27922\
        );

    \I__5194\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27919\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__27925\,
            I => \N__27916\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__27922\,
            I => \N__27911\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__27919\,
            I => \N__27911\
        );

    \I__5190\ : Span4Mux_v
    port map (
            O => \N__27916\,
            I => \N__27906\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__27911\,
            I => \N__27906\
        );

    \I__5188\ : Span4Mux_h
    port map (
            O => \N__27906\,
            I => \N__27903\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__27903\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__5186\ : InMux
    port map (
            O => \N__27900\,
            I => \N__27897\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__27897\,
            I => \N__27894\
        );

    \I__5184\ : Odrv12
    port map (
            O => \N__27894\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_14\
        );

    \I__5183\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27886\
        );

    \I__5182\ : CascadeMux
    port map (
            O => \N__27890\,
            I => \N__27883\
        );

    \I__5181\ : InMux
    port map (
            O => \N__27889\,
            I => \N__27880\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27877\
        );

    \I__5179\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27874\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__27880\,
            I => \N__27870\
        );

    \I__5177\ : Span4Mux_h
    port map (
            O => \N__27877\,
            I => \N__27867\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__27874\,
            I => \N__27864\
        );

    \I__5175\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27861\
        );

    \I__5174\ : Span4Mux_v
    port map (
            O => \N__27870\,
            I => \N__27858\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__27867\,
            I => \N__27855\
        );

    \I__5172\ : Span4Mux_v
    port map (
            O => \N__27864\,
            I => \N__27852\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__27861\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__27858\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__27855\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__27852\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__5167\ : CascadeMux
    port map (
            O => \N__27843\,
            I => \N__27836\
        );

    \I__5166\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27823\
        );

    \I__5165\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27823\
        );

    \I__5164\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27823\
        );

    \I__5163\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27813\
        );

    \I__5162\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27808\
        );

    \I__5161\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27808\
        );

    \I__5160\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27805\
        );

    \I__5159\ : CascadeMux
    port map (
            O => \N__27833\,
            I => \N__27802\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__27832\,
            I => \N__27790\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__27831\,
            I => \N__27787\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__27830\,
            I => \N__27783\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__27823\,
            I => \N__27777\
        );

    \I__5154\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27770\
        );

    \I__5153\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27770\
        );

    \I__5152\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27770\
        );

    \I__5151\ : InMux
    port map (
            O => \N__27819\,
            I => \N__27761\
        );

    \I__5150\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27761\
        );

    \I__5149\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27761\
        );

    \I__5148\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27761\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__27813\,
            I => \N__27756\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__27808\,
            I => \N__27756\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__27805\,
            I => \N__27753\
        );

    \I__5144\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27748\
        );

    \I__5143\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27748\
        );

    \I__5142\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27739\
        );

    \I__5141\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27739\
        );

    \I__5140\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27739\
        );

    \I__5139\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27739\
        );

    \I__5138\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27730\
        );

    \I__5137\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27730\
        );

    \I__5136\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27730\
        );

    \I__5135\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27730\
        );

    \I__5134\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27721\
        );

    \I__5133\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27721\
        );

    \I__5132\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27721\
        );

    \I__5131\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27721\
        );

    \I__5130\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27714\
        );

    \I__5129\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27714\
        );

    \I__5128\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27714\
        );

    \I__5127\ : Span12Mux_s3_h
    port map (
            O => \N__27777\,
            I => \N__27709\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__27770\,
            I => \N__27709\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27702\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__27756\,
            I => \N__27702\
        );

    \I__5123\ : Span4Mux_v
    port map (
            O => \N__27753\,
            I => \N__27702\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__27748\,
            I => \c0.n10009\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__27739\,
            I => \c0.n10009\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__27730\,
            I => \c0.n10009\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__27721\,
            I => \c0.n10009\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__27714\,
            I => \c0.n10009\
        );

    \I__5117\ : Odrv12
    port map (
            O => \N__27709\,
            I => \c0.n10009\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__27702\,
            I => \c0.n10009\
        );

    \I__5115\ : SRMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__5113\ : Span4Mux_h
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__27678\,
            I => \c0.n3_adj_2259\
        );

    \I__5111\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__27672\,
            I => n26_adj_2423
        );

    \I__5109\ : InMux
    port map (
            O => \N__27669\,
            I => \bfn_9_29_0_\
        );

    \I__5108\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27663\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__27663\,
            I => n25_adj_2424
        );

    \I__5106\ : InMux
    port map (
            O => \N__27660\,
            I => n16041
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__27657\,
            I => \N__27652\
        );

    \I__5104\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27649\
        );

    \I__5103\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27645\
        );

    \I__5102\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27642\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__27649\,
            I => \N__27639\
        );

    \I__5100\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27636\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27632\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27627\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__27639\,
            I => \N__27627\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27624\
        );

    \I__5095\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27621\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__27632\,
            I => \N__27616\
        );

    \I__5093\ : Span4Mux_h
    port map (
            O => \N__27627\,
            I => \N__27616\
        );

    \I__5092\ : Span12Mux_s5_h
    port map (
            O => \N__27624\,
            I => \N__27613\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__27621\,
            I => data_out_frame2_16_7
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__27616\,
            I => data_out_frame2_16_7
        );

    \I__5089\ : Odrv12
    port map (
            O => \N__27613\,
            I => data_out_frame2_16_7
        );

    \I__5088\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27603\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__27603\,
            I => \N__27600\
        );

    \I__5086\ : Span4Mux_v
    port map (
            O => \N__27600\,
            I => \N__27597\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__27597\,
            I => \N__27592\
        );

    \I__5084\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27589\
        );

    \I__5083\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27586\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__27592\,
            I => \c0.n17194\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__27589\,
            I => \c0.n17194\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__27586\,
            I => \c0.n17194\
        );

    \I__5079\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27576\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__27576\,
            I => \N__27573\
        );

    \I__5077\ : Span4Mux_h
    port map (
            O => \N__27573\,
            I => \N__27570\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__27570\,
            I => \c0.n10459\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__27567\,
            I => \N__27563\
        );

    \I__5074\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27557\
        );

    \I__5073\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27557\
        );

    \I__5072\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27554\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__27557\,
            I => \N__27551\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__27554\,
            I => data_in_0_5
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__27551\,
            I => data_in_0_5
        );

    \I__5068\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27542\
        );

    \I__5067\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27539\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27536\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__27539\,
            I => data_in_0_4
        );

    \I__5064\ : Odrv12
    port map (
            O => \N__27536\,
            I => data_in_0_4
        );

    \I__5063\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27527\
        );

    \I__5062\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27524\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__27527\,
            I => \N__27521\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__27524\,
            I => data_in_0_2
        );

    \I__5059\ : Odrv12
    port map (
            O => \N__27521\,
            I => data_in_0_2
        );

    \I__5058\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27511\
        );

    \I__5057\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27506\
        );

    \I__5056\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27506\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27503\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__27506\,
            I => data_in_1_5
        );

    \I__5053\ : Odrv12
    port map (
            O => \N__27503\,
            I => data_in_1_5
        );

    \I__5052\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27495\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27492\
        );

    \I__5050\ : Span4Mux_h
    port map (
            O => \N__27492\,
            I => \N__27489\
        );

    \I__5049\ : Span4Mux_h
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__27486\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_16\
        );

    \I__5047\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27478\
        );

    \I__5046\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27475\
        );

    \I__5045\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27472\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__27478\,
            I => \N__27467\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__27475\,
            I => \N__27467\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__27472\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__27467\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__5040\ : SRMux
    port map (
            O => \N__27462\,
            I => \N__27459\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__27459\,
            I => \N__27456\
        );

    \I__5038\ : Odrv12
    port map (
            O => \N__27456\,
            I => \c0.n16716\
        );

    \I__5037\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27444\
        );

    \I__5036\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27444\
        );

    \I__5035\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27444\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__27444\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__5033\ : SRMux
    port map (
            O => \N__27441\,
            I => \N__27438\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__27438\,
            I => \N__27435\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__27435\,
            I => \c0.n8_adj_2332\
        );

    \I__5030\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27425\
        );

    \I__5029\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27425\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__27430\,
            I => \N__27422\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__27425\,
            I => \N__27419\
        );

    \I__5026\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27416\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__27419\,
            I => \N__27413\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__27416\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__27413\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__5022\ : SRMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__27405\,
            I => \N__27402\
        );

    \I__5020\ : Span4Mux_h
    port map (
            O => \N__27402\,
            I => \N__27399\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__27399\,
            I => \c0.n8_adj_2328\
        );

    \I__5018\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27392\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__27395\,
            I => \N__27388\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__27392\,
            I => \N__27385\
        );

    \I__5015\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27382\
        );

    \I__5014\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27379\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__27385\,
            I => \N__27374\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__27382\,
            I => \N__27374\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__27379\,
            I => \N__27371\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__27374\,
            I => \N__27368\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__27371\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__27368\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__5007\ : SRMux
    port map (
            O => \N__27363\,
            I => \N__27360\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__27357\,
            I => \N__27354\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__27354\,
            I => \c0.n8_adj_2334\
        );

    \I__5003\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27348\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__27348\,
            I => \N__27343\
        );

    \I__5001\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27338\
        );

    \I__5000\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27338\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__27343\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__27338\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__4997\ : SRMux
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27327\
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__27327\,
            I => \c0.n16708\
        );

    \I__4994\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27319\
        );

    \I__4993\ : InMux
    port map (
            O => \N__27323\,
            I => \N__27316\
        );

    \I__4992\ : CascadeMux
    port map (
            O => \N__27322\,
            I => \N__27313\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__27319\,
            I => \N__27308\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__27316\,
            I => \N__27308\
        );

    \I__4989\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27305\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__27308\,
            I => \N__27302\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__27305\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__27302\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__4985\ : SRMux
    port map (
            O => \N__27297\,
            I => \N__27294\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__27294\,
            I => \N__27291\
        );

    \I__4983\ : Span4Mux_h
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__27288\,
            I => \N__27285\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__27285\,
            I => \c0.n8_adj_2331\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__27282\,
            I => \N__27278\
        );

    \I__4979\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27272\
        );

    \I__4978\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27272\
        );

    \I__4977\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27269\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__27272\,
            I => data_in_0_6
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__27269\,
            I => data_in_0_6
        );

    \I__4974\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27260\
        );

    \I__4973\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27255\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27252\
        );

    \I__4971\ : InMux
    port map (
            O => \N__27259\,
            I => \N__27249\
        );

    \I__4970\ : InMux
    port map (
            O => \N__27258\,
            I => \N__27246\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__27255\,
            I => \N__27243\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__27252\,
            I => \N__27240\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__27249\,
            I => \N__27235\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__27246\,
            I => \N__27235\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__27243\,
            I => \N__27232\
        );

    \I__4964\ : Span4Mux_h
    port map (
            O => \N__27240\,
            I => \N__27227\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__27235\,
            I => \N__27227\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__27232\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__27227\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__4960\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27219\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__4958\ : Span12Mux_s8_v
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__4957\ : Odrv12
    port map (
            O => \N__27213\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_15\
        );

    \I__4956\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27203\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \N__27199\
        );

    \I__4953\ : Span4Mux_h
    port map (
            O => \N__27203\,
            I => \N__27195\
        );

    \I__4952\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27192\
        );

    \I__4951\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27189\
        );

    \I__4950\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27186\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__27195\,
            I => \N__27179\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27179\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__27189\,
            I => \N__27179\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__27186\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__27179\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__4944\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27168\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__27165\,
            I => \N__27162\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__27162\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_13\
        );

    \I__4939\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27155\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27152\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__27155\,
            I => \N__27148\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__27152\,
            I => \N__27144\
        );

    \I__4935\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27141\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__27148\,
            I => \N__27138\
        );

    \I__4933\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27135\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__27144\,
            I => \N__27132\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__27141\,
            I => \N__27125\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__27138\,
            I => \N__27125\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__27135\,
            I => \N__27125\
        );

    \I__4928\ : Span4Mux_s0_h
    port map (
            O => \N__27132\,
            I => \N__27122\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__27125\,
            I => \N__27119\
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__27122\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__27119\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__4924\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27111\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__27102\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_11\
        );

    \I__4919\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__27096\,
            I => \N__27092\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__27095\,
            I => \N__27089\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__27092\,
            I => \N__27086\
        );

    \I__4915\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27083\
        );

    \I__4914\ : Span4Mux_h
    port map (
            O => \N__27086\,
            I => \N__27078\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27075\
        );

    \I__4912\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27070\
        );

    \I__4911\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27070\
        );

    \I__4910\ : Odrv4
    port map (
            O => \N__27078\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__27075\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__27070\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__4907\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27060\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__27060\,
            I => \N__27057\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__27057\,
            I => \N__27054\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__27054\,
            I => \N__27051\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__27051\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_7\
        );

    \I__4902\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27045\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__27045\,
            I => \N__27042\
        );

    \I__4900\ : Span4Mux_h
    port map (
            O => \N__27042\,
            I => \N__27039\
        );

    \I__4899\ : Span4Mux_h
    port map (
            O => \N__27039\,
            I => \N__27036\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__27036\,
            I => \c0.n37\
        );

    \I__4897\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27027\
        );

    \I__4895\ : Span4Mux_h
    port map (
            O => \N__27027\,
            I => \N__27021\
        );

    \I__4894\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27016\
        );

    \I__4893\ : InMux
    port map (
            O => \N__27025\,
            I => \N__27016\
        );

    \I__4892\ : InMux
    port map (
            O => \N__27024\,
            I => \N__27013\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__27021\,
            I => \N__27008\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__27016\,
            I => \N__27008\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__27005\
        );

    \I__4888\ : Span4Mux_h
    port map (
            O => \N__27008\,
            I => \N__27002\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__27005\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__27002\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__4885\ : InMux
    port map (
            O => \N__26997\,
            I => \N__26994\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__26994\,
            I => \N__26991\
        );

    \I__4883\ : Sp12to4
    port map (
            O => \N__26991\,
            I => \N__26988\
        );

    \I__4882\ : Span12Mux_s8_h
    port map (
            O => \N__26988\,
            I => \N__26985\
        );

    \I__4881\ : Odrv12
    port map (
            O => \N__26985\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_28\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__26982\,
            I => \c0.n17331_cascade_\
        );

    \I__4879\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26976\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__26976\,
            I => \c0.n17410\
        );

    \I__4877\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26970\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__26970\,
            I => \N__26967\
        );

    \I__4875\ : Span4Mux_s1_v
    port map (
            O => \N__26967\,
            I => \N__26964\
        );

    \I__4874\ : Span4Mux_v
    port map (
            O => \N__26964\,
            I => \N__26959\
        );

    \I__4873\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26956\
        );

    \I__4872\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26953\
        );

    \I__4871\ : Span4Mux_v
    port map (
            O => \N__26959\,
            I => \N__26948\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__26956\,
            I => \N__26948\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__26953\,
            I => data_in_2_6
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__26948\,
            I => data_in_2_6
        );

    \I__4867\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__26940\,
            I => \c0.n12_adj_2355\
        );

    \I__4865\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26932\
        );

    \I__4864\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26927\
        );

    \I__4863\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26927\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__26932\,
            I => data_in_2_4
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__26927\,
            I => data_in_2_4
        );

    \I__4860\ : SRMux
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__4858\ : Odrv12
    port map (
            O => \N__26916\,
            I => \c0.n4_adj_2150\
        );

    \I__4857\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26910\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__26910\,
            I => \c0.n10133\
        );

    \I__4855\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__26904\,
            I => \c0.n17406\
        );

    \I__4853\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26892\
        );

    \I__4852\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26892\
        );

    \I__4851\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26892\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__26892\,
            I => data_in_0_3
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__26889\,
            I => \c0.n10133_cascade_\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \c0.n6_adj_2356_cascade_\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__26883\,
            I => \c0.n10027_cascade_\
        );

    \I__4846\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26876\
        );

    \I__4845\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26873\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__26876\,
            I => data_in_0_7
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__26873\,
            I => data_in_0_7
        );

    \I__4842\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26861\
        );

    \I__4841\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26861\
        );

    \I__4840\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26858\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__26861\,
            I => data_in_1_3
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__26858\,
            I => data_in_1_3
        );

    \I__4837\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26849\
        );

    \I__4836\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26844\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26841\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__26848\,
            I => \N__26836\
        );

    \I__4833\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26833\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__26844\,
            I => \N__26830\
        );

    \I__4831\ : Span4Mux_h
    port map (
            O => \N__26841\,
            I => \N__26827\
        );

    \I__4830\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26823\
        );

    \I__4829\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26820\
        );

    \I__4828\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26815\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__26833\,
            I => \N__26810\
        );

    \I__4826\ : Span4Mux_h
    port map (
            O => \N__26830\,
            I => \N__26810\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__26827\,
            I => \N__26807\
        );

    \I__4824\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26804\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__26823\,
            I => \N__26799\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26799\
        );

    \I__4821\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26794\
        );

    \I__4820\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26794\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__26815\,
            I => \N__26791\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__26810\,
            I => \N__26788\
        );

    \I__4817\ : Span4Mux_v
    port map (
            O => \N__26807\,
            I => \N__26785\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__26804\,
            I => \N__26780\
        );

    \I__4815\ : Span4Mux_h
    port map (
            O => \N__26799\,
            I => \N__26780\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__26794\,
            I => \r_SM_Main_2_adj_2438\
        );

    \I__4813\ : Odrv12
    port map (
            O => \N__26791\,
            I => \r_SM_Main_2_adj_2438\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__26788\,
            I => \r_SM_Main_2_adj_2438\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__26785\,
            I => \r_SM_Main_2_adj_2438\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__26780\,
            I => \r_SM_Main_2_adj_2438\
        );

    \I__4809\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26766\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__26757\,
            I => n4_adj_2484
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__26754\,
            I => \N__26747\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__26753\,
            I => \N__26743\
        );

    \I__4802\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26735\
        );

    \I__4801\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26735\
        );

    \I__4800\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26730\
        );

    \I__4799\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26730\
        );

    \I__4798\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26727\
        );

    \I__4797\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26724\
        );

    \I__4796\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26721\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__26741\,
            I => \N__26717\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__26740\,
            I => \N__26714\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26711\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__26730\,
            I => \N__26708\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__26727\,
            I => \N__26705\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26702\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__26721\,
            I => \N__26699\
        );

    \I__4788\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26696\
        );

    \I__4787\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26691\
        );

    \I__4786\ : InMux
    port map (
            O => \N__26714\,
            I => \N__26691\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__26711\,
            I => \N__26686\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__26708\,
            I => \N__26686\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__26705\,
            I => \N__26679\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__26702\,
            I => \N__26679\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__26699\,
            I => \N__26679\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__26696\,
            I => \r_SM_Main_1_adj_2439\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__26691\,
            I => \r_SM_Main_1_adj_2439\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__26686\,
            I => \r_SM_Main_1_adj_2439\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__26679\,
            I => \r_SM_Main_1_adj_2439\
        );

    \I__4776\ : InMux
    port map (
            O => \N__26670\,
            I => \c0.n15977\
        );

    \I__4775\ : InMux
    port map (
            O => \N__26667\,
            I => \c0.n15978\
        );

    \I__4774\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26661\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__26661\,
            I => \N__26658\
        );

    \I__4772\ : Span4Mux_h
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__26655\,
            I => \c0.n17714\
        );

    \I__4770\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26649\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__26649\,
            I => \c0.n17589\
        );

    \I__4768\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26640\
        );

    \I__4767\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26640\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__26640\,
            I => \N__26636\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__26639\,
            I => \N__26633\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__26636\,
            I => \N__26629\
        );

    \I__4763\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26626\
        );

    \I__4762\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26623\
        );

    \I__4761\ : Sp12to4
    port map (
            O => \N__26629\,
            I => \N__26618\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__26626\,
            I => \N__26618\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__26623\,
            I => data_out_frame2_7_1
        );

    \I__4758\ : Odrv12
    port map (
            O => \N__26618\,
            I => data_out_frame2_7_1
        );

    \I__4757\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26602\
        );

    \I__4756\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26602\
        );

    \I__4755\ : CEMux
    port map (
            O => \N__26611\,
            I => \N__26593\
        );

    \I__4754\ : CEMux
    port map (
            O => \N__26610\,
            I => \N__26590\
        );

    \I__4753\ : CEMux
    port map (
            O => \N__26609\,
            I => \N__26568\
        );

    \I__4752\ : CEMux
    port map (
            O => \N__26608\,
            I => \N__26551\
        );

    \I__4751\ : CEMux
    port map (
            O => \N__26607\,
            I => \N__26548\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__26602\,
            I => \N__26539\
        );

    \I__4749\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26531\
        );

    \I__4748\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26531\
        );

    \I__4747\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26531\
        );

    \I__4746\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26524\
        );

    \I__4745\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26524\
        );

    \I__4744\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26524\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__26593\,
            I => \N__26519\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__26590\,
            I => \N__26519\
        );

    \I__4741\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26501\
        );

    \I__4740\ : InMux
    port map (
            O => \N__26588\,
            I => \N__26501\
        );

    \I__4739\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26501\
        );

    \I__4738\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26494\
        );

    \I__4737\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26494\
        );

    \I__4736\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26494\
        );

    \I__4735\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26491\
        );

    \I__4734\ : InMux
    port map (
            O => \N__26582\,
            I => \N__26484\
        );

    \I__4733\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26484\
        );

    \I__4732\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26484\
        );

    \I__4731\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26475\
        );

    \I__4730\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26475\
        );

    \I__4729\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26475\
        );

    \I__4728\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26475\
        );

    \I__4727\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26464\
        );

    \I__4726\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26464\
        );

    \I__4725\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26464\
        );

    \I__4724\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26464\
        );

    \I__4723\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26464\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__26568\,
            I => \N__26461\
        );

    \I__4721\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26452\
        );

    \I__4720\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26452\
        );

    \I__4719\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26452\
        );

    \I__4718\ : CEMux
    port map (
            O => \N__26564\,
            I => \N__26449\
        );

    \I__4717\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26446\
        );

    \I__4716\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26443\
        );

    \I__4715\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26440\
        );

    \I__4714\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26433\
        );

    \I__4713\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26433\
        );

    \I__4712\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26433\
        );

    \I__4711\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26424\
        );

    \I__4710\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26424\
        );

    \I__4709\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26424\
        );

    \I__4708\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26424\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__26551\,
            I => \N__26419\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__26548\,
            I => \N__26419\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__26547\,
            I => \N__26416\
        );

    \I__4704\ : InMux
    port map (
            O => \N__26546\,
            I => \N__26410\
        );

    \I__4703\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26410\
        );

    \I__4702\ : CEMux
    port map (
            O => \N__26544\,
            I => \N__26407\
        );

    \I__4701\ : CEMux
    port map (
            O => \N__26543\,
            I => \N__26404\
        );

    \I__4700\ : CEMux
    port map (
            O => \N__26542\,
            I => \N__26401\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__26539\,
            I => \N__26398\
        );

    \I__4698\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26395\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__26531\,
            I => \N__26390\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__26524\,
            I => \N__26390\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__26519\,
            I => \N__26387\
        );

    \I__4694\ : CEMux
    port map (
            O => \N__26518\,
            I => \N__26330\
        );

    \I__4693\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26327\
        );

    \I__4692\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26318\
        );

    \I__4691\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26318\
        );

    \I__4690\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26318\
        );

    \I__4689\ : InMux
    port map (
            O => \N__26513\,
            I => \N__26318\
        );

    \I__4688\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26307\
        );

    \I__4687\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26307\
        );

    \I__4686\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26307\
        );

    \I__4685\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26307\
        );

    \I__4684\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26307\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26304\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26301\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__26491\,
            I => \N__26290\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__26484\,
            I => \N__26290\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26290\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__26464\,
            I => \N__26290\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__26461\,
            I => \N__26290\
        );

    \I__4676\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26285\
        );

    \I__4675\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26285\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26282\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26279\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__26446\,
            I => \N__26270\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__26443\,
            I => \N__26270\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26270\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__26433\,
            I => \N__26270\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__26424\,
            I => \N__26265\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__26419\,
            I => \N__26265\
        );

    \I__4666\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26260\
        );

    \I__4665\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26260\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__26410\,
            I => \N__26255\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__26407\,
            I => \N__26255\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26250\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__26401\,
            I => \N__26250\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__26398\,
            I => \N__26241\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__26395\,
            I => \N__26241\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__26390\,
            I => \N__26241\
        );

    \I__4657\ : Span4Mux_s0_h
    port map (
            O => \N__26387\,
            I => \N__26241\
        );

    \I__4656\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26236\
        );

    \I__4655\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26236\
        );

    \I__4654\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26219\
        );

    \I__4653\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26219\
        );

    \I__4652\ : InMux
    port map (
            O => \N__26382\,
            I => \N__26219\
        );

    \I__4651\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26219\
        );

    \I__4650\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26219\
        );

    \I__4649\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26219\
        );

    \I__4648\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26219\
        );

    \I__4647\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26219\
        );

    \I__4646\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26208\
        );

    \I__4645\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26208\
        );

    \I__4644\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26208\
        );

    \I__4643\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26208\
        );

    \I__4642\ : InMux
    port map (
            O => \N__26372\,
            I => \N__26208\
        );

    \I__4641\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26193\
        );

    \I__4640\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26193\
        );

    \I__4639\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26193\
        );

    \I__4638\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26193\
        );

    \I__4637\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26193\
        );

    \I__4636\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26193\
        );

    \I__4635\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26193\
        );

    \I__4634\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26180\
        );

    \I__4633\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26180\
        );

    \I__4632\ : InMux
    port map (
            O => \N__26362\,
            I => \N__26180\
        );

    \I__4631\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26180\
        );

    \I__4630\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26180\
        );

    \I__4629\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26180\
        );

    \I__4628\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26167\
        );

    \I__4627\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26167\
        );

    \I__4626\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26167\
        );

    \I__4625\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26167\
        );

    \I__4624\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26167\
        );

    \I__4623\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26167\
        );

    \I__4622\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26152\
        );

    \I__4621\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26152\
        );

    \I__4620\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26152\
        );

    \I__4619\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26152\
        );

    \I__4618\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26152\
        );

    \I__4617\ : InMux
    port map (
            O => \N__26347\,
            I => \N__26152\
        );

    \I__4616\ : InMux
    port map (
            O => \N__26346\,
            I => \N__26152\
        );

    \I__4615\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26135\
        );

    \I__4614\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26135\
        );

    \I__4613\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26135\
        );

    \I__4612\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26135\
        );

    \I__4611\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26135\
        );

    \I__4610\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26135\
        );

    \I__4609\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26135\
        );

    \I__4608\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26135\
        );

    \I__4607\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26124\
        );

    \I__4606\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26124\
        );

    \I__4605\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26124\
        );

    \I__4604\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26124\
        );

    \I__4603\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26124\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__26330\,
            I => \N__26121\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__26327\,
            I => \N__26118\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__26318\,
            I => \N__26115\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26106\
        );

    \I__4598\ : Span4Mux_s3_h
    port map (
            O => \N__26304\,
            I => \N__26106\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__26301\,
            I => \N__26106\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__26290\,
            I => \N__26106\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26095\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__26282\,
            I => \N__26095\
        );

    \I__4593\ : Span4Mux_v
    port map (
            O => \N__26279\,
            I => \N__26095\
        );

    \I__4592\ : Span4Mux_v
    port map (
            O => \N__26270\,
            I => \N__26095\
        );

    \I__4591\ : Span4Mux_s2_h
    port map (
            O => \N__26265\,
            I => \N__26095\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__26260\,
            I => \N__26086\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26086\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__26250\,
            I => \N__26086\
        );

    \I__4587\ : Span4Mux_h
    port map (
            O => \N__26241\,
            I => \N__26086\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__26236\,
            I => n10725
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__26219\,
            I => n10725
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__26208\,
            I => n10725
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__26193\,
            I => n10725
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__26180\,
            I => n10725
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__26167\,
            I => n10725
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__26152\,
            I => n10725
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__26135\,
            I => n10725
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__26124\,
            I => n10725
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__26121\,
            I => n10725
        );

    \I__4576\ : Odrv12
    port map (
            O => \N__26118\,
            I => n10725
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__26115\,
            I => n10725
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__26106\,
            I => n10725
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__26095\,
            I => n10725
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__26086\,
            I => n10725
        );

    \I__4571\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26049\
        );

    \I__4570\ : InMux
    port map (
            O => \N__26054\,
            I => \N__26046\
        );

    \I__4569\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26043\
        );

    \I__4568\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26039\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__26049\,
            I => \N__26036\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__26046\,
            I => \N__26033\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__26043\,
            I => \N__26029\
        );

    \I__4564\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26026\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__26039\,
            I => \N__26023\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__26036\,
            I => \N__26017\
        );

    \I__4561\ : Span4Mux_h
    port map (
            O => \N__26033\,
            I => \N__26017\
        );

    \I__4560\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26014\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__26029\,
            I => \N__26011\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__26026\,
            I => \N__26006\
        );

    \I__4557\ : Span4Mux_h
    port map (
            O => \N__26023\,
            I => \N__26006\
        );

    \I__4556\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26003\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__26017\,
            I => \N__26000\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__26014\,
            I => \N__25993\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__26011\,
            I => \N__25993\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__26006\,
            I => \N__25993\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__26003\,
            I => data_out_frame2_12_0
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__26000\,
            I => data_out_frame2_12_0
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__25993\,
            I => data_out_frame2_12_0
        );

    \I__4548\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25978\
        );

    \I__4547\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25978\
        );

    \I__4546\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25975\
        );

    \I__4545\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25972\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__25978\,
            I => \N__25969\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__25975\,
            I => \N__25963\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__25972\,
            I => \N__25963\
        );

    \I__4541\ : Span4Mux_v
    port map (
            O => \N__25969\,
            I => \N__25959\
        );

    \I__4540\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25956\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__25963\,
            I => \N__25953\
        );

    \I__4538\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25950\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__25959\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__25956\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__25953\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__25950\,
            I => \r_SM_Main_2_N_2031_1\
        );

    \I__4533\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25931\
        );

    \I__4532\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25928\
        );

    \I__4531\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25925\
        );

    \I__4530\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25920\
        );

    \I__4529\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25920\
        );

    \I__4528\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25917\
        );

    \I__4527\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25912\
        );

    \I__4526\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25912\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25907\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__25928\,
            I => \N__25907\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__25925\,
            I => \N__25904\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__25920\,
            I => \N__25901\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__25917\,
            I => \N__25898\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25893\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__25907\,
            I => \N__25893\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__25904\,
            I => \r_SM_Main_0\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__25901\,
            I => \r_SM_Main_0\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__25898\,
            I => \r_SM_Main_0\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__25893\,
            I => \r_SM_Main_0\
        );

    \I__4514\ : InMux
    port map (
            O => \N__25884\,
            I => \N__25881\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__25881\,
            I => \N__25878\
        );

    \I__4512\ : Span4Mux_h
    port map (
            O => \N__25878\,
            I => \N__25875\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__25875\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_12\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__25872\,
            I => \N__25869\
        );

    \I__4509\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25863\
        );

    \I__4508\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25858\
        );

    \I__4507\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25858\
        );

    \I__4506\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25855\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__25863\,
            I => \N__25852\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25849\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25846\
        );

    \I__4502\ : Span4Mux_h
    port map (
            O => \N__25852\,
            I => \N__25843\
        );

    \I__4501\ : Span12Mux_v
    port map (
            O => \N__25849\,
            I => \N__25840\
        );

    \I__4500\ : Odrv12
    port map (
            O => \N__25846\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__25843\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__4498\ : Odrv12
    port map (
            O => \N__25840\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__4497\ : SRMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__4495\ : Span4Mux_s2_v
    port map (
            O => \N__25827\,
            I => \N__25824\
        );

    \I__4494\ : Span4Mux_v
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__25821\,
            I => \c0.n3_adj_2268\
        );

    \I__4492\ : InMux
    port map (
            O => \N__25818\,
            I => \bfn_9_17_0_\
        );

    \I__4491\ : InMux
    port map (
            O => \N__25815\,
            I => \c0.n15972\
        );

    \I__4490\ : InMux
    port map (
            O => \N__25812\,
            I => \c0.n15973\
        );

    \I__4489\ : InMux
    port map (
            O => \N__25809\,
            I => \c0.n15974\
        );

    \I__4488\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__25803\,
            I => \c0.n17606\
        );

    \I__4486\ : InMux
    port map (
            O => \N__25800\,
            I => \c0.n15975\
        );

    \I__4485\ : InMux
    port map (
            O => \N__25797\,
            I => \c0.n15976\
        );

    \I__4484\ : CascadeMux
    port map (
            O => \N__25794\,
            I => \N__25788\
        );

    \I__4483\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25785\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__25792\,
            I => \N__25782\
        );

    \I__4481\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25777\
        );

    \I__4480\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25777\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__25785\,
            I => \N__25774\
        );

    \I__4478\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25768\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__25777\,
            I => \N__25765\
        );

    \I__4476\ : Span12Mux_s4_v
    port map (
            O => \N__25774\,
            I => \N__25762\
        );

    \I__4475\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25759\
        );

    \I__4474\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25754\
        );

    \I__4473\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25754\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25749\
        );

    \I__4471\ : Span4Mux_v
    port map (
            O => \N__25765\,
            I => \N__25749\
        );

    \I__4470\ : Odrv12
    port map (
            O => \N__25762\,
            I => \r_Bit_Index_1_adj_2441\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__25759\,
            I => \r_Bit_Index_1_adj_2441\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__25754\,
            I => \r_Bit_Index_1_adj_2441\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__25749\,
            I => \r_Bit_Index_1_adj_2441\
        );

    \I__4466\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__25737\,
            I => \N__25731\
        );

    \I__4464\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25726\
        );

    \I__4463\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25721\
        );

    \I__4462\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25721\
        );

    \I__4461\ : Span12Mux_s6_v
    port map (
            O => \N__25731\,
            I => \N__25718\
        );

    \I__4460\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25713\
        );

    \I__4459\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25713\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__25726\,
            I => \N__25710\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__25721\,
            I => \r_Bit_Index_0_adj_2442\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__25718\,
            I => \r_Bit_Index_0_adj_2442\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__25713\,
            I => \r_Bit_Index_0_adj_2442\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__25710\,
            I => \r_Bit_Index_0_adj_2442\
        );

    \I__4453\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__25698\,
            I => \N__25695\
        );

    \I__4451\ : Span12Mux_v
    port map (
            O => \N__25695\,
            I => \N__25692\
        );

    \I__4450\ : Odrv12
    port map (
            O => \N__25692\,
            I => n5266
        );

    \I__4449\ : IoInMux
    port map (
            O => \N__25689\,
            I => \N__25686\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__4447\ : Span4Mux_s3_v
    port map (
            O => \N__25683\,
            I => \N__25680\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__25680\,
            I => tx_enable
        );

    \I__4445\ : CEMux
    port map (
            O => \N__25677\,
            I => \N__25673\
        );

    \I__4444\ : CEMux
    port map (
            O => \N__25676\,
            I => \N__25669\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25666\
        );

    \I__4442\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25663\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25660\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__25666\,
            I => \N__25655\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__25663\,
            I => \N__25655\
        );

    \I__4438\ : Sp12to4
    port map (
            O => \N__25660\,
            I => \N__25650\
        );

    \I__4437\ : Sp12to4
    port map (
            O => \N__25655\,
            I => \N__25650\
        );

    \I__4436\ : Odrv12
    port map (
            O => \N__25650\,
            I => n10674
        );

    \I__4435\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__25644\,
            I => \N__25641\
        );

    \I__4433\ : Odrv12
    port map (
            O => \N__25641\,
            I => \c0.n17574\
        );

    \I__4432\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25635\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__4430\ : Span4Mux_s2_v
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__25629\,
            I => \c0.rx.n10620\
        );

    \I__4428\ : InMux
    port map (
            O => \N__25626\,
            I => \N__25620\
        );

    \I__4427\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25613\
        );

    \I__4426\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25613\
        );

    \I__4425\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25613\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__25620\,
            I => \N__25608\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__25613\,
            I => \N__25608\
        );

    \I__4422\ : Span4Mux_s2_v
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__25605\,
            I => n17361
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__4419\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25595\
        );

    \I__4418\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25592\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__25595\,
            I => \N__25588\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25585\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__25591\,
            I => \N__25581\
        );

    \I__4414\ : Span4Mux_s2_v
    port map (
            O => \N__25588\,
            I => \N__25578\
        );

    \I__4413\ : Span4Mux_s2_v
    port map (
            O => \N__25585\,
            I => \N__25575\
        );

    \I__4412\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25570\
        );

    \I__4411\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25570\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__25578\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__25575\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__25570\,
            I => \c0.rx.r_SM_Main_2_N_2088_2\
        );

    \I__4407\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25553\
        );

    \I__4406\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25553\
        );

    \I__4405\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25553\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__25560\,
            I => \N__25547\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__25553\,
            I => \N__25541\
        );

    \I__4402\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25534\
        );

    \I__4401\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25534\
        );

    \I__4400\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25534\
        );

    \I__4399\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25531\
        );

    \I__4398\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25524\
        );

    \I__4397\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25524\
        );

    \I__4396\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25524\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__25541\,
            I => \N__25521\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__25534\,
            I => \r_SM_Main_1\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__25531\,
            I => \r_SM_Main_1\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__25524\,
            I => \r_SM_Main_1\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__25521\,
            I => \r_SM_Main_1\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__25512\,
            I => \c0.rx.r_SM_Main_2_N_2088_2_cascade_\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__25509\,
            I => \N__25504\
        );

    \I__4388\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25499\
        );

    \I__4387\ : InMux
    port map (
            O => \N__25507\,
            I => \N__25496\
        );

    \I__4386\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25489\
        );

    \I__4385\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25489\
        );

    \I__4384\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25489\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__25499\,
            I => \N__25479\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__25496\,
            I => \N__25479\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__25489\,
            I => \N__25476\
        );

    \I__4380\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25469\
        );

    \I__4379\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25469\
        );

    \I__4378\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25469\
        );

    \I__4377\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25464\
        );

    \I__4376\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25464\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__25479\,
            I => \N__25461\
        );

    \I__4374\ : Span4Mux_h
    port map (
            O => \N__25476\,
            I => \N__25458\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__25469\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__25464\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__25461\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__25458\,
            I => \c0.rx.r_SM_Main_0\
        );

    \I__4369\ : SRMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__25440\,
            I => \c0.n3_adj_2254\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__25437\,
            I => \N__25434\
        );

    \I__4364\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25426\
        );

    \I__4363\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25426\
        );

    \I__4362\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25423\
        );

    \I__4361\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25420\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__25426\,
            I => \N__25417\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__25423\,
            I => \N__25414\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__25420\,
            I => \N__25411\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__25417\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__4356\ : Odrv12
    port map (
            O => \N__25414\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__25411\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__4354\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__25395\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_18\
        );

    \I__4350\ : SRMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__25389\,
            I => \N__25386\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__25380\,
            I => \c0.n3_adj_2288\
        );

    \I__4345\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__4343\ : Span4Mux_h
    port map (
            O => \N__25371\,
            I => \N__25368\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__25368\,
            I => \N__25365\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__25365\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_1\
        );

    \I__4340\ : SRMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__25353\,
            I => \N__25350\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__25350\,
            I => \c0.n3_adj_2246\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__4334\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25337\
        );

    \I__4333\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25337\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__25342\,
            I => \N__25334\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__25337\,
            I => \N__25331\
        );

    \I__4330\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25328\
        );

    \I__4329\ : Span4Mux_v
    port map (
            O => \N__25331\,
            I => \N__25322\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__25328\,
            I => \N__25322\
        );

    \I__4327\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25319\
        );

    \I__4326\ : Span4Mux_h
    port map (
            O => \N__25322\,
            I => \N__25316\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__25319\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__25316\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__4323\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25308\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__25308\,
            I => \N__25305\
        );

    \I__4321\ : Span4Mux_v
    port map (
            O => \N__25305\,
            I => \N__25302\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__25302\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_22\
        );

    \I__4319\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25295\
        );

    \I__4318\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25292\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__25295\,
            I => \N__25289\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__25292\,
            I => \N__25285\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__25289\,
            I => \N__25282\
        );

    \I__4314\ : InMux
    port map (
            O => \N__25288\,
            I => \N__25278\
        );

    \I__4313\ : Span4Mux_h
    port map (
            O => \N__25285\,
            I => \N__25275\
        );

    \I__4312\ : Span4Mux_v
    port map (
            O => \N__25282\,
            I => \N__25272\
        );

    \I__4311\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25269\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__25278\,
            I => \N__25266\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__25275\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__25272\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__25269\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__4306\ : Odrv12
    port map (
            O => \N__25266\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__4305\ : SRMux
    port map (
            O => \N__25257\,
            I => \N__25254\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__25254\,
            I => \N__25251\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__4302\ : Span4Mux_v
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__25245\,
            I => \c0.n3_adj_2238\
        );

    \I__4300\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__25236\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_10\
        );

    \I__4297\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25230\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__25230\,
            I => \N__25227\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__25224\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_26\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__25221\,
            I => \N__25215\
        );

    \I__4292\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25212\
        );

    \I__4291\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25207\
        );

    \I__4290\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25207\
        );

    \I__4289\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25204\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25201\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25198\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__25204\,
            I => \N__25195\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__25201\,
            I => \N__25192\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__25198\,
            I => \N__25189\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__25195\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__25192\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__25189\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__4280\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__25179\,
            I => \N__25176\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__25176\,
            I => \N__25173\
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__25173\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_25\
        );

    \I__4276\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25166\
        );

    \I__4275\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25163\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25160\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__25163\,
            I => \N__25155\
        );

    \I__4272\ : Span4Mux_h
    port map (
            O => \N__25160\,
            I => \N__25152\
        );

    \I__4271\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25147\
        );

    \I__4270\ : InMux
    port map (
            O => \N__25158\,
            I => \N__25147\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__25155\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__25152\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__25147\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__4266\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25137\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__25134\,
            I => \N__25131\
        );

    \I__4263\ : Span4Mux_s3_h
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__25128\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_24\
        );

    \I__4261\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25121\
        );

    \I__4260\ : CascadeMux
    port map (
            O => \N__25124\,
            I => \N__25116\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__25121\,
            I => \N__25113\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__25120\,
            I => \N__25110\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__25119\,
            I => \N__25107\
        );

    \I__4256\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25104\
        );

    \I__4255\ : Span4Mux_v
    port map (
            O => \N__25113\,
            I => \N__25101\
        );

    \I__4254\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25096\
        );

    \I__4253\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25096\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__25104\,
            I => \N__25093\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__25101\,
            I => \N__25090\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__25096\,
            I => \N__25087\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__25093\,
            I => \N__25082\
        );

    \I__4248\ : Span4Mux_h
    port map (
            O => \N__25090\,
            I => \N__25082\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__25087\,
            I => \N__25079\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__25082\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__25079\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__4244\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__4242\ : Span4Mux_h
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__25065\,
            I => \N__25062\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__25062\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_23\
        );

    \I__4239\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25050\
        );

    \I__4237\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25045\
        );

    \I__4236\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25045\
        );

    \I__4235\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25042\
        );

    \I__4234\ : Span4Mux_v
    port map (
            O => \N__25050\,
            I => \N__25039\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__25045\,
            I => \N__25036\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__25042\,
            I => \N__25033\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__25039\,
            I => \N__25030\
        );

    \I__4230\ : Span4Mux_h
    port map (
            O => \N__25036\,
            I => \N__25027\
        );

    \I__4229\ : Odrv12
    port map (
            O => \N__25033\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__25030\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__25027\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__4226\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__4224\ : Span4Mux_h
    port map (
            O => \N__25014\,
            I => \N__25011\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__25011\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_20\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__25008\,
            I => \N__25004\
        );

    \I__4221\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25001\
        );

    \I__4220\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24998\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__25001\,
            I => \N__24995\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__24998\,
            I => \N__24990\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__24995\,
            I => \N__24987\
        );

    \I__4216\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24982\
        );

    \I__4215\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24982\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__24990\,
            I => \N__24979\
        );

    \I__4213\ : Sp12to4
    port map (
            O => \N__24987\,
            I => \N__24974\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__24982\,
            I => \N__24974\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__24979\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__4210\ : Odrv12
    port map (
            O => \N__24974\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__4209\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__4207\ : Span4Mux_h
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__4206\ : Span4Mux_h
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__24957\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_19\
        );

    \I__4204\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24951\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__4202\ : Span12Mux_s6_v
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__4201\ : Odrv12
    port map (
            O => \N__24945\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_16\
        );

    \I__4200\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24938\
        );

    \I__4199\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24933\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__24938\,
            I => \N__24930\
        );

    \I__4197\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24927\
        );

    \I__4196\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24924\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__24933\,
            I => \N__24921\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__24930\,
            I => \N__24916\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24916\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24912\
        );

    \I__4191\ : Span4Mux_h
    port map (
            O => \N__24921\,
            I => \N__24909\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__24916\,
            I => \N__24906\
        );

    \I__4189\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24901\
        );

    \I__4188\ : Span4Mux_h
    port map (
            O => \N__24912\,
            I => \N__24896\
        );

    \I__4187\ : Span4Mux_v
    port map (
            O => \N__24909\,
            I => \N__24896\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__24906\,
            I => \N__24893\
        );

    \I__4185\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24888\
        );

    \I__4184\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24888\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__24901\,
            I => data_out_frame2_16_0
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__24896\,
            I => data_out_frame2_16_0
        );

    \I__4181\ : Odrv4
    port map (
            O => \N__24893\,
            I => data_out_frame2_16_0
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__24888\,
            I => data_out_frame2_16_0
        );

    \I__4179\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__24870\,
            I => \N__24866\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__24869\,
            I => \N__24863\
        );

    \I__4174\ : Span4Mux_v
    port map (
            O => \N__24866\,
            I => \N__24860\
        );

    \I__4173\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24857\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__24860\,
            I => \c0.n17098\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__24857\,
            I => \c0.n17098\
        );

    \I__4170\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24847\
        );

    \I__4169\ : InMux
    port map (
            O => \N__24851\,
            I => \N__24842\
        );

    \I__4168\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24839\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24836\
        );

    \I__4166\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24833\
        );

    \I__4165\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24829\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__24842\,
            I => \N__24826\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24823\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__24836\,
            I => \N__24818\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24818\
        );

    \I__4160\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24815\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24812\
        );

    \I__4158\ : Span4Mux_h
    port map (
            O => \N__24826\,
            I => \N__24805\
        );

    \I__4157\ : Span4Mux_h
    port map (
            O => \N__24823\,
            I => \N__24805\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__24818\,
            I => \N__24805\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__24815\,
            I => data_out_frame2_8_3
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__24812\,
            I => data_out_frame2_8_3
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__24805\,
            I => data_out_frame2_8_3
        );

    \I__4152\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24795\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__4150\ : Span4Mux_h
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__24789\,
            I => \c0.n17_adj_2321\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__24786\,
            I => \c0.n30_cascade_\
        );

    \I__4147\ : InMux
    port map (
            O => \N__24783\,
            I => \N__24779\
        );

    \I__4146\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24775\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24771\
        );

    \I__4144\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24768\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__24775\,
            I => \N__24765\
        );

    \I__4142\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24762\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__24771\,
            I => \N__24759\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__24768\,
            I => data_out_frame2_14_4
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__24765\,
            I => data_out_frame2_14_4
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__24762\,
            I => data_out_frame2_14_4
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__24759\,
            I => data_out_frame2_14_4
        );

    \I__4136\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24745\
        );

    \I__4135\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24740\
        );

    \I__4134\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24737\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__24745\,
            I => \N__24734\
        );

    \I__4132\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24731\
        );

    \I__4131\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24728\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__24740\,
            I => \N__24725\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__24737\,
            I => \N__24722\
        );

    \I__4128\ : Span4Mux_v
    port map (
            O => \N__24734\,
            I => \N__24719\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24716\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__24728\,
            I => data_out_frame2_11_0
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__24725\,
            I => data_out_frame2_11_0
        );

    \I__4124\ : Odrv12
    port map (
            O => \N__24722\,
            I => data_out_frame2_11_0
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__24719\,
            I => data_out_frame2_11_0
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__24716\,
            I => data_out_frame2_11_0
        );

    \I__4121\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__4119\ : Span4Mux_v
    port map (
            O => \N__24699\,
            I => \N__24695\
        );

    \I__4118\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24692\
        );

    \I__4117\ : IoSpan4Mux
    port map (
            O => \N__24695\,
            I => \N__24689\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__24692\,
            I => \N__24686\
        );

    \I__4115\ : Span4Mux_s2_h
    port map (
            O => \N__24689\,
            I => \N__24681\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__24686\,
            I => \N__24681\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__24681\,
            I => \N__24678\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__24678\,
            I => \c0.n17276\
        );

    \I__4111\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24669\
        );

    \I__4110\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24662\
        );

    \I__4109\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24662\
        );

    \I__4108\ : InMux
    port map (
            O => \N__24672\,
            I => \N__24662\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24657\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__24662\,
            I => \N__24657\
        );

    \I__4105\ : Odrv12
    port map (
            O => \N__24657\,
            I => n17412
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__24654\,
            I => \N__24648\
        );

    \I__4103\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24643\
        );

    \I__4102\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24643\
        );

    \I__4101\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24640\
        );

    \I__4100\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24637\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__24643\,
            I => \N__24633\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24630\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__24637\,
            I => \N__24627\
        );

    \I__4096\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24624\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__24633\,
            I => \N__24621\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__24630\,
            I => \N__24616\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__24627\,
            I => \N__24616\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__24624\,
            I => data_out_frame2_9_3
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__24621\,
            I => data_out_frame2_9_3
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__24616\,
            I => data_out_frame2_9_3
        );

    \I__4089\ : InMux
    port map (
            O => \N__24609\,
            I => \N__24606\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__24606\,
            I => \N__24603\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__24603\,
            I => \N__24600\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__24600\,
            I => \c0.n6_adj_2197\
        );

    \I__4085\ : InMux
    port map (
            O => \N__24597\,
            I => \N__24593\
        );

    \I__4084\ : InMux
    port map (
            O => \N__24596\,
            I => \N__24590\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__24593\,
            I => \N__24587\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__24590\,
            I => \N__24584\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__24587\,
            I => \N__24579\
        );

    \I__4080\ : Span4Mux_v
    port map (
            O => \N__24584\,
            I => \N__24576\
        );

    \I__4079\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24573\
        );

    \I__4078\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24570\
        );

    \I__4077\ : Span4Mux_h
    port map (
            O => \N__24579\,
            I => \N__24567\
        );

    \I__4076\ : Span4Mux_h
    port map (
            O => \N__24576\,
            I => \N__24562\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__24573\,
            I => \N__24562\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__24570\,
            I => data_out_frame2_15_7
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__24567\,
            I => data_out_frame2_15_7
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__24562\,
            I => data_out_frame2_15_7
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__4070\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24548\
        );

    \I__4069\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24545\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__24548\,
            I => \N__24542\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__24545\,
            I => \N__24539\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__24542\,
            I => \N__24536\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__24539\,
            I => \N__24533\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__24536\,
            I => \c0.n17123\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__24533\,
            I => \c0.n17123\
        );

    \I__4062\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24522\
        );

    \I__4061\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24519\
        );

    \I__4060\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24516\
        );

    \I__4059\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24513\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__24522\,
            I => \N__24510\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__24519\,
            I => \N__24507\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__24516\,
            I => data_out_frame2_14_6
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__24513\,
            I => data_out_frame2_14_6
        );

    \I__4054\ : Odrv12
    port map (
            O => \N__24510\,
            I => data_out_frame2_14_6
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__24507\,
            I => data_out_frame2_14_6
        );

    \I__4052\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__4050\ : Span4Mux_v
    port map (
            O => \N__24492\,
            I => \N__24489\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__24489\,
            I => \N__24486\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__24486\,
            I => \c0.n10434\
        );

    \I__4047\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24478\
        );

    \I__4046\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24475\
        );

    \I__4045\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24472\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24468\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__24475\,
            I => \N__24465\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__24472\,
            I => \N__24461\
        );

    \I__4041\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24458\
        );

    \I__4040\ : Span4Mux_v
    port map (
            O => \N__24468\,
            I => \N__24453\
        );

    \I__4039\ : Span4Mux_s3_h
    port map (
            O => \N__24465\,
            I => \N__24453\
        );

    \I__4038\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24450\
        );

    \I__4037\ : Span4Mux_h
    port map (
            O => \N__24461\,
            I => \N__24447\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__24458\,
            I => \N__24442\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__24453\,
            I => \N__24442\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__24450\,
            I => data_out_frame2_16_3
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__24447\,
            I => data_out_frame2_16_3
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__24442\,
            I => data_out_frame2_16_3
        );

    \I__4031\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24430\
        );

    \I__4030\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24427\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__24433\,
            I => \N__24423\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24419\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24416\
        );

    \I__4026\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24411\
        );

    \I__4025\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24411\
        );

    \I__4024\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24408\
        );

    \I__4023\ : Span4Mux_v
    port map (
            O => \N__24419\,
            I => \N__24401\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__24416\,
            I => \N__24401\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24401\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__24408\,
            I => data_out_frame2_15_3
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__24401\,
            I => data_out_frame2_15_3
        );

    \I__4018\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__4016\ : Span4Mux_s3_h
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__24384\,
            I => \c0.n10482\
        );

    \I__4013\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24377\
        );

    \I__4012\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__24377\,
            I => \N__24371\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24368\
        );

    \I__4009\ : Span4Mux_s3_h
    port map (
            O => \N__24371\,
            I => \N__24362\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__24368\,
            I => \N__24362\
        );

    \I__4007\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24359\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__24362\,
            I => \N__24354\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24351\
        );

    \I__4004\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24347\
        );

    \I__4003\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24344\
        );

    \I__4002\ : Span4Mux_s3_h
    port map (
            O => \N__24354\,
            I => \N__24339\
        );

    \I__4001\ : Span4Mux_v
    port map (
            O => \N__24351\,
            I => \N__24339\
        );

    \I__4000\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24336\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__24347\,
            I => data_out_frame2_8_4
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__24344\,
            I => data_out_frame2_8_4
        );

    \I__3997\ : Odrv4
    port map (
            O => \N__24339\,
            I => data_out_frame2_8_4
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__24336\,
            I => data_out_frame2_8_4
        );

    \I__3995\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24324\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__24324\,
            I => \N__24320\
        );

    \I__3993\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24317\
        );

    \I__3992\ : Span4Mux_s2_h
    port map (
            O => \N__24320\,
            I => \N__24312\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__24317\,
            I => \N__24309\
        );

    \I__3990\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24305\
        );

    \I__3989\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24302\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__24312\,
            I => \N__24299\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__24309\,
            I => \N__24296\
        );

    \I__3986\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24293\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__24305\,
            I => data_out_frame2_8_0
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__24302\,
            I => data_out_frame2_8_0
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__24299\,
            I => data_out_frame2_8_0
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__24296\,
            I => data_out_frame2_8_0
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__24293\,
            I => data_out_frame2_8_0
        );

    \I__3980\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24279\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__3978\ : Odrv12
    port map (
            O => \N__24276\,
            I => \c0.n10513\
        );

    \I__3977\ : CEMux
    port map (
            O => \N__24273\,
            I => \N__24266\
        );

    \I__3976\ : CEMux
    port map (
            O => \N__24272\,
            I => \N__24261\
        );

    \I__3975\ : CEMux
    port map (
            O => \N__24271\,
            I => \N__24258\
        );

    \I__3974\ : CEMux
    port map (
            O => \N__24270\,
            I => \N__24255\
        );

    \I__3973\ : CEMux
    port map (
            O => \N__24269\,
            I => \N__24251\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__24266\,
            I => \N__24248\
        );

    \I__3971\ : CEMux
    port map (
            O => \N__24265\,
            I => \N__24245\
        );

    \I__3970\ : CEMux
    port map (
            O => \N__24264\,
            I => \N__24242\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__24261\,
            I => \N__24239\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24236\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24233\
        );

    \I__3966\ : CEMux
    port map (
            O => \N__24254\,
            I => \N__24230\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24227\
        );

    \I__3964\ : Span4Mux_v
    port map (
            O => \N__24248\,
            I => \N__24224\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24221\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__24242\,
            I => \N__24218\
        );

    \I__3961\ : Span4Mux_s3_h
    port map (
            O => \N__24239\,
            I => \N__24209\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__24236\,
            I => \N__24209\
        );

    \I__3959\ : Span4Mux_s3_h
    port map (
            O => \N__24233\,
            I => \N__24209\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24209\
        );

    \I__3957\ : Sp12to4
    port map (
            O => \N__24227\,
            I => \N__24206\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__24224\,
            I => \N__24201\
        );

    \I__3955\ : Span4Mux_v
    port map (
            O => \N__24221\,
            I => \N__24201\
        );

    \I__3954\ : Span4Mux_v
    port map (
            O => \N__24218\,
            I => \N__24198\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__24209\,
            I => \N__24195\
        );

    \I__3952\ : Span12Mux_v
    port map (
            O => \N__24206\,
            I => \N__24192\
        );

    \I__3951\ : Sp12to4
    port map (
            O => \N__24201\,
            I => \N__24189\
        );

    \I__3950\ : Span4Mux_h
    port map (
            O => \N__24198\,
            I => \N__24184\
        );

    \I__3949\ : Span4Mux_h
    port map (
            O => \N__24195\,
            I => \N__24184\
        );

    \I__3948\ : Odrv12
    port map (
            O => \N__24192\,
            I => \c0.tx2.n9269\
        );

    \I__3947\ : Odrv12
    port map (
            O => \N__24189\,
            I => \c0.tx2.n9269\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__24184\,
            I => \c0.tx2.n9269\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__24177\,
            I => \N__24173\
        );

    \I__3944\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24170\
        );

    \I__3943\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24167\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24164\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__24167\,
            I => \N__24160\
        );

    \I__3940\ : Span4Mux_h
    port map (
            O => \N__24164\,
            I => \N__24157\
        );

    \I__3939\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24153\
        );

    \I__3938\ : Span4Mux_v
    port map (
            O => \N__24160\,
            I => \N__24148\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__24157\,
            I => \N__24148\
        );

    \I__3936\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24145\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__24153\,
            I => data_out_frame2_5_2
        );

    \I__3934\ : Odrv4
    port map (
            O => \N__24148\,
            I => data_out_frame2_5_2
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__24145\,
            I => data_out_frame2_5_2
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__24138\,
            I => \N__24134\
        );

    \I__3931\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24130\
        );

    \I__3930\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24126\
        );

    \I__3929\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24123\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24120\
        );

    \I__3927\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24117\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__24126\,
            I => \N__24114\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__24123\,
            I => data_out_frame2_10_4
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__24120\,
            I => data_out_frame2_10_4
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__24117\,
            I => data_out_frame2_10_4
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__24114\,
            I => data_out_frame2_10_4
        );

    \I__3921\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24102\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24099\
        );

    \I__3919\ : Span4Mux_s2_h
    port map (
            O => \N__24099\,
            I => \N__24095\
        );

    \I__3918\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24092\
        );

    \I__3917\ : Span4Mux_h
    port map (
            O => \N__24095\,
            I => \N__24089\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__24092\,
            I => \N__24086\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__24089\,
            I => \c0.n10456\
        );

    \I__3914\ : Odrv12
    port map (
            O => \N__24086\,
            I => \c0.n10456\
        );

    \I__3913\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24074\
        );

    \I__3912\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24074\
        );

    \I__3911\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24070\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24067\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__24073\,
            I => \N__24064\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24060\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__24067\,
            I => \N__24057\
        );

    \I__3906\ : InMux
    port map (
            O => \N__24064\,
            I => \N__24054\
        );

    \I__3905\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24051\
        );

    \I__3904\ : Span4Mux_h
    port map (
            O => \N__24060\,
            I => \N__24048\
        );

    \I__3903\ : Sp12to4
    port map (
            O => \N__24057\,
            I => \N__24043\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24043\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__24051\,
            I => data_out_frame2_10_5
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__24048\,
            I => data_out_frame2_10_5
        );

    \I__3899\ : Odrv12
    port map (
            O => \N__24043\,
            I => data_out_frame2_10_5
        );

    \I__3898\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24033\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__24033\,
            I => \N__24028\
        );

    \I__3896\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24025\
        );

    \I__3895\ : InMux
    port map (
            O => \N__24031\,
            I => \N__24021\
        );

    \I__3894\ : Span4Mux_h
    port map (
            O => \N__24028\,
            I => \N__24018\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24015\
        );

    \I__3892\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24012\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__24021\,
            I => data_out_frame2_11_3
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__24018\,
            I => data_out_frame2_11_3
        );

    \I__3889\ : Odrv12
    port map (
            O => \N__24015\,
            I => data_out_frame2_11_3
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__24012\,
            I => data_out_frame2_11_3
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__3886\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23996\
        );

    \I__3885\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23993\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23989\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__23993\,
            I => \N__23986\
        );

    \I__3882\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23982\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__23989\,
            I => \N__23979\
        );

    \I__3880\ : Span4Mux_h
    port map (
            O => \N__23986\,
            I => \N__23976\
        );

    \I__3879\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23973\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__23982\,
            I => data_out_frame2_14_1
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__23979\,
            I => data_out_frame2_14_1
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__23976\,
            I => data_out_frame2_14_1
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__23973\,
            I => data_out_frame2_14_1
        );

    \I__3874\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__23961\,
            I => \N__23955\
        );

    \I__3872\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23952\
        );

    \I__3871\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23949\
        );

    \I__3870\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23946\
        );

    \I__3869\ : Span4Mux_h
    port map (
            O => \N__23955\,
            I => \N__23943\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23940\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__23949\,
            I => data_out_frame2_15_1
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__23946\,
            I => data_out_frame2_15_1
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__23943\,
            I => data_out_frame2_15_1
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__23940\,
            I => data_out_frame2_15_1
        );

    \I__3863\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23928\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__23925\,
            I => \c0.n18016\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__23922\,
            I => \N__23919\
        );

    \I__3859\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23911\
        );

    \I__3858\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23911\
        );

    \I__3857\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23907\
        );

    \I__3856\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23904\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__23911\,
            I => \N__23899\
        );

    \I__3854\ : InMux
    port map (
            O => \N__23910\,
            I => \N__23896\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__23907\,
            I => \N__23893\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23890\
        );

    \I__3851\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23887\
        );

    \I__3850\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23884\
        );

    \I__3849\ : Span4Mux_v
    port map (
            O => \N__23899\,
            I => \N__23881\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__23896\,
            I => \N__23878\
        );

    \I__3847\ : Span4Mux_s3_h
    port map (
            O => \N__23893\,
            I => \N__23873\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__23890\,
            I => \N__23873\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23870\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__23884\,
            I => data_out_frame2_12_2
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__23881\,
            I => data_out_frame2_12_2
        );

    \I__3842\ : Odrv12
    port map (
            O => \N__23878\,
            I => data_out_frame2_12_2
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__23873\,
            I => data_out_frame2_12_2
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__23870\,
            I => data_out_frame2_12_2
        );

    \I__3839\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__23856\,
            I => \N__23853\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__23853\,
            I => \N__23848\
        );

    \I__3836\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23845\
        );

    \I__3835\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23841\
        );

    \I__3834\ : Span4Mux_h
    port map (
            O => \N__23848\,
            I => \N__23836\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__23845\,
            I => \N__23836\
        );

    \I__3832\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23833\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__23841\,
            I => \N__23830\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__23836\,
            I => \N__23827\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__23833\,
            I => data_out_frame2_7_2
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__23830\,
            I => data_out_frame2_7_2
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__23827\,
            I => data_out_frame2_7_2
        );

    \I__3826\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23816\
        );

    \I__3825\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23811\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23808\
        );

    \I__3823\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23805\
        );

    \I__3822\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23802\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__23811\,
            I => \N__23799\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__23808\,
            I => \N__23794\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__23805\,
            I => \N__23794\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__23802\,
            I => data_out_frame2_6_2
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__23799\,
            I => data_out_frame2_6_2
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__23794\,
            I => data_out_frame2_6_2
        );

    \I__3815\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__23781\,
            I => \N__23778\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__23778\,
            I => \N__23775\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__23775\,
            I => \c0.n5_adj_2290\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__23772\,
            I => \N__23768\
        );

    \I__3809\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23763\
        );

    \I__3808\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23763\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__23763\,
            I => \N__23759\
        );

    \I__3806\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23756\
        );

    \I__3805\ : Span4Mux_h
    port map (
            O => \N__23759\,
            I => \N__23751\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23751\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__23751\,
            I => \c0.n10563\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__23748\,
            I => \N__23745\
        );

    \I__3801\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23741\
        );

    \I__3800\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23738\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__23741\,
            I => \N__23735\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23732\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__23735\,
            I => \N__23729\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__23732\,
            I => \N__23726\
        );

    \I__3795\ : Span4Mux_h
    port map (
            O => \N__23729\,
            I => \N__23718\
        );

    \I__3794\ : Span4Mux_v
    port map (
            O => \N__23726\,
            I => \N__23718\
        );

    \I__3793\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23715\
        );

    \I__3792\ : InMux
    port map (
            O => \N__23724\,
            I => \N__23712\
        );

    \I__3791\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23709\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__23718\,
            I => \N__23706\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23703\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__23712\,
            I => data_out_frame2_13_5
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__23709\,
            I => data_out_frame2_13_5
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__23706\,
            I => data_out_frame2_13_5
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__23703\,
            I => data_out_frame2_13_5
        );

    \I__3784\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__23688\,
            I => \N__23684\
        );

    \I__3781\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23681\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__23684\,
            I => \c0.n17095\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__23681\,
            I => \c0.n17095\
        );

    \I__3778\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__3776\ : Odrv12
    port map (
            O => \N__23670\,
            I => \c0.n31\
        );

    \I__3775\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23663\
        );

    \I__3774\ : InMux
    port map (
            O => \N__23666\,
            I => \N__23660\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23655\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23655\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__23655\,
            I => \N__23649\
        );

    \I__3770\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23646\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__23653\,
            I => \N__23643\
        );

    \I__3768\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23640\
        );

    \I__3767\ : Span4Mux_s3_h
    port map (
            O => \N__23649\,
            I => \N__23637\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23634\
        );

    \I__3765\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23631\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__23640\,
            I => data_out_frame2_13_1
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__23637\,
            I => data_out_frame2_13_1
        );

    \I__3762\ : Odrv12
    port map (
            O => \N__23634\,
            I => data_out_frame2_13_1
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__23631\,
            I => data_out_frame2_13_1
        );

    \I__3760\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23618\
        );

    \I__3759\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23615\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23609\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23606\
        );

    \I__3756\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23603\
        );

    \I__3755\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23599\
        );

    \I__3754\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23596\
        );

    \I__3753\ : Span4Mux_v
    port map (
            O => \N__23609\,
            I => \N__23589\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__23606\,
            I => \N__23589\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23589\
        );

    \I__3750\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23586\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__23599\,
            I => data_out_frame2_12_1
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__23596\,
            I => data_out_frame2_12_1
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__23589\,
            I => data_out_frame2_12_1
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__23586\,
            I => data_out_frame2_12_1
        );

    \I__3745\ : InMux
    port map (
            O => \N__23577\,
            I => \N__23574\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__23574\,
            I => \N__23571\
        );

    \I__3743\ : Span4Mux_v
    port map (
            O => \N__23571\,
            I => \N__23568\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__23568\,
            I => \c0.n18019\
        );

    \I__3741\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23558\
        );

    \I__3740\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23558\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__23563\,
            I => \N__23555\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23551\
        );

    \I__3737\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23548\
        );

    \I__3736\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23543\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__23551\,
            I => \N__23540\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__23548\,
            I => \N__23537\
        );

    \I__3733\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23532\
        );

    \I__3732\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23532\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__23543\,
            I => data_out_frame2_12_3
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__23540\,
            I => data_out_frame2_12_3
        );

    \I__3729\ : Odrv12
    port map (
            O => \N__23537\,
            I => data_out_frame2_12_3
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__23532\,
            I => data_out_frame2_12_3
        );

    \I__3727\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23519\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__23522\,
            I => \N__23516\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__23519\,
            I => \N__23513\
        );

    \I__3724\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23510\
        );

    \I__3723\ : Span4Mux_v
    port map (
            O => \N__23513\,
            I => \N__23505\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__23510\,
            I => \N__23505\
        );

    \I__3721\ : Span4Mux_h
    port map (
            O => \N__23505\,
            I => \N__23500\
        );

    \I__3720\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23495\
        );

    \I__3719\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23495\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__23500\,
            I => data_out_frame2_5_3
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__23495\,
            I => data_out_frame2_5_3
        );

    \I__3716\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23487\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__23487\,
            I => \c0.n18142\
        );

    \I__3714\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23479\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__23483\,
            I => \N__23476\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__23482\,
            I => \N__23472\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23469\
        );

    \I__3710\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23462\
        );

    \I__3709\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23462\
        );

    \I__3708\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23462\
        );

    \I__3707\ : Span4Mux_h
    port map (
            O => \N__23469\,
            I => \N__23459\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__23462\,
            I => data_out_frame2_8_7
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__23459\,
            I => data_out_frame2_8_7
        );

    \I__3704\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23450\
        );

    \I__3703\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23444\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23441\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__23449\,
            I => \N__23438\
        );

    \I__3700\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23435\
        );

    \I__3699\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23432\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23429\
        );

    \I__3697\ : Span12Mux_v
    port map (
            O => \N__23441\,
            I => \N__23426\
        );

    \I__3696\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23423\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__23435\,
            I => data_out_frame2_9_7
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__23432\,
            I => data_out_frame2_9_7
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__23429\,
            I => data_out_frame2_9_7
        );

    \I__3692\ : Odrv12
    port map (
            O => \N__23426\,
            I => data_out_frame2_9_7
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__23423\,
            I => data_out_frame2_9_7
        );

    \I__3690\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23409\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23406\
        );

    \I__3688\ : Span4Mux_s2_h
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__23400\,
            I => \c0.n18145\
        );

    \I__3685\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23393\
        );

    \I__3684\ : InMux
    port map (
            O => \N__23396\,
            I => \N__23390\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23385\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23382\
        );

    \I__3681\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23378\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__23388\,
            I => \N__23375\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__23385\,
            I => \N__23370\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__23382\,
            I => \N__23370\
        );

    \I__3677\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23367\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23364\
        );

    \I__3675\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23361\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__23370\,
            I => \N__23358\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__23367\,
            I => data_out_frame2_5_1
        );

    \I__3672\ : Odrv12
    port map (
            O => \N__23364\,
            I => data_out_frame2_5_1
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__23361\,
            I => data_out_frame2_5_1
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__23358\,
            I => data_out_frame2_5_1
        );

    \I__3669\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23346\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__3667\ : Span12Mux_v
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__3666\ : Odrv12
    port map (
            O => \N__23340\,
            I => \c0.n6_adj_2142\
        );

    \I__3665\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23334\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__23334\,
            I => \N__23331\
        );

    \I__3663\ : Span4Mux_h
    port map (
            O => \N__23331\,
            I => \N__23328\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__23328\,
            I => \N__23325\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__23325\,
            I => \c0.n18064\
        );

    \I__3660\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23319\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__23319\,
            I => \c0.n18067\
        );

    \I__3658\ : InMux
    port map (
            O => \N__23316\,
            I => \N__23313\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__23310\,
            I => n8191
        );

    \I__3655\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__23304\,
            I => \N__23300\
        );

    \I__3653\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23297\
        );

    \I__3652\ : Span4Mux_h
    port map (
            O => \N__23300\,
            I => \N__23292\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__23297\,
            I => \N__23289\
        );

    \I__3650\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23286\
        );

    \I__3649\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23283\
        );

    \I__3648\ : Span4Mux_v
    port map (
            O => \N__23292\,
            I => \N__23280\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__23289\,
            I => \N__23275\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23275\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__23283\,
            I => data_out_frame2_6_1
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__23280\,
            I => data_out_frame2_6_1
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__23275\,
            I => data_out_frame2_6_1
        );

    \I__3642\ : InMux
    port map (
            O => \N__23268\,
            I => \N__23265\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__23265\,
            I => \c0.n5_adj_2289\
        );

    \I__3640\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23256\
        );

    \I__3639\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23250\
        );

    \I__3638\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23250\
        );

    \I__3637\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23247\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23244\
        );

    \I__3635\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23241\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23234\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__23247\,
            I => \N__23234\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__23244\,
            I => \N__23229\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__23241\,
            I => \N__23229\
        );

    \I__3630\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23226\
        );

    \I__3629\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23223\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__23234\,
            I => \N__23218\
        );

    \I__3627\ : Span4Mux_h
    port map (
            O => \N__23229\,
            I => \N__23218\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__23226\,
            I => data_out_frame2_11_7
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__23223\,
            I => data_out_frame2_11_7
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__23218\,
            I => data_out_frame2_11_7
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__23211\,
            I => \c0.n10413_cascade_\
        );

    \I__3622\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23202\
        );

    \I__3621\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23202\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__3619\ : Span4Mux_s2_h
    port map (
            O => \N__23199\,
            I => \N__23196\
        );

    \I__3618\ : Span4Mux_h
    port map (
            O => \N__23196\,
            I => \N__23193\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__23193\,
            I => \c0.n17282\
        );

    \I__3616\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23187\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__23187\,
            I => \N__23181\
        );

    \I__3614\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23177\
        );

    \I__3613\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23174\
        );

    \I__3612\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23171\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__23181\,
            I => \N__23168\
        );

    \I__3610\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23165\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23160\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23160\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__23171\,
            I => data_out_frame2_10_6
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__23168\,
            I => data_out_frame2_10_6
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__23165\,
            I => data_out_frame2_10_6
        );

    \I__3604\ : Odrv12
    port map (
            O => \N__23160\,
            I => data_out_frame2_10_6
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__23151\,
            I => \N__23147\
        );

    \I__3602\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23144\
        );

    \I__3601\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23141\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23138\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23131\
        );

    \I__3598\ : Span4Mux_v
    port map (
            O => \N__23138\,
            I => \N__23131\
        );

    \I__3597\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23128\
        );

    \I__3596\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23125\
        );

    \I__3595\ : Sp12to4
    port map (
            O => \N__23131\,
            I => \N__23120\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23115\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__23125\,
            I => \N__23115\
        );

    \I__3592\ : InMux
    port map (
            O => \N__23124\,
            I => \N__23110\
        );

    \I__3591\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23110\
        );

    \I__3590\ : Odrv12
    port map (
            O => \N__23120\,
            I => data_out_frame2_11_6
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__23115\,
            I => data_out_frame2_11_6
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__23110\,
            I => data_out_frame2_11_6
        );

    \I__3587\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23100\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__23100\,
            I => \c0.n18124\
        );

    \I__3585\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23094\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__23094\,
            I => \N__23091\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__23091\,
            I => \N__23088\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__23088\,
            I => \c0.data_out_frame2_19_0\
        );

    \I__3581\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23081\
        );

    \I__3580\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23078\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__23081\,
            I => data_out_frame2_18_0
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__23078\,
            I => data_out_frame2_18_0
        );

    \I__3577\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23070\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__23070\,
            I => \N__23067\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__23067\,
            I => \c0.n18160\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__23064\,
            I => \c0.tx2.n13614_cascade_\
        );

    \I__3573\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__3571\ : Span4Mux_v
    port map (
            O => \N__23055\,
            I => \N__23052\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__23052\,
            I => \N__23049\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__23049\,
            I => \c0.n17587\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__23046\,
            I => \N__23042\
        );

    \I__3567\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23039\
        );

    \I__3566\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23036\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__23039\,
            I => \N__23031\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__23031\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__23028\,
            I => \c0.n17107\
        );

    \I__3561\ : InMux
    port map (
            O => \N__23025\,
            I => \N__23020\
        );

    \I__3560\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23016\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__23023\,
            I => \N__23013\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__23020\,
            I => \N__23009\
        );

    \I__3557\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23006\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__23016\,
            I => \N__23003\
        );

    \I__3555\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23000\
        );

    \I__3554\ : InMux
    port map (
            O => \N__23012\,
            I => \N__22997\
        );

    \I__3553\ : Span4Mux_h
    port map (
            O => \N__23009\,
            I => \N__22994\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__22991\
        );

    \I__3551\ : Span4Mux_h
    port map (
            O => \N__23003\,
            I => \N__22988\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22985\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__22997\,
            I => data_out_frame2_15_6
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__22994\,
            I => data_out_frame2_15_6
        );

    \I__3547\ : Odrv12
    port map (
            O => \N__22991\,
            I => data_out_frame2_15_6
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__22988\,
            I => data_out_frame2_15_6
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__22985\,
            I => data_out_frame2_15_6
        );

    \I__3544\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22969\
        );

    \I__3543\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22966\
        );

    \I__3542\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22963\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22959\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22954\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22954\
        );

    \I__3538\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22951\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__22959\,
            I => \N__22946\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__22954\,
            I => \N__22946\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__22951\,
            I => data_out_frame2_12_6
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__22946\,
            I => data_out_frame2_12_6
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__22941\,
            I => \c0.n18118_cascade_\
        );

    \I__3532\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22934\
        );

    \I__3531\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22931\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22928\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__22931\,
            I => \N__22922\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__22928\,
            I => \N__22922\
        );

    \I__3527\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22918\
        );

    \I__3526\ : Span4Mux_v
    port map (
            O => \N__22922\,
            I => \N__22915\
        );

    \I__3525\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22912\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__22918\,
            I => data_out_frame2_13_6
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__22915\,
            I => data_out_frame2_13_6
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__22912\,
            I => data_out_frame2_13_6
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__22905\,
            I => \N__22902\
        );

    \I__3520\ : InMux
    port map (
            O => \N__22902\,
            I => \N__22899\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__22896\,
            I => \N__22893\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__22893\,
            I => \c0.n18121\
        );

    \I__3516\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__22884\,
            I => \c0.tx2.n13614\
        );

    \I__3513\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22875\
        );

    \I__3512\ : InMux
    port map (
            O => \N__22880\,
            I => \N__22875\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__22875\,
            I => n10976
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__22872\,
            I => \n10976_cascade_\
        );

    \I__3509\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22864\
        );

    \I__3508\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22859\
        );

    \I__3507\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22859\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__22864\,
            I => \r_Bit_Index_2_adj_2440\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__22859\,
            I => \r_Bit_Index_2_adj_2440\
        );

    \I__3504\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22849\
        );

    \I__3503\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22844\
        );

    \I__3502\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22844\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__22849\,
            I => \c0.rx.r_SM_Main_2_N_2094_0\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__22844\,
            I => \c0.rx.r_SM_Main_2_N_2094_0\
        );

    \I__3499\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__22836\,
            I => \c0.rx.n6_adj_2130\
        );

    \I__3497\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__22830\,
            I => \c0.n18247\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__22827\,
            I => \N__22824\
        );

    \I__3494\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22821\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22818\
        );

    \I__3492\ : Span4Mux_h
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__22815\,
            I => \c0.n22_adj_2372\
        );

    \I__3490\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22809\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__22809\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__3488\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__3486\ : Span4Mux_h
    port map (
            O => \N__22800\,
            I => \N__22797\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__22797\,
            I => \c0.n17620\
        );

    \I__3484\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__3482\ : Span12Mux_v
    port map (
            O => \N__22788\,
            I => \N__22785\
        );

    \I__3481\ : Odrv12
    port map (
            O => \N__22785\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__22782\,
            I => \N__22779\
        );

    \I__3479\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22776\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__22773\,
            I => \N__22770\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__22767\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__3474\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22758\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__22758\,
            I => \N__22755\
        );

    \I__3471\ : Span4Mux_h
    port map (
            O => \N__22755\,
            I => \N__22752\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__22752\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__22749\,
            I => \c0.tx2.n18082_cascade_\
        );

    \I__3468\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__3464\ : Odrv4
    port map (
            O => \N__22734\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__22731\,
            I => \c0.tx2.n18085_cascade_\
        );

    \I__3462\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22725\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__22725\,
            I => \c0.tx2.n18235\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__22722\,
            I => \c0.tx2.o_Tx_Serial_N_2062_cascade_\
        );

    \I__3459\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__3457\ : Span4Mux_v
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__22710\,
            I => n3
        );

    \I__3455\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22701\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__22701\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_27\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__3451\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22690\
        );

    \I__3450\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22687\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__22693\,
            I => \N__22684\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__22690\,
            I => \N__22680\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22677\
        );

    \I__3446\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22672\
        );

    \I__3445\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22672\
        );

    \I__3444\ : Sp12to4
    port map (
            O => \N__22680\,
            I => \N__22669\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__22677\,
            I => \N__22666\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__22672\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__3441\ : Odrv12
    port map (
            O => \N__22669\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__22666\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__3439\ : SRMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__3436\ : Span4Mux_s2_v
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__22647\,
            I => \c0.n3_adj_2236\
        );

    \I__3434\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22641\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__3432\ : Span4Mux_v
    port map (
            O => \N__22638\,
            I => \N__22635\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__22635\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_9\
        );

    \I__3430\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22627\
        );

    \I__3429\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22621\
        );

    \I__3428\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22621\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22618\
        );

    \I__3426\ : InMux
    port map (
            O => \N__22626\,
            I => \N__22615\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__22621\,
            I => \N__22612\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__22618\,
            I => \N__22609\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22606\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__22612\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__22609\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__22606\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__3419\ : SRMux
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__3417\ : Span4Mux_h
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__22590\,
            I => \c0.n3_adj_2274\
        );

    \I__3415\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__22584\,
            I => \c0.rx.n17636\
        );

    \I__3413\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__22578\,
            I => n17707
        );

    \I__3411\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22571\
        );

    \I__3410\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22568\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22565\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__22568\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__22565\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__3406\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22556\
        );

    \I__3405\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22550\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__22553\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__22550\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__3400\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22538\
        );

    \I__3399\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22535\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22532\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__22535\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__22532\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__3395\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22524\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__22524\,
            I => \c0.rx.n6\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__22521\,
            I => \c0.rx.n17022_cascade_\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__22518\,
            I => \c0.rx.r_SM_Main_2_N_2094_0_cascade_\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__22515\,
            I => \c0.rx.n17380_cascade_\
        );

    \I__3390\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22509\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__22509\,
            I => \c0.rx.n17635\
        );

    \I__3388\ : InMux
    port map (
            O => \N__22506\,
            I => \N__22503\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22500\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__22500\,
            I => \c0.n40\
        );

    \I__3385\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22494\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22491\
        );

    \I__3383\ : Span4Mux_h
    port map (
            O => \N__22491\,
            I => \N__22488\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__22488\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_24\
        );

    \I__3381\ : SRMux
    port map (
            O => \N__22485\,
            I => \N__22482\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__22482\,
            I => \N__22479\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__22479\,
            I => \c0.n3_adj_2242\
        );

    \I__3378\ : SRMux
    port map (
            O => \N__22476\,
            I => \N__22473\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__3376\ : Span4Mux_v
    port map (
            O => \N__22470\,
            I => \N__22467\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__22467\,
            I => \c0.n3_adj_2240\
        );

    \I__3374\ : SRMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__22458\,
            I => \N__22455\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__22455\,
            I => \c0.n3_adj_2234\
        );

    \I__3370\ : SRMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22446\
        );

    \I__3368\ : Span4Mux_h
    port map (
            O => \N__22446\,
            I => \N__22443\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__22443\,
            I => \c0.n3_adj_2230\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__22440\,
            I => \c0.n10009_cascade_\
        );

    \I__3365\ : SRMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__3363\ : Span4Mux_v
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__22428\,
            I => \c0.n3_adj_2181\
        );

    \I__3361\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22422\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__22419\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_18\
        );

    \I__3358\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22413\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__22413\,
            I => \N__22410\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__22410\,
            I => \c0.n42\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__22407\,
            I => \c0.n41_adj_2376_cascade_\
        );

    \I__3354\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22401\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__22401\,
            I => \c0.n39_adj_2377\
        );

    \I__3352\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22395\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__22389\,
            I => \c0.n43_adj_2380\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__22386\,
            I => \c0.n48_adj_2379_cascade_\
        );

    \I__3347\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22380\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__22380\,
            I => \c0.n44_adj_2378\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__22377\,
            I => \c0.n9995_cascade_\
        );

    \I__3344\ : InMux
    port map (
            O => \N__22374\,
            I => \N__22370\
        );

    \I__3343\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22367\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__22370\,
            I => \c0.n9995\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__22367\,
            I => \c0.n9995\
        );

    \I__3340\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22359\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__22356\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_2\
        );

    \I__3337\ : SRMux
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__22350\,
            I => \N__22347\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__22347\,
            I => \c0.n3_adj_2286\
        );

    \I__3334\ : SRMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__3332\ : Span4Mux_v
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__3331\ : Odrv4
    port map (
            O => \N__22335\,
            I => \c0.n3_adj_2226\
        );

    \I__3330\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__22326\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_2\
        );

    \I__3327\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22319\
        );

    \I__3326\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22316\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22313\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__22316\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__22313\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__3322\ : InMux
    port map (
            O => \N__22308\,
            I => \c0.tx2.n16134\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__22305\,
            I => \N__22301\
        );

    \I__3320\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22298\
        );

    \I__3319\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22295\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__22298\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__22295\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__3316\ : InMux
    port map (
            O => \N__22290\,
            I => \c0.tx2.n16135\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__3314\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22277\
        );

    \I__3313\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22277\
        );

    \I__3312\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22274\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22271\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__22274\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__22271\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__3308\ : InMux
    port map (
            O => \N__22266\,
            I => \c0.tx2.n16136\
        );

    \I__3307\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22259\
        );

    \I__3306\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22256\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__22259\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__22256\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__3303\ : InMux
    port map (
            O => \N__22251\,
            I => \c0.tx2.n16137\
        );

    \I__3302\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22244\
        );

    \I__3301\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22241\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__22244\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__22241\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__3298\ : InMux
    port map (
            O => \N__22236\,
            I => \c0.tx2.n16138\
        );

    \I__3297\ : InMux
    port map (
            O => \N__22233\,
            I => \bfn_6_25_0_\
        );

    \I__3296\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22226\
        );

    \I__3295\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22223\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__22226\,
            I => \N__22220\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__22223\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__22220\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__3291\ : SRMux
    port map (
            O => \N__22215\,
            I => \N__22211\
        );

    \I__3290\ : SRMux
    port map (
            O => \N__22214\,
            I => \N__22208\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__22211\,
            I => \N__22205\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__22208\,
            I => \N__22202\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__22205\,
            I => \N__22199\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__22202\,
            I => \c0.tx2.n10852\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__22199\,
            I => \c0.tx2.n10852\
        );

    \I__3284\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22189\
        );

    \I__3283\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22186\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__22192\,
            I => \N__22183\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22177\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__22186\,
            I => \N__22177\
        );

    \I__3279\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22174\
        );

    \I__3278\ : InMux
    port map (
            O => \N__22182\,
            I => \N__22171\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__22177\,
            I => \N__22166\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__22174\,
            I => \N__22166\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22163\
        );

    \I__3274\ : Span4Mux_h
    port map (
            O => \N__22166\,
            I => \N__22160\
        );

    \I__3273\ : Span4Mux_v
    port map (
            O => \N__22163\,
            I => \N__22157\
        );

    \I__3272\ : Span4Mux_s0_h
    port map (
            O => \N__22160\,
            I => \N__22154\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__22157\,
            I => \N__22151\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__22154\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__22151\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__22146\,
            I => \N__22142\
        );

    \I__3267\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22139\
        );

    \I__3266\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22136\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__22139\,
            I => \c0.tx2.n10\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__22136\,
            I => \c0.tx2.n10\
        );

    \I__3263\ : IoInMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__3261\ : IoSpan4Mux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__3260\ : Span4Mux_s2_h
    port map (
            O => \N__22122\,
            I => \N__22118\
        );

    \I__3259\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22115\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__22118\,
            I => \N__22109\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22109\
        );

    \I__3256\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22106\
        );

    \I__3255\ : Span4Mux_v
    port map (
            O => \N__22109\,
            I => \N__22103\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__22106\,
            I => \N__22100\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__22103\,
            I => tx2_o
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__22100\,
            I => tx2_o
        );

    \I__3251\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22090\
        );

    \I__3250\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22087\
        );

    \I__3249\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22084\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__22090\,
            I => \N__22081\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__22087\,
            I => data_out_frame2_14_7
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__22084\,
            I => data_out_frame2_14_7
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__22081\,
            I => data_out_frame2_14_7
        );

    \I__3244\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22071\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__22071\,
            I => \c0.tx2.n17322\
        );

    \I__3242\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22062\
        );

    \I__3241\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22062\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__22062\,
            I => \c0.tx2.n17018\
        );

    \I__3239\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22055\
        );

    \I__3238\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22052\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__22055\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__22052\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__3235\ : InMux
    port map (
            O => \N__22047\,
            I => \bfn_6_24_0_\
        );

    \I__3234\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22037\
        );

    \I__3233\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22037\
        );

    \I__3232\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22034\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22031\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__22034\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__22031\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__3228\ : InMux
    port map (
            O => \N__22026\,
            I => \c0.tx2.n16132\
        );

    \I__3227\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22019\
        );

    \I__3226\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22016\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__22019\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__22016\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__3223\ : InMux
    port map (
            O => \N__22011\,
            I => \c0.tx2.n16133\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__22008\,
            I => \c0.tx2.n13748_cascade_\
        );

    \I__3221\ : InMux
    port map (
            O => \N__22005\,
            I => \N__22002\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__22002\,
            I => \N__21998\
        );

    \I__3219\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21995\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__21998\,
            I => \N__21992\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__21995\,
            I => \N__21987\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__21992\,
            I => \N__21987\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__21987\,
            I => data_out_frame2_18_7
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__21984\,
            I => \N__21981\
        );

    \I__3213\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21974\
        );

    \I__3211\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21971\
        );

    \I__3210\ : Span4Mux_h
    port map (
            O => \N__21974\,
            I => \N__21968\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__21971\,
            I => data_out_frame2_17_2
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__21968\,
            I => data_out_frame2_17_2
        );

    \I__3207\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21959\
        );

    \I__3206\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21952\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21949\
        );

    \I__3204\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21946\
        );

    \I__3203\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21943\
        );

    \I__3202\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21940\
        );

    \I__3201\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21937\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__21952\,
            I => \N__21934\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__21949\,
            I => \N__21931\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__21946\,
            I => \N__21928\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__21943\,
            I => \N__21925\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__21940\,
            I => \N__21922\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__21937\,
            I => \N__21919\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__21934\,
            I => \N__21914\
        );

    \I__3193\ : Span4Mux_v
    port map (
            O => \N__21931\,
            I => \N__21914\
        );

    \I__3192\ : Span12Mux_v
    port map (
            O => \N__21928\,
            I => \N__21911\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__21925\,
            I => \N__21906\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__21922\,
            I => \N__21906\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__21919\,
            I => data_out_frame2_7_5
        );

    \I__3188\ : Odrv4
    port map (
            O => \N__21914\,
            I => data_out_frame2_7_5
        );

    \I__3187\ : Odrv12
    port map (
            O => \N__21911\,
            I => data_out_frame2_7_5
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__21906\,
            I => data_out_frame2_7_5
        );

    \I__3185\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21890\
        );

    \I__3184\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21887\
        );

    \I__3183\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21882\
        );

    \I__3182\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21882\
        );

    \I__3181\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21879\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__21890\,
            I => data_out_frame2_11_4
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__21887\,
            I => data_out_frame2_11_4
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__21882\,
            I => data_out_frame2_11_4
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__21879\,
            I => data_out_frame2_11_4
        );

    \I__3176\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21861\
        );

    \I__3175\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21861\
        );

    \I__3174\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21857\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__21867\,
            I => \N__21854\
        );

    \I__3172\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21851\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21848\
        );

    \I__3170\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21845\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21842\
        );

    \I__3168\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21839\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__21851\,
            I => data_out_frame2_11_5
        );

    \I__3166\ : Odrv12
    port map (
            O => \N__21848\,
            I => data_out_frame2_11_5
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__21845\,
            I => data_out_frame2_11_5
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__21842\,
            I => data_out_frame2_11_5
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__21839\,
            I => data_out_frame2_11_5
        );

    \I__3162\ : InMux
    port map (
            O => \N__21828\,
            I => \N__21825\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__21825\,
            I => \N__21821\
        );

    \I__3160\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21817\
        );

    \I__3159\ : Span4Mux_s1_h
    port map (
            O => \N__21821\,
            I => \N__21814\
        );

    \I__3158\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21811\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__21817\,
            I => \N__21808\
        );

    \I__3156\ : Span4Mux_h
    port map (
            O => \N__21814\,
            I => \N__21805\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21800\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__21808\,
            I => \N__21800\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__21805\,
            I => \c0.n10359\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__21800\,
            I => \c0.n10359\
        );

    \I__3151\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21791\
        );

    \I__3150\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21788\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__21791\,
            I => \N__21784\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21780\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__21787\,
            I => \N__21777\
        );

    \I__3146\ : Span4Mux_s2_h
    port map (
            O => \N__21784\,
            I => \N__21774\
        );

    \I__3145\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21771\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__21780\,
            I => \N__21768\
        );

    \I__3143\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21765\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__21774\,
            I => \N__21762\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__21771\,
            I => data_out_frame2_5_4
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__21768\,
            I => data_out_frame2_5_4
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__21765\,
            I => data_out_frame2_5_4
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__21762\,
            I => data_out_frame2_5_4
        );

    \I__3137\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21749\
        );

    \I__3136\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21746\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21742\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__21746\,
            I => \N__21737\
        );

    \I__3133\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21734\
        );

    \I__3132\ : Span4Mux_h
    port map (
            O => \N__21742\,
            I => \N__21731\
        );

    \I__3131\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21726\
        );

    \I__3130\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21726\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__21737\,
            I => data_out_frame2_10_7
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__21734\,
            I => data_out_frame2_10_7
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__21731\,
            I => data_out_frame2_10_7
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__21726\,
            I => data_out_frame2_10_7
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__21717\,
            I => \N__21714\
        );

    \I__3124\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21710\
        );

    \I__3123\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21707\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21704\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__21707\,
            I => data_out_frame2_17_0
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__21704\,
            I => data_out_frame2_17_0
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__21699\,
            I => \N__21696\
        );

    \I__3118\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21693\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__3116\ : Odrv12
    port map (
            O => \N__21690\,
            I => \c0.n18163\
        );

    \I__3115\ : InMux
    port map (
            O => \N__21687\,
            I => \N__21684\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__21684\,
            I => \c0.n18208\
        );

    \I__3113\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21677\
        );

    \I__3112\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21674\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21671\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__21674\,
            I => data_out_frame2_17_3
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__21671\,
            I => data_out_frame2_17_3
        );

    \I__3108\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21661\
        );

    \I__3107\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21657\
        );

    \I__3106\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21654\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21651\
        );

    \I__3104\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21648\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__21657\,
            I => \N__21645\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__21654\,
            I => \N__21642\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__21651\,
            I => \N__21639\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__21648\,
            I => data_out_frame2_14_2
        );

    \I__3099\ : Odrv12
    port map (
            O => \N__21645\,
            I => data_out_frame2_14_2
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__21642\,
            I => data_out_frame2_14_2
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__21639\,
            I => data_out_frame2_14_2
        );

    \I__3096\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21627\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__3094\ : Span4Mux_h
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__3093\ : Span4Mux_h
    port map (
            O => \N__21621\,
            I => \N__21618\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__21618\,
            I => \c0.n10_adj_2207\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__3090\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21609\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__21609\,
            I => \N__21606\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__21606\,
            I => \N__21603\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__21603\,
            I => \c0.n18061\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__21600\,
            I => \c0.n18256_cascade_\
        );

    \I__3085\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21594\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__21594\,
            I => \c0.n6_adj_2139\
        );

    \I__3083\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21588\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__21588\,
            I => \c0.n22_adj_2371\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__21585\,
            I => \c0.n18259_cascade_\
        );

    \I__3080\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21579\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__21576\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__3077\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21568\
        );

    \I__3076\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21565\
        );

    \I__3075\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21561\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__21568\,
            I => \N__21558\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__21565\,
            I => \N__21555\
        );

    \I__3072\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21552\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21547\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__21558\,
            I => \N__21547\
        );

    \I__3069\ : Span4Mux_h
    port map (
            O => \N__21555\,
            I => \N__21544\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__21552\,
            I => data_out_frame2_10_1
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__21547\,
            I => data_out_frame2_10_1
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__21544\,
            I => data_out_frame2_10_1
        );

    \I__3065\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21534\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__21534\,
            I => \N__21531\
        );

    \I__3063\ : Span4Mux_h
    port map (
            O => \N__21531\,
            I => \N__21528\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__21528\,
            I => \c0.n17203\
        );

    \I__3061\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21519\
        );

    \I__3060\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21516\
        );

    \I__3059\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21513\
        );

    \I__3058\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21510\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__21519\,
            I => \N__21506\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__21516\,
            I => \N__21503\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__21513\,
            I => \N__21500\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__21510\,
            I => \N__21497\
        );

    \I__3053\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21494\
        );

    \I__3052\ : Span4Mux_h
    port map (
            O => \N__21506\,
            I => \N__21491\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__21503\,
            I => \N__21486\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__21500\,
            I => \N__21486\
        );

    \I__3049\ : Span4Mux_h
    port map (
            O => \N__21497\,
            I => \N__21483\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__21494\,
            I => data_out_frame2_8_6
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__21491\,
            I => data_out_frame2_8_6
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__21486\,
            I => data_out_frame2_8_6
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__21483\,
            I => data_out_frame2_8_6
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__21474\,
            I => \N__21471\
        );

    \I__3043\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21468\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21464\
        );

    \I__3041\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21461\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__21464\,
            I => \N__21458\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21453\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__21458\,
            I => \N__21450\
        );

    \I__3037\ : InMux
    port map (
            O => \N__21457\,
            I => \N__21447\
        );

    \I__3036\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21444\
        );

    \I__3035\ : Span4Mux_s3_h
    port map (
            O => \N__21453\,
            I => \N__21441\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__21450\,
            I => \N__21436\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__21447\,
            I => \N__21436\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__21444\,
            I => data_out_frame2_9_6
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__21441\,
            I => data_out_frame2_9_6
        );

    \I__3030\ : Odrv4
    port map (
            O => \N__21436\,
            I => data_out_frame2_9_6
        );

    \I__3029\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21426\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__21423\,
            I => \N__21420\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__21420\,
            I => \c0.n18127\
        );

    \I__3025\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21413\
        );

    \I__3024\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21410\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__21413\,
            I => data_out_frame2_18_3
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__21410\,
            I => data_out_frame2_18_3
        );

    \I__3021\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21402\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__21402\,
            I => \c0.n22_adj_2387\
        );

    \I__3019\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21396\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__21396\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__3017\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21390\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__3015\ : Odrv12
    port map (
            O => \N__21387\,
            I => \c0.n18157\
        );

    \I__3014\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__21381\,
            I => \c0.n17603\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__21378\,
            I => \c0.n18226_cascade_\
        );

    \I__3011\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21372\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__21372\,
            I => \c0.n18229\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__21369\,
            I => \N__21365\
        );

    \I__3008\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21361\
        );

    \I__3007\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21354\
        );

    \I__3006\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21354\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21350\
        );

    \I__3004\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21347\
        );

    \I__3003\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21344\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__21354\,
            I => \N__21341\
        );

    \I__3001\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21338\
        );

    \I__3000\ : Span4Mux_v
    port map (
            O => \N__21350\,
            I => \N__21335\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__21347\,
            I => data_out_frame2_10_0
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__21344\,
            I => data_out_frame2_10_0
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__21341\,
            I => data_out_frame2_10_0
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__21338\,
            I => data_out_frame2_10_0
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__21335\,
            I => data_out_frame2_10_0
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__21324\,
            I => \c0.n18148_cascade_\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__21321\,
            I => \N__21318\
        );

    \I__2992\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21315\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__21315\,
            I => \c0.n18151\
        );

    \I__2990\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21308\
        );

    \I__2989\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21305\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21301\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21297\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__21304\,
            I => \N__21294\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__21301\,
            I => \N__21290\
        );

    \I__2984\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21287\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__21297\,
            I => \N__21284\
        );

    \I__2982\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21279\
        );

    \I__2981\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21279\
        );

    \I__2980\ : Span4Mux_v
    port map (
            O => \N__21290\,
            I => \N__21274\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21274\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__21284\,
            I => data_out_frame2_5_0
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__21279\,
            I => data_out_frame2_5_0
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__21274\,
            I => data_out_frame2_5_0
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__2974\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21261\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__21261\,
            I => \N__21258\
        );

    \I__2972\ : Span4Mux_h
    port map (
            O => \N__21258\,
            I => \N__21255\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__21252\,
            I => \N__21249\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__21249\,
            I => \c0.n5_adj_2217\
        );

    \I__2968\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21243\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__21243\,
            I => \c0.n6_adj_2143\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__2965\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__2963\ : Odrv12
    port map (
            O => \N__21231\,
            I => \c0.data_out_frame2_19_3\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__21228\,
            I => \c0.n18052_cascade_\
        );

    \I__2961\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__2959\ : Odrv12
    port map (
            O => \N__21219\,
            I => \c0.data_out_frame2_20_3\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__21216\,
            I => \c0.n18055_cascade_\
        );

    \I__2957\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21207\
        );

    \I__2956\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21204\
        );

    \I__2955\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21200\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21196\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21191\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__21204\,
            I => \N__21188\
        );

    \I__2951\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21185\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__21200\,
            I => \N__21182\
        );

    \I__2949\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21179\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21176\
        );

    \I__2947\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21173\
        );

    \I__2946\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21170\
        );

    \I__2945\ : Span4Mux_v
    port map (
            O => \N__21191\,
            I => \N__21167\
        );

    \I__2944\ : Span4Mux_s3_h
    port map (
            O => \N__21188\,
            I => \N__21162\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__21185\,
            I => \N__21162\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__21182\,
            I => \N__21153\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21153\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__21176\,
            I => \N__21153\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__21173\,
            I => \N__21153\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N__21150\
        );

    \I__2937\ : Span4Mux_s3_h
    port map (
            O => \N__21167\,
            I => \N__21145\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__21162\,
            I => \N__21145\
        );

    \I__2935\ : Span4Mux_h
    port map (
            O => \N__21153\,
            I => \N__21142\
        );

    \I__2934\ : Odrv12
    port map (
            O => \N__21150\,
            I => \c0.n9157\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__21145\,
            I => \c0.n9157\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__21142\,
            I => \c0.n9157\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__21135\,
            I => \n17708_cascade_\
        );

    \I__2930\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21128\
        );

    \I__2929\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21125\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__21128\,
            I => n5244
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__21125\,
            I => n5244
        );

    \I__2926\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21116\
        );

    \I__2925\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21113\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__21116\,
            I => n11018
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__21113\,
            I => n11018
        );

    \I__2922\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__21105\,
            I => \c0.data_out_frame2_20_0\
        );

    \I__2920\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__21090\,
            I => \c0.n18049\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__2914\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21081\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__21081\,
            I => \N__21078\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__21078\,
            I => \N__21075\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__21075\,
            I => \c0.n18043\
        );

    \I__2910\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21069\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__2908\ : Span4Mux_h
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__21063\,
            I => \c0.n17586\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__21060\,
            I => \c0.n18244_cascade_\
        );

    \I__2905\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__21054\,
            I => \c0.n6_adj_2140\
        );

    \I__2903\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__2901\ : Odrv12
    port map (
            O => \N__21045\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__21042\,
            I => \c0.tx2.n18232_cascade_\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__2898\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__21033\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_31\
        );

    \I__2896\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21027\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__21027\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_25\
        );

    \I__2894\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__21021\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_26\
        );

    \I__2892\ : SRMux
    port map (
            O => \N__21018\,
            I => \N__21015\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__21012\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__21012\,
            I => \c0.rx.n10845\
        );

    \I__2889\ : InMux
    port map (
            O => \N__21009\,
            I => \N__21006\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__21006\,
            I => n1
        );

    \I__2887\ : InMux
    port map (
            O => \N__21003\,
            I => \N__20999\
        );

    \I__2886\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20996\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__20999\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__20996\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__2883\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20987\
        );

    \I__2882\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20984\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__20987\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__20984\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__2879\ : CEMux
    port map (
            O => \N__20979\,
            I => \N__20976\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__20976\,
            I => \N__20973\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__20973\,
            I => \N__20970\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__20970\,
            I => \c0.rx.n10656\
        );

    \I__2875\ : SRMux
    port map (
            O => \N__20967\,
            I => \N__20964\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__20964\,
            I => \N__20961\
        );

    \I__2873\ : Span4Mux_s1_h
    port map (
            O => \N__20961\,
            I => \N__20958\
        );

    \I__2872\ : Span4Mux_h
    port map (
            O => \N__20958\,
            I => \N__20955\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__20955\,
            I => \c0.n3_adj_2244\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__20952\,
            I => \N__20949\
        );

    \I__2869\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20943\
        );

    \I__2868\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20936\
        );

    \I__2867\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20936\
        );

    \I__2866\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20936\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20933\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20930\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__20933\,
            I => \N__20927\
        );

    \I__2862\ : Span12Mux_h
    port map (
            O => \N__20930\,
            I => \N__20924\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__20927\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__2860\ : Odrv12
    port map (
            O => \N__20924\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__2859\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20916\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__20916\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_21\
        );

    \I__2857\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20910\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__20910\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_27\
        );

    \I__2855\ : SRMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__20901\,
            I => \N__20898\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__20895\,
            I => \c0.n3_adj_2276\
        );

    \I__2850\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__20889\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_8\
        );

    \I__2848\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20883\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__20883\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_9\
        );

    \I__2846\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20874\
        );

    \I__2845\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20867\
        );

    \I__2844\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20867\
        );

    \I__2843\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20867\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__20874\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__20867\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__2840\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__20859\,
            I => \c0.n41\
        );

    \I__2838\ : SRMux
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__2836\ : Span4Mux_s1_h
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__20844\,
            I => \c0.n3_adj_2261\
        );

    \I__2833\ : SRMux
    port map (
            O => \N__20841\,
            I => \N__20838\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__20838\,
            I => \N__20835\
        );

    \I__2831\ : Span4Mux_s1_h
    port map (
            O => \N__20835\,
            I => \N__20832\
        );

    \I__2830\ : Span4Mux_h
    port map (
            O => \N__20832\,
            I => \N__20829\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__20829\,
            I => \c0.n3_adj_2270\
        );

    \I__2828\ : SRMux
    port map (
            O => \N__20826\,
            I => \N__20823\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__2826\ : Span4Mux_s2_h
    port map (
            O => \N__20820\,
            I => \N__20817\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__20817\,
            I => \c0.n3_adj_2252\
        );

    \I__2824\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__20811\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_17\
        );

    \I__2822\ : SRMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__20802\,
            I => \c0.n3_adj_2257\
        );

    \I__2819\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20793\
        );

    \I__2818\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20786\
        );

    \I__2817\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20786\
        );

    \I__2816\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20786\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__20793\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__20786\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__2813\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20775\
        );

    \I__2811\ : Span4Mux_v
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__20772\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_17\
        );

    \I__2809\ : SRMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__20766\,
            I => \N__20763\
        );

    \I__2807\ : Span12Mux_s4_h
    port map (
            O => \N__20763\,
            I => \N__20760\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__20760\,
            I => \c0.n3_adj_2248\
        );

    \I__2805\ : SRMux
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__20754\,
            I => \N__20751\
        );

    \I__2803\ : Span4Mux_s1_h
    port map (
            O => \N__20751\,
            I => \N__20748\
        );

    \I__2802\ : Span4Mux_h
    port map (
            O => \N__20748\,
            I => \N__20745\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__20745\,
            I => \c0.n3_adj_2250\
        );

    \I__2800\ : InMux
    port map (
            O => \N__20742\,
            I => n16005
        );

    \I__2799\ : InMux
    port map (
            O => \N__20739\,
            I => n16006
        );

    \I__2798\ : InMux
    port map (
            O => \N__20736\,
            I => n16007
        );

    \I__2797\ : InMux
    port map (
            O => \N__20733\,
            I => n16008
        );

    \I__2796\ : InMux
    port map (
            O => \N__20730\,
            I => n16009
        );

    \I__2795\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20724\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__20724\,
            I => \c0.n3\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__20721\,
            I => \c0.n26_adj_2373_cascade_\
        );

    \I__2792\ : SRMux
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__20715\,
            I => \N__20712\
        );

    \I__2790\ : Sp12to4
    port map (
            O => \N__20712\,
            I => \N__20709\
        );

    \I__2789\ : Odrv12
    port map (
            O => \N__20709\,
            I => \c0.n3_adj_2280\
        );

    \I__2788\ : InMux
    port map (
            O => \N__20706\,
            I => n15996
        );

    \I__2787\ : InMux
    port map (
            O => \N__20703\,
            I => n15997
        );

    \I__2786\ : InMux
    port map (
            O => \N__20700\,
            I => n15998
        );

    \I__2785\ : InMux
    port map (
            O => \N__20697\,
            I => n15999
        );

    \I__2784\ : InMux
    port map (
            O => \N__20694\,
            I => n16000
        );

    \I__2783\ : InMux
    port map (
            O => \N__20691\,
            I => n16001
        );

    \I__2782\ : InMux
    port map (
            O => \N__20688\,
            I => \bfn_5_26_0_\
        );

    \I__2781\ : InMux
    port map (
            O => \N__20685\,
            I => n16003
        );

    \I__2780\ : InMux
    port map (
            O => \N__20682\,
            I => n16004
        );

    \I__2779\ : InMux
    port map (
            O => \N__20679\,
            I => n15987
        );

    \I__2778\ : InMux
    port map (
            O => \N__20676\,
            I => n15988
        );

    \I__2777\ : InMux
    port map (
            O => \N__20673\,
            I => n15989
        );

    \I__2776\ : InMux
    port map (
            O => \N__20670\,
            I => n15990
        );

    \I__2775\ : InMux
    port map (
            O => \N__20667\,
            I => n15991
        );

    \I__2774\ : InMux
    port map (
            O => \N__20664\,
            I => n15992
        );

    \I__2773\ : InMux
    port map (
            O => \N__20661\,
            I => n15993
        );

    \I__2772\ : InMux
    port map (
            O => \N__20658\,
            I => \bfn_5_25_0_\
        );

    \I__2771\ : InMux
    port map (
            O => \N__20655\,
            I => n15995
        );

    \I__2770\ : InMux
    port map (
            O => \N__20652\,
            I => \bfn_5_23_0_\
        );

    \I__2769\ : InMux
    port map (
            O => \N__20649\,
            I => n15979
        );

    \I__2768\ : InMux
    port map (
            O => \N__20646\,
            I => n15980
        );

    \I__2767\ : InMux
    port map (
            O => \N__20643\,
            I => n15981
        );

    \I__2766\ : InMux
    port map (
            O => \N__20640\,
            I => n15982
        );

    \I__2765\ : InMux
    port map (
            O => \N__20637\,
            I => n15983
        );

    \I__2764\ : InMux
    port map (
            O => \N__20634\,
            I => n15984
        );

    \I__2763\ : InMux
    port map (
            O => \N__20631\,
            I => n15985
        );

    \I__2762\ : InMux
    port map (
            O => \N__20628\,
            I => \bfn_5_24_0_\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__20625\,
            I => \N__20621\
        );

    \I__2760\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20616\
        );

    \I__2759\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20613\
        );

    \I__2758\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20609\
        );

    \I__2757\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20606\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20601\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__20613\,
            I => \N__20601\
        );

    \I__2754\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20598\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20595\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__20606\,
            I => \N__20592\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20589\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__20598\,
            I => data_out_frame2_15_2
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__20595\,
            I => data_out_frame2_15_2
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__20592\,
            I => data_out_frame2_15_2
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__20589\,
            I => data_out_frame2_15_2
        );

    \I__2746\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20573\
        );

    \I__2744\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20570\
        );

    \I__2743\ : Span4Mux_s3_h
    port map (
            O => \N__20573\,
            I => \N__20567\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__20570\,
            I => data_out_frame2_18_2
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__20567\,
            I => data_out_frame2_18_2
        );

    \I__2740\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20558\
        );

    \I__2739\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20554\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__20558\,
            I => \N__20551\
        );

    \I__2737\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20548\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__20554\,
            I => \N__20544\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__20551\,
            I => \N__20539\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20539\
        );

    \I__2733\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20536\
        );

    \I__2732\ : Span4Mux_h
    port map (
            O => \N__20544\,
            I => \N__20531\
        );

    \I__2731\ : Span4Mux_h
    port map (
            O => \N__20539\,
            I => \N__20531\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__20536\,
            I => data_out_frame2_16_5
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__20531\,
            I => data_out_frame2_16_5
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__20526\,
            I => \N__20522\
        );

    \I__2727\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20518\
        );

    \I__2726\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20514\
        );

    \I__2725\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20510\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__20518\,
            I => \N__20507\
        );

    \I__2723\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20504\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20501\
        );

    \I__2721\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20498\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__20510\,
            I => \N__20495\
        );

    \I__2719\ : Span4Mux_s2_h
    port map (
            O => \N__20507\,
            I => \N__20490\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20490\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__20501\,
            I => \N__20487\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__20498\,
            I => data_out_frame2_15_4
        );

    \I__2715\ : Odrv12
    port map (
            O => \N__20495\,
            I => data_out_frame2_15_4
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__20490\,
            I => data_out_frame2_15_4
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__20487\,
            I => data_out_frame2_15_4
        );

    \I__2712\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20475\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__20475\,
            I => \N__20471\
        );

    \I__2710\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20468\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__20471\,
            I => \c0.n17156\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__20468\,
            I => \c0.n17156\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__20463\,
            I => \c0.n6_adj_2182_cascade_\
        );

    \I__2706\ : InMux
    port map (
            O => \N__20460\,
            I => \N__20457\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__20454\,
            I => \N__20450\
        );

    \I__2703\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20447\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__20450\,
            I => \c0.n10229\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__20447\,
            I => \c0.n10229\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__20442\,
            I => \n10725_cascade_\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__20439\,
            I => \N__20435\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__20438\,
            I => \N__20432\
        );

    \I__2697\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20428\
        );

    \I__2696\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20425\
        );

    \I__2695\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20421\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__20428\,
            I => \N__20418\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__20425\,
            I => \N__20415\
        );

    \I__2692\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20412\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__20421\,
            I => \N__20409\
        );

    \I__2690\ : Span4Mux_s1_h
    port map (
            O => \N__20418\,
            I => \N__20404\
        );

    \I__2689\ : Span4Mux_v
    port map (
            O => \N__20415\,
            I => \N__20404\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__20412\,
            I => data_out_frame2_12_7
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__20409\,
            I => data_out_frame2_12_7
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__20404\,
            I => data_out_frame2_12_7
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20392\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20389\
        );

    \I__2683\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20386\
        );

    \I__2682\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20383\
        );

    \I__2681\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20380\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__20386\,
            I => \N__20376\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__20383\,
            I => \N__20373\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__20380\,
            I => \N__20370\
        );

    \I__2677\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20367\
        );

    \I__2676\ : Span4Mux_h
    port map (
            O => \N__20376\,
            I => \N__20364\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__20373\,
            I => \N__20359\
        );

    \I__2674\ : Span4Mux_s1_h
    port map (
            O => \N__20370\,
            I => \N__20359\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__20367\,
            I => data_out_frame2_10_3
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__20364\,
            I => data_out_frame2_10_3
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__20359\,
            I => data_out_frame2_10_3
        );

    \I__2670\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20349\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20346\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__20343\,
            I => \c0.n18106\
        );

    \I__2666\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20336\
        );

    \I__2665\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20333\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20327\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__20333\,
            I => \N__20327\
        );

    \I__2662\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20324\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__20327\,
            I => \N__20319\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20316\
        );

    \I__2659\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20313\
        );

    \I__2658\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20310\
        );

    \I__2657\ : Span4Mux_s2_h
    port map (
            O => \N__20319\,
            I => \N__20307\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__20316\,
            I => \N__20304\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__20313\,
            I => \N__20301\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__20310\,
            I => data_out_frame2_16_2
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__20307\,
            I => data_out_frame2_16_2
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__20304\,
            I => data_out_frame2_16_2
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__20301\,
            I => data_out_frame2_16_2
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__2649\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20285\
        );

    \I__2648\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20281\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__20285\,
            I => \N__20278\
        );

    \I__2646\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20275\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20272\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__20278\,
            I => \c0.n10263\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__20275\,
            I => \c0.n10263\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__20272\,
            I => \c0.n10263\
        );

    \I__2641\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20262\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__20262\,
            I => \N__20259\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__20259\,
            I => \c0.n15_adj_2205\
        );

    \I__2638\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20250\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__20250\,
            I => \N__20247\
        );

    \I__2635\ : Span4Mux_h
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__20244\,
            I => \c0.n5_adj_2337\
        );

    \I__2633\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20235\
        );

    \I__2632\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20235\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__20235\,
            I => \N__20231\
        );

    \I__2630\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20226\
        );

    \I__2629\ : Span4Mux_s3_h
    port map (
            O => \N__20231\,
            I => \N__20223\
        );

    \I__2628\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20220\
        );

    \I__2627\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20217\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__20226\,
            I => data_out_frame2_10_2
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__20223\,
            I => data_out_frame2_10_2
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__20220\,
            I => data_out_frame2_10_2
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__20217\,
            I => data_out_frame2_10_2
        );

    \I__2622\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20204\
        );

    \I__2621\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20201\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__20204\,
            I => \N__20198\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__20201\,
            I => \N__20195\
        );

    \I__2618\ : Span4Mux_s3_h
    port map (
            O => \N__20198\,
            I => \N__20190\
        );

    \I__2617\ : Span4Mux_v
    port map (
            O => \N__20195\,
            I => \N__20190\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__20190\,
            I => \c0.n10492\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__2614\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20179\
        );

    \I__2613\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20174\
        );

    \I__2612\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20174\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__20179\,
            I => \N__20171\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__20174\,
            I => \N__20168\
        );

    \I__2609\ : Span4Mux_s2_h
    port map (
            O => \N__20171\,
            I => \N__20161\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__20168\,
            I => \N__20161\
        );

    \I__2607\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20158\
        );

    \I__2606\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20155\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__20161\,
            I => \N__20152\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__20158\,
            I => data_out_frame2_12_5
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__20155\,
            I => data_out_frame2_12_5
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__20152\,
            I => data_out_frame2_12_5
        );

    \I__2601\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20142\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__20139\,
            I => \N__20135\
        );

    \I__2598\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20132\
        );

    \I__2597\ : Span4Mux_s1_h
    port map (
            O => \N__20135\,
            I => \N__20129\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__20132\,
            I => \c0.n17255\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__20129\,
            I => \c0.n17255\
        );

    \I__2594\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20120\
        );

    \I__2593\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20117\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__20120\,
            I => \N__20114\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20110\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__20114\,
            I => \N__20107\
        );

    \I__2589\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20103\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__20110\,
            I => \N__20098\
        );

    \I__2587\ : Span4Mux_s2_h
    port map (
            O => \N__20107\,
            I => \N__20098\
        );

    \I__2586\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20095\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__20103\,
            I => data_out_frame2_16_4
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__20098\,
            I => data_out_frame2_16_4
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__20095\,
            I => data_out_frame2_16_4
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__20088\,
            I => \N__20084\
        );

    \I__2581\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20081\
        );

    \I__2580\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20077\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20074\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__20080\,
            I => \N__20071\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__20077\,
            I => \N__20068\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__20074\,
            I => \N__20065\
        );

    \I__2575\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20061\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__20068\,
            I => \N__20058\
        );

    \I__2573\ : Span4Mux_h
    port map (
            O => \N__20065\,
            I => \N__20055\
        );

    \I__2572\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20052\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__20061\,
            I => data_out_frame2_11_1
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__20058\,
            I => data_out_frame2_11_1
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__20055\,
            I => data_out_frame2_11_1
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__20052\,
            I => data_out_frame2_11_1
        );

    \I__2567\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__20037\,
            I => \c0.n17288\
        );

    \I__2564\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__20027\
        );

    \I__2562\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20023\
        );

    \I__2561\ : Span4Mux_v
    port map (
            O => \N__20027\,
            I => \N__20020\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__20026\,
            I => \N__20016\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20013\
        );

    \I__2558\ : Sp12to4
    port map (
            O => \N__20020\,
            I => \N__20008\
        );

    \I__2557\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20005\
        );

    \I__2556\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20002\
        );

    \I__2555\ : Span4Mux_s2_h
    port map (
            O => \N__20013\,
            I => \N__19999\
        );

    \I__2554\ : InMux
    port map (
            O => \N__20012\,
            I => \N__19994\
        );

    \I__2553\ : InMux
    port map (
            O => \N__20011\,
            I => \N__19994\
        );

    \I__2552\ : Span12Mux_h
    port map (
            O => \N__20008\,
            I => \N__19989\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__20005\,
            I => \N__19989\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__20002\,
            I => data_out_frame2_12_4
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__19999\,
            I => data_out_frame2_12_4
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__19994\,
            I => data_out_frame2_12_4
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__19989\,
            I => data_out_frame2_12_4
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__19980\,
            I => \c0.n17288_cascade_\
        );

    \I__2545\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__19974\,
            I => \c0.n14_adj_2292\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__19971\,
            I => \N__19967\
        );

    \I__2542\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19964\
        );

    \I__2541\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19961\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__19964\,
            I => \c0.n17294\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__19961\,
            I => \c0.n17294\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__19956\,
            I => \c0.n10428_cascade_\
        );

    \I__2537\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19950\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__19947\,
            I => \N__19944\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__19944\,
            I => \c0.n12_adj_2178\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__2532\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__19929\,
            I => \c0.n10504\
        );

    \I__2528\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__19923\,
            I => \N__19919\
        );

    \I__2526\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19916\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__19919\,
            I => \N__19913\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19908\
        );

    \I__2523\ : Span4Mux_s3_h
    port map (
            O => \N__19913\,
            I => \N__19908\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__19908\,
            I => data_out_frame2_17_1
        );

    \I__2521\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19900\
        );

    \I__2520\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19897\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__19903\,
            I => \N__19894\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19891\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19888\
        );

    \I__2516\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19885\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__19891\,
            I => \N__19881\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__19888\,
            I => \N__19875\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19875\
        );

    \I__2512\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19872\
        );

    \I__2511\ : Span4Mux_s2_h
    port map (
            O => \N__19881\,
            I => \N__19869\
        );

    \I__2510\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19866\
        );

    \I__2509\ : Span4Mux_v
    port map (
            O => \N__19875\,
            I => \N__19863\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19858\
        );

    \I__2507\ : Sp12to4
    port map (
            O => \N__19869\,
            I => \N__19858\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__19866\,
            I => \N__19855\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__19863\,
            I => data_out_frame2_9_4
        );

    \I__2504\ : Odrv12
    port map (
            O => \N__19858\,
            I => data_out_frame2_9_4
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__19855\,
            I => data_out_frame2_9_4
        );

    \I__2502\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19845\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__19839\,
            I => \c0.n17568\
        );

    \I__2498\ : InMux
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__19833\,
            I => \c0.n10554\
        );

    \I__2496\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19826\
        );

    \I__2495\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19823\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__19826\,
            I => \N__19820\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19812\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__19820\,
            I => \N__19812\
        );

    \I__2491\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19809\
        );

    \I__2490\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19806\
        );

    \I__2489\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19803\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__19812\,
            I => \N__19796\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__19809\,
            I => \N__19796\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__19806\,
            I => \N__19796\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__19803\,
            I => data_out_frame2_5_6
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__19796\,
            I => data_out_frame2_5_6
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__19791\,
            I => \c0.n14_adj_2188_cascade_\
        );

    \I__2482\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__19776\,
            I => \c0.n15_adj_2185\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__2476\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__19767\,
            I => \c0.data_out_frame2_20_2\
        );

    \I__2474\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19759\
        );

    \I__2473\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19756\
        );

    \I__2472\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19753\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__19759\,
            I => \N__19749\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__19756\,
            I => \N__19746\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__19753\,
            I => \N__19743\
        );

    \I__2468\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19740\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__19749\,
            I => \N__19737\
        );

    \I__2466\ : Span4Mux_s3_h
    port map (
            O => \N__19746\,
            I => \N__19734\
        );

    \I__2465\ : Span4Mux_s3_h
    port map (
            O => \N__19743\,
            I => \N__19731\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__19740\,
            I => data_out_frame2_7_4
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__19737\,
            I => data_out_frame2_7_4
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__19734\,
            I => data_out_frame2_7_4
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__19731\,
            I => data_out_frame2_7_4
        );

    \I__2460\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__19719\,
            I => \c0.n17240\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__19716\,
            I => \c0.n17240_cascade_\
        );

    \I__2457\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__19710\,
            I => \N__19707\
        );

    \I__2455\ : Span12Mux_v
    port map (
            O => \N__19707\,
            I => \N__19704\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__19704\,
            I => \c0.n14_adj_2206\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__2452\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__19695\,
            I => \N__19692\
        );

    \I__2450\ : Span12Mux_v
    port map (
            O => \N__19692\,
            I => \N__19689\
        );

    \I__2449\ : Odrv12
    port map (
            O => \N__19689\,
            I => \c0.n17439\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__2447\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19680\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__19680\,
            I => \c0.n17249\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__19677\,
            I => \N__19674\
        );

    \I__2444\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19671\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__19671\,
            I => \N__19668\
        );

    \I__2442\ : Span12Mux_v
    port map (
            O => \N__19668\,
            I => \N__19665\
        );

    \I__2441\ : Odrv12
    port map (
            O => \N__19665\,
            I => \c0.data_out_frame2_19_5\
        );

    \I__2440\ : InMux
    port map (
            O => \N__19662\,
            I => \N__19658\
        );

    \I__2439\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19655\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19649\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__19652\,
            I => \N__19646\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__19649\,
            I => \N__19643\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__19646\,
            I => \c0.n17116\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__19643\,
            I => \c0.n17116\
        );

    \I__2432\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__19632\,
            I => \N__19628\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__19631\,
            I => \N__19625\
        );

    \I__2428\ : Span4Mux_h
    port map (
            O => \N__19628\,
            I => \N__19622\
        );

    \I__2427\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19619\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__19622\,
            I => \c0.n17234\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__19619\,
            I => \c0.n17234\
        );

    \I__2424\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19611\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__19611\,
            I => \c0.n15_adj_2291\
        );

    \I__2422\ : InMux
    port map (
            O => \N__19608\,
            I => \c0.rx.n16125\
        );

    \I__2421\ : InMux
    port map (
            O => \N__19605\,
            I => \c0.rx.n16126\
        );

    \I__2420\ : InMux
    port map (
            O => \N__19602\,
            I => \c0.rx.n16127\
        );

    \I__2419\ : InMux
    port map (
            O => \N__19599\,
            I => \c0.rx.n16128\
        );

    \I__2418\ : InMux
    port map (
            O => \N__19596\,
            I => \c0.rx.n16129\
        );

    \I__2417\ : InMux
    port map (
            O => \N__19593\,
            I => \c0.rx.n16130\
        );

    \I__2416\ : InMux
    port map (
            O => \N__19590\,
            I => \c0.rx.n16131\
        );

    \I__2415\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19583\
        );

    \I__2414\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19580\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19577\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__19580\,
            I => \N__19572\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__19577\,
            I => \N__19572\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__19572\,
            I => data_out_frame2_18_1
        );

    \I__2409\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__19566\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_31\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \n5244_cascade_\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__19560\,
            I => \n11018_cascade_\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__19557\,
            I => \N__19538\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__19556\,
            I => \N__19534\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__19555\,
            I => \N__19530\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__19554\,
            I => \N__19526\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__19553\,
            I => \N__19523\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__19552\,
            I => \N__19520\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__19551\,
            I => \N__19516\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__19550\,
            I => \N__19512\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__19549\,
            I => \N__19508\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__19548\,
            I => \N__19503\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__19547\,
            I => \N__19499\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__19546\,
            I => \N__19495\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__19545\,
            I => \N__19491\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__19544\,
            I => \N__19487\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__19543\,
            I => \N__19483\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__19542\,
            I => \N__19479\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__19541\,
            I => \N__19475\
        );

    \I__2388\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19472\
        );

    \I__2387\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19457\
        );

    \I__2386\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19457\
        );

    \I__2385\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19457\
        );

    \I__2384\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19457\
        );

    \I__2383\ : InMux
    port map (
            O => \N__19529\,
            I => \N__19457\
        );

    \I__2382\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19457\
        );

    \I__2381\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19457\
        );

    \I__2380\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19440\
        );

    \I__2379\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19440\
        );

    \I__2378\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19440\
        );

    \I__2377\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19440\
        );

    \I__2376\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19440\
        );

    \I__2375\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19440\
        );

    \I__2374\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19440\
        );

    \I__2373\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19440\
        );

    \I__2372\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19423\
        );

    \I__2371\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19423\
        );

    \I__2370\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19423\
        );

    \I__2369\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19423\
        );

    \I__2368\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19423\
        );

    \I__2367\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19423\
        );

    \I__2366\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19423\
        );

    \I__2365\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19423\
        );

    \I__2364\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19406\
        );

    \I__2363\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19406\
        );

    \I__2362\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19406\
        );

    \I__2361\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19406\
        );

    \I__2360\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19406\
        );

    \I__2359\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19406\
        );

    \I__2358\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19406\
        );

    \I__2357\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19406\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__19472\,
            I => \N__19397\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__19457\,
            I => \N__19397\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__19440\,
            I => \N__19397\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__19423\,
            I => \N__19397\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__19406\,
            I => \c0.n18008\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__19397\,
            I => \c0.n18008\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__19392\,
            I => \n13692_cascade_\
        );

    \I__2349\ : InMux
    port map (
            O => \N__19389\,
            I => \bfn_4_32_0_\
        );

    \I__2348\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19383\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19380\
        );

    \I__2346\ : Span4Mux_s3_h
    port map (
            O => \N__19380\,
            I => \N__19377\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__19377\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_23\
        );

    \I__2344\ : InMux
    port map (
            O => \N__19374\,
            I => \c0.n16101\
        );

    \I__2343\ : InMux
    port map (
            O => \N__19371\,
            I => \bfn_4_30_0_\
        );

    \I__2342\ : InMux
    port map (
            O => \N__19368\,
            I => \c0.n16103\
        );

    \I__2341\ : InMux
    port map (
            O => \N__19365\,
            I => \c0.n16104\
        );

    \I__2340\ : InMux
    port map (
            O => \N__19362\,
            I => \c0.n16105\
        );

    \I__2339\ : InMux
    port map (
            O => \N__19359\,
            I => \N__19356\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__19356\,
            I => \N__19353\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__19353\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_28\
        );

    \I__2336\ : InMux
    port map (
            O => \N__19350\,
            I => \c0.n16106\
        );

    \I__2335\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__19344\,
            I => \N__19341\
        );

    \I__2333\ : Span4Mux_s3_v
    port map (
            O => \N__19341\,
            I => \N__19338\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__19338\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_29\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__19335\,
            I => \N__19332\
        );

    \I__2330\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19323\
        );

    \I__2328\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19316\
        );

    \I__2327\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19316\
        );

    \I__2326\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19316\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__19323\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__19316\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__2323\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19308\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__19308\,
            I => \N__19305\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__19305\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_29\
        );

    \I__2320\ : InMux
    port map (
            O => \N__19302\,
            I => \c0.n16107\
        );

    \I__2319\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19296\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__19296\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_30\
        );

    \I__2317\ : InMux
    port map (
            O => \N__19293\,
            I => \c0.n16108\
        );

    \I__2316\ : InMux
    port map (
            O => \N__19290\,
            I => \c0.n16109\
        );

    \I__2315\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19284\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__19281\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_14\
        );

    \I__2312\ : InMux
    port map (
            O => \N__19278\,
            I => \c0.n16092\
        );

    \I__2311\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19272\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__2309\ : Span4Mux_s3_h
    port map (
            O => \N__19269\,
            I => \N__19266\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__19266\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_15\
        );

    \I__2307\ : InMux
    port map (
            O => \N__19263\,
            I => \c0.n16093\
        );

    \I__2306\ : InMux
    port map (
            O => \N__19260\,
            I => \bfn_4_29_0_\
        );

    \I__2305\ : InMux
    port map (
            O => \N__19257\,
            I => \c0.n16095\
        );

    \I__2304\ : InMux
    port map (
            O => \N__19254\,
            I => \c0.n16096\
        );

    \I__2303\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__19242\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_19\
        );

    \I__2299\ : InMux
    port map (
            O => \N__19239\,
            I => \c0.n16097\
        );

    \I__2298\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__19227\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_20\
        );

    \I__2294\ : InMux
    port map (
            O => \N__19224\,
            I => \c0.n16098\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__19215\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_21\
        );

    \I__2290\ : InMux
    port map (
            O => \N__19212\,
            I => \c0.n16099\
        );

    \I__2289\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__19206\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_22\
        );

    \I__2287\ : InMux
    port map (
            O => \N__19203\,
            I => \c0.n16100\
        );

    \I__2286\ : InMux
    port map (
            O => \N__19200\,
            I => \c0.n16084\
        );

    \I__2285\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__19194\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_7\
        );

    \I__2283\ : InMux
    port map (
            O => \N__19191\,
            I => \c0.n16085\
        );

    \I__2282\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__19182\,
            I => \N__19179\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__19179\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_8\
        );

    \I__2278\ : InMux
    port map (
            O => \N__19176\,
            I => \bfn_4_28_0_\
        );

    \I__2277\ : InMux
    port map (
            O => \N__19173\,
            I => \c0.n16087\
        );

    \I__2276\ : InMux
    port map (
            O => \N__19170\,
            I => \c0.n16088\
        );

    \I__2275\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19164\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__19158\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_11\
        );

    \I__2271\ : InMux
    port map (
            O => \N__19155\,
            I => \c0.n16089\
        );

    \I__2270\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__19149\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_12\
        );

    \I__2268\ : InMux
    port map (
            O => \N__19146\,
            I => \c0.n16090\
        );

    \I__2267\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__19137\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_13\
        );

    \I__2264\ : InMux
    port map (
            O => \N__19134\,
            I => \c0.n16091\
        );

    \I__2263\ : SRMux
    port map (
            O => \N__19131\,
            I => \N__19128\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__19128\,
            I => \N__19125\
        );

    \I__2261\ : Span4Mux_s3_h
    port map (
            O => \N__19125\,
            I => \N__19122\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__19122\,
            I => \c0.n3_adj_2179\
        );

    \I__2259\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19116\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19113\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__19113\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_0\
        );

    \I__2256\ : InMux
    port map (
            O => \N__19110\,
            I => \bfn_4_27_0_\
        );

    \I__2255\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19101\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__19101\,
            I => \N__19098\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__19098\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_1\
        );

    \I__2251\ : InMux
    port map (
            O => \N__19095\,
            I => \c0.n16079\
        );

    \I__2250\ : InMux
    port map (
            O => \N__19092\,
            I => \c0.n16080\
        );

    \I__2249\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19086\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__19086\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_3\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__19083\,
            I => \N__19080\
        );

    \I__2246\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19076\
        );

    \I__2245\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19071\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19068\
        );

    \I__2243\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19063\
        );

    \I__2242\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19063\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__19071\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__19068\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__19063\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__2238\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19053\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__19053\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_3\
        );

    \I__2236\ : InMux
    port map (
            O => \N__19050\,
            I => \c0.n16081\
        );

    \I__2235\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__19044\,
            I => \c0.FRAME_MATCHER_i_31_N_1310_4\
        );

    \I__2233\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19035\
        );

    \I__2232\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19032\
        );

    \I__2231\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19027\
        );

    \I__2230\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19027\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__19024\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__19032\,
            I => \N__19019\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__19027\,
            I => \N__19019\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__19024\,
            I => \N__19016\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__19019\,
            I => \N__19013\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__19016\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__19013\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__2222\ : InMux
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__19005\,
            I => \N__19002\
        );

    \I__2220\ : Span4Mux_s3_h
    port map (
            O => \N__19002\,
            I => \N__18999\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__18999\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_4\
        );

    \I__2218\ : InMux
    port map (
            O => \N__18996\,
            I => \c0.n16082\
        );

    \I__2217\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18990\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__18990\,
            I => \c0.n43\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__2214\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18978\
        );

    \I__2213\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18971\
        );

    \I__2212\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18971\
        );

    \I__2211\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18971\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__18978\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__18971\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__2208\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__18963\,
            I => \c0.FRAME_MATCHER_i_31_N_1278_5\
        );

    \I__2206\ : InMux
    port map (
            O => \N__18960\,
            I => \c0.n16083\
        );

    \I__2205\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18953\
        );

    \I__2204\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18947\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__18953\,
            I => \N__18944\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__18952\,
            I => \N__18941\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__18951\,
            I => \N__18938\
        );

    \I__2200\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18935\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18932\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__18944\,
            I => \N__18929\
        );

    \I__2197\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18926\
        );

    \I__2196\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18923\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__18935\,
            I => data_out_frame2_9_2
        );

    \I__2194\ : Odrv12
    port map (
            O => \N__18932\,
            I => data_out_frame2_9_2
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__18929\,
            I => data_out_frame2_9_2
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__18926\,
            I => data_out_frame2_9_2
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__18923\,
            I => data_out_frame2_9_2
        );

    \I__2190\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18909\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__18909\,
            I => \N__18906\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__18903\,
            I => \c0.n18046\
        );

    \I__2186\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18897\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__18897\,
            I => \N__18894\
        );

    \I__2184\ : Span4Mux_h
    port map (
            O => \N__18894\,
            I => \N__18890\
        );

    \I__2183\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18887\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__18890\,
            I => \c0.n17165\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__18887\,
            I => \c0.n17165\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__18882\,
            I => \N__18879\
        );

    \I__2179\ : InMux
    port map (
            O => \N__18879\,
            I => \N__18876\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__18876\,
            I => \c0.n10334\
        );

    \I__2177\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18870\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__18870\,
            I => \c0.n10223\
        );

    \I__2175\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18864\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__18864\,
            I => \N__18861\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__18861\,
            I => \N__18858\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__18858\,
            I => \c0.n10_adj_2190\
        );

    \I__2171\ : SRMux
    port map (
            O => \N__18855\,
            I => \N__18852\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__18852\,
            I => \N__18849\
        );

    \I__2169\ : Span4Mux_h
    port map (
            O => \N__18849\,
            I => \N__18846\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__18846\,
            I => \c0.n3_adj_2282\
        );

    \I__2167\ : SRMux
    port map (
            O => \N__18843\,
            I => \N__18840\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__18840\,
            I => \c0.n3_adj_2227\
        );

    \I__2165\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18832\
        );

    \I__2164\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18829\
        );

    \I__2163\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18825\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__18832\,
            I => \N__18822\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__18829\,
            I => \N__18819\
        );

    \I__2160\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18815\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__18825\,
            I => \N__18812\
        );

    \I__2158\ : Span4Mux_s3_h
    port map (
            O => \N__18822\,
            I => \N__18809\
        );

    \I__2157\ : Span4Mux_s3_h
    port map (
            O => \N__18819\,
            I => \N__18806\
        );

    \I__2156\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18803\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__18815\,
            I => data_out_frame2_7_6
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__18812\,
            I => data_out_frame2_7_6
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__18809\,
            I => data_out_frame2_7_6
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__18806\,
            I => data_out_frame2_7_6
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__18803\,
            I => data_out_frame2_7_6
        );

    \I__2150\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18788\
        );

    \I__2149\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18784\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__18788\,
            I => \N__18781\
        );

    \I__2147\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18777\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__18784\,
            I => \N__18774\
        );

    \I__2145\ : Span4Mux_h
    port map (
            O => \N__18781\,
            I => \N__18771\
        );

    \I__2144\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18768\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__18777\,
            I => data_out_frame2_6_4
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__18774\,
            I => data_out_frame2_6_4
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__18771\,
            I => data_out_frame2_6_4
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__18768\,
            I => data_out_frame2_6_4
        );

    \I__2139\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18756\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__18756\,
            I => \c0.n6_adj_2339\
        );

    \I__2137\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18750\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__18747\,
            I => \N__18744\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__18744\,
            I => \N__18740\
        );

    \I__2133\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18737\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__18740\,
            I => \c0.n10507\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__18737\,
            I => \c0.n10507\
        );

    \I__2130\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18727\
        );

    \I__2129\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18723\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__18730\,
            I => \N__18719\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__18727\,
            I => \N__18716\
        );

    \I__2126\ : InMux
    port map (
            O => \N__18726\,
            I => \N__18713\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__18723\,
            I => \N__18709\
        );

    \I__2124\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18706\
        );

    \I__2123\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18703\
        );

    \I__2122\ : Span4Mux_s2_h
    port map (
            O => \N__18716\,
            I => \N__18700\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18697\
        );

    \I__2120\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18694\
        );

    \I__2119\ : Span4Mux_h
    port map (
            O => \N__18709\,
            I => \N__18691\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18682\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__18703\,
            I => \N__18682\
        );

    \I__2116\ : Sp12to4
    port map (
            O => \N__18700\,
            I => \N__18682\
        );

    \I__2115\ : Sp12to4
    port map (
            O => \N__18697\,
            I => \N__18682\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__18694\,
            I => data_out_frame2_15_0
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__18691\,
            I => data_out_frame2_15_0
        );

    \I__2112\ : Odrv12
    port map (
            O => \N__18682\,
            I => data_out_frame2_15_0
        );

    \I__2111\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__18672\,
            I => \N__18669\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__18669\,
            I => \c0.n17273\
        );

    \I__2108\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18661\
        );

    \I__2107\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18658\
        );

    \I__2106\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18655\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__18661\,
            I => \N__18650\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__18658\,
            I => \N__18650\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18646\
        );

    \I__2102\ : Sp12to4
    port map (
            O => \N__18650\,
            I => \N__18643\
        );

    \I__2101\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18640\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__18646\,
            I => \N__18637\
        );

    \I__2099\ : Span12Mux_v
    port map (
            O => \N__18643\,
            I => \N__18634\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__18640\,
            I => data_out_frame2_6_7
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__18637\,
            I => data_out_frame2_6_7
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__18634\,
            I => data_out_frame2_6_7
        );

    \I__2095\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18623\
        );

    \I__2094\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18620\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__18623\,
            I => \N__18614\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__18620\,
            I => \N__18611\
        );

    \I__2091\ : InMux
    port map (
            O => \N__18619\,
            I => \N__18606\
        );

    \I__2090\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18606\
        );

    \I__2089\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18603\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__18614\,
            I => \N__18598\
        );

    \I__2087\ : Span4Mux_s3_h
    port map (
            O => \N__18611\,
            I => \N__18598\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18595\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__18603\,
            I => data_out_frame2_16_1
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__18598\,
            I => data_out_frame2_16_1
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__18595\,
            I => data_out_frame2_16_1
        );

    \I__2082\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18585\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__18582\,
            I => \c0.n17153\
        );

    \I__2079\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18576\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__18576\,
            I => \c0.n17168\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__18573\,
            I => \c0.n17153_cascade_\
        );

    \I__2076\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18567\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__18567\,
            I => \c0.n26_adj_2203\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__18564\,
            I => \N__18561\
        );

    \I__2073\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18557\
        );

    \I__2072\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18553\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18550\
        );

    \I__2070\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18547\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18542\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__18550\,
            I => \N__18542\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18539\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18534\
        );

    \I__2065\ : Span4Mux_s3_h
    port map (
            O => \N__18539\,
            I => \N__18531\
        );

    \I__2064\ : InMux
    port map (
            O => \N__18538\,
            I => \N__18526\
        );

    \I__2063\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18526\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__18534\,
            I => data_out_frame2_5_7
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__18531\,
            I => data_out_frame2_5_7
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__18526\,
            I => data_out_frame2_5_7
        );

    \I__2059\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18513\
        );

    \I__2058\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18510\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__18517\,
            I => \N__18507\
        );

    \I__2056\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18504\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__18513\,
            I => \N__18501\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__18510\,
            I => \N__18498\
        );

    \I__2053\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18495\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__18504\,
            I => data_out_frame2_13_3
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__18501\,
            I => data_out_frame2_13_3
        );

    \I__2050\ : Odrv12
    port map (
            O => \N__18498\,
            I => data_out_frame2_13_3
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__18495\,
            I => data_out_frame2_13_3
        );

    \I__2048\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18483\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__18483\,
            I => \N__18479\
        );

    \I__2046\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18476\
        );

    \I__2045\ : Span12Mux_s3_h
    port map (
            O => \N__18479\,
            I => \N__18473\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__18476\,
            I => data_out_frame2_18_4
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__18473\,
            I => data_out_frame2_18_4
        );

    \I__2042\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18465\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__18465\,
            I => \N__18460\
        );

    \I__2040\ : InMux
    port map (
            O => \N__18464\,
            I => \N__18457\
        );

    \I__2039\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18454\
        );

    \I__2038\ : Span4Mux_s2_h
    port map (
            O => \N__18460\,
            I => \N__18450\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__18457\,
            I => \N__18447\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__18454\,
            I => \N__18444\
        );

    \I__2035\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18441\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__18450\,
            I => \N__18436\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__18447\,
            I => \N__18436\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__18444\,
            I => \N__18433\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__18441\,
            I => data_out_frame2_5_5
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__18436\,
            I => data_out_frame2_5_5
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__18433\,
            I => data_out_frame2_5_5
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__18426\,
            I => \N__18422\
        );

    \I__2027\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18418\
        );

    \I__2026\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18415\
        );

    \I__2025\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18412\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__18418\,
            I => \N__18408\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__18415\,
            I => \N__18405\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__18412\,
            I => \N__18402\
        );

    \I__2021\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18399\
        );

    \I__2020\ : Span4Mux_s3_h
    port map (
            O => \N__18408\,
            I => \N__18396\
        );

    \I__2019\ : Span4Mux_s3_h
    port map (
            O => \N__18405\,
            I => \N__18391\
        );

    \I__2018\ : Span4Mux_s3_h
    port map (
            O => \N__18402\,
            I => \N__18391\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__18399\,
            I => data_out_frame2_7_3
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__18396\,
            I => data_out_frame2_7_3
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__18391\,
            I => data_out_frame2_7_3
        );

    \I__2014\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18378\
        );

    \I__2012\ : Sp12to4
    port map (
            O => \N__18378\,
            I => \N__18374\
        );

    \I__2011\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__2010\ : Span12Mux_v
    port map (
            O => \N__18374\,
            I => \N__18368\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__18371\,
            I => data_out_frame2_17_4
        );

    \I__2008\ : Odrv12
    port map (
            O => \N__18368\,
            I => data_out_frame2_17_4
        );

    \I__2007\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__18360\,
            I => \N__18356\
        );

    \I__2005\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__18356\,
            I => \N__18350\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__18353\,
            I => data_out_frame2_17_7
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__18350\,
            I => data_out_frame2_17_7
        );

    \I__2001\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18339\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__18339\,
            I => \N__18336\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__18336\,
            I => \c0.n10356\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__1996\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18327\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18324\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__18324\,
            I => \N__18320\
        );

    \I__1993\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18317\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__18320\,
            I => \c0.n10572\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__18317\,
            I => \c0.n10572\
        );

    \I__1990\ : InMux
    port map (
            O => \N__18312\,
            I => \N__18309\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__18309\,
            I => \N__18306\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__18306\,
            I => \c0.n16_adj_2170\
        );

    \I__1987\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18300\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__18300\,
            I => \N__18296\
        );

    \I__1985\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18292\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__18296\,
            I => \N__18289\
        );

    \I__1983\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18285\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__18292\,
            I => \N__18280\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__18289\,
            I => \N__18280\
        );

    \I__1980\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18277\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__18285\,
            I => data_out_frame2_6_5
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__18280\,
            I => data_out_frame2_6_5
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__18277\,
            I => data_out_frame2_6_5
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__18270\,
            I => \c0.n16_adj_2320_cascade_\
        );

    \I__1975\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18264\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__18264\,
            I => \N__18261\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__18261\,
            I => \N__18257\
        );

    \I__1972\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18254\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__18257\,
            I => \c0.n17216\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__18254\,
            I => \c0.n17216\
        );

    \I__1969\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18246\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__18243\,
            I => \c0.data_out_frame2_19_1\
        );

    \I__1966\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18237\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__18237\,
            I => \c0.n18058\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__18234\,
            I => \c0.n6_adj_2175_cascade_\
        );

    \I__1963\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18227\
        );

    \I__1962\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18224\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18221\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__18224\,
            I => \N__18218\
        );

    \I__1959\ : Span4Mux_s3_h
    port map (
            O => \N__18221\,
            I => \N__18215\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__18218\,
            I => \c0.n17258\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__18215\,
            I => \c0.n17258\
        );

    \I__1956\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18207\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__18207\,
            I => \N__18203\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__18206\,
            I => \N__18198\
        );

    \I__1953\ : Span4Mux_s3_h
    port map (
            O => \N__18203\,
            I => \N__18194\
        );

    \I__1952\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18189\
        );

    \I__1951\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18189\
        );

    \I__1950\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18184\
        );

    \I__1949\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18184\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__18194\,
            I => data_out_frame2_11_2
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__18189\,
            I => data_out_frame2_11_2
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__18184\,
            I => data_out_frame2_11_2
        );

    \I__1945\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18173\
        );

    \I__1944\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18170\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18165\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18165\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__18165\,
            I => \N__18162\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__18162\,
            I => \c0.n17171\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__18159\,
            I => \N__18156\
        );

    \I__1938\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18153\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__18153\,
            I => \N__18150\
        );

    \I__1936\ : Span4Mux_h
    port map (
            O => \N__18150\,
            I => \N__18147\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__18147\,
            I => \c0.n17132\
        );

    \I__1934\ : InMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__18141\,
            I => \N__18137\
        );

    \I__1932\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18134\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__18137\,
            I => \N__18131\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18128\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__18131\,
            I => \c0.n17184\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__18128\,
            I => \c0.n17184\
        );

    \I__1927\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__18120\,
            I => \c0.n32\
        );

    \I__1925\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__1922\ : Span4Mux_s1_h
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__18105\,
            I => \c0.n10437\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__18102\,
            I => \c0.n17249_cascade_\
        );

    \I__1919\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18096\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__18096\,
            I => \N__18093\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__18090\,
            I => \c0.n12_adj_2298\
        );

    \I__1915\ : InMux
    port map (
            O => \N__18087\,
            I => \N__18081\
        );

    \I__1914\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18077\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__18085\,
            I => \N__18074\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__18084\,
            I => \N__18071\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__18081\,
            I => \N__18068\
        );

    \I__1910\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18065\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__18077\,
            I => \N__18062\
        );

    \I__1908\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18058\
        );

    \I__1907\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18055\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__18068\,
            I => \N__18052\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__18065\,
            I => \N__18049\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__18062\,
            I => \N__18046\
        );

    \I__1903\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18043\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__18058\,
            I => data_out_frame2_8_1
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__18055\,
            I => data_out_frame2_8_1
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__18052\,
            I => data_out_frame2_8_1
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__18049\,
            I => data_out_frame2_8_1
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__18046\,
            I => data_out_frame2_8_1
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__18043\,
            I => data_out_frame2_8_1
        );

    \I__1896\ : InMux
    port map (
            O => \N__18030\,
            I => \N__18027\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__18027\,
            I => \N__18024\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__18024\,
            I => \N__18021\
        );

    \I__1893\ : Span4Mux_s0_h
    port map (
            O => \N__18021\,
            I => \N__18018\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__18018\,
            I => \c0.n20\
        );

    \I__1891\ : InMux
    port map (
            O => \N__18015\,
            I => \N__18012\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__18012\,
            I => \N__18009\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__18009\,
            I => \N__18006\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__18006\,
            I => \N__18003\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__18003\,
            I => \c0.n17678\
        );

    \I__1886\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17996\
        );

    \I__1885\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17993\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__17996\,
            I => \N__17990\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17987\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__17990\,
            I => \N__17984\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__17987\,
            I => \N__17981\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__17984\,
            I => \N__17978\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__17981\,
            I => \c0.n17279\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__17978\,
            I => \c0.n17279\
        );

    \I__1877\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17970\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__1875\ : Sp12to4
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__1874\ : Odrv12
    port map (
            O => \N__17964\,
            I => \c0.data_out_frame2_20_1\
        );

    \I__1873\ : InMux
    port map (
            O => \N__17961\,
            I => \N__17953\
        );

    \I__1872\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17953\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__17959\,
            I => \N__17950\
        );

    \I__1870\ : InMux
    port map (
            O => \N__17958\,
            I => \N__17947\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__17953\,
            I => \N__17944\
        );

    \I__1868\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17941\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__17947\,
            I => \N__17935\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__17944\,
            I => \N__17935\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__17941\,
            I => \N__17932\
        );

    \I__1864\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17929\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__17935\,
            I => \N__17926\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__17932\,
            I => \N__17923\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__17929\,
            I => data_out_frame2_13_0
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__17926\,
            I => data_out_frame2_13_0
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__17923\,
            I => data_out_frame2_13_0
        );

    \I__1858\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17913\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__17913\,
            I => \N__17910\
        );

    \I__1856\ : Span4Mux_h
    port map (
            O => \N__17910\,
            I => \N__17906\
        );

    \I__1855\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17903\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__17906\,
            I => \c0.n10424\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__17903\,
            I => \c0.n10424\
        );

    \I__1852\ : InMux
    port map (
            O => \N__17898\,
            I => \N__17895\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__17895\,
            I => \N__17892\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__17892\,
            I => \N__17889\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__17889\,
            I => \c0.n14_adj_2346\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__17886\,
            I => \c0.n15_adj_2341_cascade_\
        );

    \I__1847\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17879\
        );

    \I__1846\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17876\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__17879\,
            I => \N__17870\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__17876\,
            I => \N__17870\
        );

    \I__1843\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17866\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__17870\,
            I => \N__17863\
        );

    \I__1841\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17860\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__17866\,
            I => data_out_frame2_14_5
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__17863\,
            I => data_out_frame2_14_5
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__17860\,
            I => data_out_frame2_14_5
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__17853\,
            I => \c0.n18178_cascade_\
        );

    \I__1836\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17847\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17844\
        );

    \I__1834\ : Span4Mux_h
    port map (
            O => \N__17844\,
            I => \N__17841\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__17838\,
            I => \c0.n6_adj_2161\
        );

    \I__1831\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17832\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__17832\,
            I => \c0.n18181\
        );

    \I__1829\ : InMux
    port map (
            O => \N__17829\,
            I => \N__17825\
        );

    \I__1828\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17822\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__17825\,
            I => \N__17819\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17814\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__17819\,
            I => \N__17811\
        );

    \I__1824\ : InMux
    port map (
            O => \N__17818\,
            I => \N__17806\
        );

    \I__1823\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17806\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__17814\,
            I => data_out_frame2_16_6
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__17811\,
            I => data_out_frame2_16_6
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__17806\,
            I => data_out_frame2_16_6
        );

    \I__1819\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__17796\,
            I => \c0.n18112\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \N__17789\
        );

    \I__1816\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17784\
        );

    \I__1815\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17784\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__17784\,
            I => data_out_frame2_17_6
        );

    \I__1813\ : InMux
    port map (
            O => \N__17781\,
            I => \N__17778\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__17778\,
            I => \N__17775\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__17775\,
            I => \N__17772\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__17772\,
            I => \c0.data_out_frame2_20_6\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__17769\,
            I => \c0.n18115_cascade_\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__17766\,
            I => \N__17763\
        );

    \I__1807\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17760\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__17760\,
            I => \c0.n22_adj_2364\
        );

    \I__1805\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17753\
        );

    \I__1804\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17750\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__17753\,
            I => data_out_frame2_18_6
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__17750\,
            I => data_out_frame2_18_6
        );

    \I__1801\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17742\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__17742\,
            I => \c0.n18031\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__17739\,
            I => \N__17736\
        );

    \I__1798\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17733\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__17733\,
            I => \N__17730\
        );

    \I__1796\ : Span4Mux_s3_h
    port map (
            O => \N__17730\,
            I => \N__17727\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__17727\,
            I => \c0.n10548\
        );

    \I__1794\ : SRMux
    port map (
            O => \N__17724\,
            I => \N__17721\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__17721\,
            I => \c0.n3_adj_2278\
        );

    \I__1792\ : SRMux
    port map (
            O => \N__17718\,
            I => \N__17715\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__17715\,
            I => \N__17712\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__17712\,
            I => \c0.n3_adj_2266\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__17709\,
            I => \N__17706\
        );

    \I__1788\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17703\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__17703\,
            I => \N__17700\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__17700\,
            I => \N__17697\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__17697\,
            I => \c0.data_out_frame2_19_6\
        );

    \I__1784\ : IoInMux
    port map (
            O => \N__17694\,
            I => \N__17691\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__17691\,
            I => \N__17688\
        );

    \I__1782\ : Span4Mux_s2_h
    port map (
            O => \N__17688\,
            I => \N__17685\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__17685\,
            I => tx2_enable
        );

    \I__1780\ : SRMux
    port map (
            O => \N__17682\,
            I => \N__17679\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__17679\,
            I => \N__17676\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__17676\,
            I => \c0.n3_adj_2232\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__17673\,
            I => \N__17667\
        );

    \I__1776\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17664\
        );

    \I__1775\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17660\
        );

    \I__1774\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17657\
        );

    \I__1773\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17654\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__17664\,
            I => \N__17651\
        );

    \I__1771\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17648\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__17660\,
            I => \N__17645\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17640\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__17654\,
            I => \N__17640\
        );

    \I__1767\ : Span4Mux_h
    port map (
            O => \N__17651\,
            I => \N__17637\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__17648\,
            I => data_out_frame2_9_1
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__17645\,
            I => data_out_frame2_9_1
        );

    \I__1764\ : Odrv12
    port map (
            O => \N__17640\,
            I => data_out_frame2_9_1
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__17637\,
            I => data_out_frame2_9_1
        );

    \I__1762\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17625\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17621\
        );

    \I__1760\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17618\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__17621\,
            I => \c0.n10346\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__17618\,
            I => \c0.n10346\
        );

    \I__1757\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17610\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__17610\,
            I => \N__17606\
        );

    \I__1755\ : InMux
    port map (
            O => \N__17609\,
            I => \N__17603\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__17606\,
            I => \c0.n17231\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__17603\,
            I => \c0.n17231\
        );

    \I__1752\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17595\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__17595\,
            I => \N__17592\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__17592\,
            I => \c0.n18076\
        );

    \I__1749\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17584\
        );

    \I__1748\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17581\
        );

    \I__1747\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17578\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__17584\,
            I => \N__17571\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__17581\,
            I => \N__17571\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17568\
        );

    \I__1743\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17563\
        );

    \I__1742\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17563\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__17571\,
            I => data_out_frame2_9_5
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__17568\,
            I => data_out_frame2_9_5
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__17563\,
            I => data_out_frame2_9_5
        );

    \I__1738\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17553\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__17553\,
            I => \N__17550\
        );

    \I__1736\ : Span4Mux_s2_h
    port map (
            O => \N__17550\,
            I => \N__17547\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__17547\,
            I => \N__17544\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__17544\,
            I => \c0.n18109\
        );

    \I__1733\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17537\
        );

    \I__1732\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17534\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17530\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__17534\,
            I => \N__17526\
        );

    \I__1729\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17523\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__17530\,
            I => \N__17520\
        );

    \I__1727\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17517\
        );

    \I__1726\ : Span4Mux_s1_h
    port map (
            O => \N__17526\,
            I => \N__17514\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__17523\,
            I => data_out_frame2_6_3
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__17520\,
            I => data_out_frame2_6_3
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__17517\,
            I => data_out_frame2_6_3
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__17514\,
            I => data_out_frame2_6_3
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__17505\,
            I => \c0.n10334_cascade_\
        );

    \I__1720\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17498\
        );

    \I__1719\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__17498\,
            I => \c0.n10533\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__17495\,
            I => \c0.n10533\
        );

    \I__1716\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17487\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__17487\,
            I => \c0.n10_adj_2297\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__17484\,
            I => \c0.n14_adj_2296_cascade_\
        );

    \I__1713\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17478\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__17478\,
            I => \N__17474\
        );

    \I__1711\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17471\
        );

    \I__1710\ : Sp12to4
    port map (
            O => \N__17474\,
            I => \N__17468\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__17471\,
            I => \N__17465\
        );

    \I__1708\ : Odrv12
    port map (
            O => \N__17468\,
            I => \c0.n17267\
        );

    \I__1707\ : Odrv12
    port map (
            O => \N__17465\,
            I => \c0.n17267\
        );

    \I__1706\ : InMux
    port map (
            O => \N__17460\,
            I => \N__17457\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__17457\,
            I => \N__17453\
        );

    \I__1704\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17450\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__17453\,
            I => \N__17447\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17444\
        );

    \I__1701\ : Span4Mux_v
    port map (
            O => \N__17447\,
            I => \N__17438\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__17444\,
            I => \N__17435\
        );

    \I__1699\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17428\
        );

    \I__1698\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17428\
        );

    \I__1697\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17428\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__17438\,
            I => data_out_frame2_13_2
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__17435\,
            I => data_out_frame2_13_2
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__17428\,
            I => data_out_frame2_13_2
        );

    \I__1693\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17418\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__17418\,
            I => \N__17415\
        );

    \I__1691\ : Span4Mux_s2_h
    port map (
            O => \N__17415\,
            I => \N__17411\
        );

    \I__1690\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17408\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__17411\,
            I => \c0.n17309\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__17408\,
            I => \c0.n17309\
        );

    \I__1687\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17399\
        );

    \I__1686\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17396\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__17399\,
            I => \N__17393\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__17396\,
            I => \c0.n17291\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__17393\,
            I => \c0.n17291\
        );

    \I__1682\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17385\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__17385\,
            I => \N__17382\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__17382\,
            I => \N__17378\
        );

    \I__1679\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17375\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__17378\,
            I => \c0.n17303\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__17375\,
            I => \c0.n17303\
        );

    \I__1676\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17367\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__17367\,
            I => \c0.n25\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__17364\,
            I => \c0.n28_adj_2200_cascade_\
        );

    \I__1673\ : InMux
    port map (
            O => \N__17361\,
            I => \N__17358\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__17358\,
            I => \c0.n27_adj_2204\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__17355\,
            I => \c0.n10223_cascade_\
        );

    \I__1670\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17349\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__17349\,
            I => \c0.n6_adj_2318\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__17346\,
            I => \N__17343\
        );

    \I__1667\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17340\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17337\
        );

    \I__1665\ : Span4Mux_s2_h
    port map (
            O => \N__17337\,
            I => \N__17334\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__17334\,
            I => \c0.n17569\
        );

    \I__1663\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17324\
        );

    \I__1661\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17321\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__17324\,
            I => \N__17318\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__17321\,
            I => data_out_frame2_17_5
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__17318\,
            I => data_out_frame2_17_5
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__17313\,
            I => \N__17309\
        );

    \I__1656\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17306\
        );

    \I__1655\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17303\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__17306\,
            I => \N__17298\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__17303\,
            I => \N__17298\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__17298\,
            I => \c0.n17138\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__17295\,
            I => \c0.n6_adj_2228_cascade_\
        );

    \I__1650\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17289\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__1648\ : Span4Mux_s3_h
    port map (
            O => \N__17286\,
            I => \N__17282\
        );

    \I__1647\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17279\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__17282\,
            I => \c0.n17312\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__17279\,
            I => \c0.n17312\
        );

    \I__1644\ : InMux
    port map (
            O => \N__17274\,
            I => \N__17266\
        );

    \I__1643\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17266\
        );

    \I__1642\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17262\
        );

    \I__1641\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17259\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__17266\,
            I => \N__17256\
        );

    \I__1639\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17253\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__17262\,
            I => \N__17250\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__17259\,
            I => data_out_frame2_14_3
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__17256\,
            I => data_out_frame2_14_3
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__17253\,
            I => data_out_frame2_14_3
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__17250\,
            I => data_out_frame2_14_3
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__17241\,
            I => \c0.n33_cascade_\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__17238\,
            I => \N__17235\
        );

    \I__1631\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17232\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__17232\,
            I => \N__17229\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__17229\,
            I => \c0.data_out_frame2_19_7\
        );

    \I__1628\ : InMux
    port map (
            O => \N__17226\,
            I => \N__17223\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__17223\,
            I => \c0.n30_adj_2218\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__17220\,
            I => \c0.n17300_cascade_\
        );

    \I__1625\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17214\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__17214\,
            I => \c0.n34\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__17211\,
            I => \N__17208\
        );

    \I__1622\ : InMux
    port map (
            O => \N__17208\,
            I => \N__17205\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__17205\,
            I => \N__17202\
        );

    \I__1620\ : Odrv12
    port map (
            O => \N__17202\,
            I => \c0.n17237\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__17199\,
            I => \N__17196\
        );

    \I__1618\ : InMux
    port map (
            O => \N__17196\,
            I => \N__17193\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__17193\,
            I => \N__17190\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__17190\,
            I => \N__17187\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__17187\,
            I => \c0.n10440\
        );

    \I__1614\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17181\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__17181\,
            I => \c0.n6_adj_2215\
        );

    \I__1612\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17175\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__17175\,
            I => \c0.n17219\
        );

    \I__1610\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17169\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__17169\,
            I => \N__17166\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__17166\,
            I => \c0.n17141\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__17163\,
            I => \c0.n17219_cascade_\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__17160\,
            I => \c0.n17_cascade_\
        );

    \I__1605\ : InMux
    port map (
            O => \N__17157\,
            I => \N__17153\
        );

    \I__1604\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17150\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__17153\,
            I => \N__17147\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__17150\,
            I => \N__17144\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__17147\,
            I => \c0.n17228\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__17144\,
            I => \c0.n17228\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__17139\,
            I => \c0.n17246_cascade_\
        );

    \I__1598\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17133\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__17133\,
            I => \N__17130\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__17130\,
            I => \N__17127\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__17127\,
            I => \c0.n17187\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__17124\,
            I => \c0.n18238_cascade_\
        );

    \I__1593\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17118\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__17118\,
            I => \c0.n18241\
        );

    \I__1591\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17112\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__17112\,
            I => \N__17109\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__17109\,
            I => \N__17106\
        );

    \I__1588\ : Span4Mux_v
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__1587\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17097\
        );

    \I__1586\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17092\
        );

    \I__1585\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17092\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__17100\,
            I => data_out_frame2_7_7
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__17097\,
            I => data_out_frame2_7_7
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__17092\,
            I => data_out_frame2_7_7
        );

    \I__1581\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17082\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__17082\,
            I => \N__17079\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__17079\,
            I => \c0.n5_adj_2137\
        );

    \I__1578\ : InMux
    port map (
            O => \N__17076\,
            I => \N__17073\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__17073\,
            I => \c0.n18154\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__17070\,
            I => \c0.n18130_cascade_\
        );

    \I__1575\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17064\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__17064\,
            I => \N__17061\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__17061\,
            I => \N__17058\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__17058\,
            I => \N__17055\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__17055\,
            I => \c0.data_out_frame2_20_7\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__17052\,
            I => \c0.n18133_cascade_\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__17049\,
            I => \N__17046\
        );

    \I__1568\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17043\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__17043\,
            I => \N__17040\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__17040\,
            I => \c0.n22_adj_2363\
        );

    \I__1565\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17034\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__17034\,
            I => \N__17031\
        );

    \I__1563\ : Span4Mux_h
    port map (
            O => \N__17031\,
            I => \N__17028\
        );

    \I__1562\ : Span4Mux_s1_h
    port map (
            O => \N__17028\,
            I => \N__17025\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__17025\,
            I => \N__17022\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__17022\,
            I => \c0.n18028\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__17019\,
            I => \c0.n18040_cascade_\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__17016\,
            I => \c0.n18010_cascade_\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__17013\,
            I => \c0.n18013_cascade_\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__17010\,
            I => \N__17007\
        );

    \I__1555\ : InMux
    port map (
            O => \N__17007\,
            I => \N__17004\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__17004\,
            I => \c0.n22_adj_2375\
        );

    \I__1553\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16998\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__16998\,
            I => \N__16995\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__16995\,
            I => \c0.n18025\
        );

    \I__1550\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16989\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16986\
        );

    \I__1548\ : Odrv12
    port map (
            O => \N__16986\,
            I => \c0.n10530\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__16983\,
            I => \c0.n10530_cascade_\
        );

    \I__1546\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16976\
        );

    \I__1545\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16973\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__16976\,
            I => \N__16970\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__16973\,
            I => \N__16967\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__16970\,
            I => \c0.n10371\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__16967\,
            I => \c0.n10371\
        );

    \I__1540\ : InMux
    port map (
            O => \N__16962\,
            I => \N__16956\
        );

    \I__1539\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16953\
        );

    \I__1538\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16948\
        );

    \I__1537\ : InMux
    port map (
            O => \N__16959\,
            I => \N__16948\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__16956\,
            I => \N__16945\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__16953\,
            I => data_out_frame2_7_0
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__16948\,
            I => data_out_frame2_7_0
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__16945\,
            I => data_out_frame2_7_0
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__16938\,
            I => \N__16934\
        );

    \I__1531\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16927\
        );

    \I__1530\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16927\
        );

    \I__1529\ : InMux
    port map (
            O => \N__16933\,
            I => \N__16922\
        );

    \I__1528\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16922\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__16927\,
            I => \N__16919\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__16922\,
            I => data_out_frame2_6_0
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__16919\,
            I => data_out_frame2_6_0
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__16914\,
            I => \N__16911\
        );

    \I__1523\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16908\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__16908\,
            I => \N__16905\
        );

    \I__1521\ : Span4Mux_s1_h
    port map (
            O => \N__16905\,
            I => \N__16902\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__16902\,
            I => \c0.n5_adj_2343\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__16899\,
            I => \N__16895\
        );

    \I__1518\ : InMux
    port map (
            O => \N__16898\,
            I => \N__16892\
        );

    \I__1517\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16887\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__16892\,
            I => \N__16884\
        );

    \I__1515\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16881\
        );

    \I__1514\ : InMux
    port map (
            O => \N__16890\,
            I => \N__16878\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__16887\,
            I => \N__16871\
        );

    \I__1512\ : Span4Mux_v
    port map (
            O => \N__16884\,
            I => \N__16871\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__16881\,
            I => \N__16871\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__16878\,
            I => data_out_frame2_15_5
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__16871\,
            I => data_out_frame2_15_5
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__16866\,
            I => \c0.n18100_cascade_\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__16863\,
            I => \N__16860\
        );

    \I__1506\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16857\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__16857\,
            I => \N__16854\
        );

    \I__1504\ : Span12Mux_s1_h
    port map (
            O => \N__16854\,
            I => \N__16851\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__16851\,
            I => \c0.n18103\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__16848\,
            I => \c0.n10520_cascade_\
        );

    \I__1501\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16842\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__16842\,
            I => \N__16838\
        );

    \I__1499\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16835\
        );

    \I__1498\ : Odrv12
    port map (
            O => \N__16838\,
            I => \c0.n10349\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__16835\,
            I => \c0.n10349\
        );

    \I__1496\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16827\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__16827\,
            I => \N__16824\
        );

    \I__1494\ : Odrv12
    port map (
            O => \N__16824\,
            I => \c0.n10462\
        );

    \I__1493\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16818\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__16818\,
            I => \N__16815\
        );

    \I__1491\ : Odrv12
    port map (
            O => \N__16815\,
            I => \c0.n15_adj_2312\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__16812\,
            I => \N__16808\
        );

    \I__1489\ : InMux
    port map (
            O => \N__16811\,
            I => \N__16805\
        );

    \I__1488\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16802\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16799\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__16802\,
            I => \N__16796\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__16799\,
            I => \c0.n17285\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__16796\,
            I => \c0.n17285\
        );

    \I__1483\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16788\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__16788\,
            I => \c0.n18136\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__16785\,
            I => \N__16782\
        );

    \I__1480\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16779\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__16779\,
            I => \N__16776\
        );

    \I__1478\ : Span4Mux_v
    port map (
            O => \N__16776\,
            I => \N__16773\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__16773\,
            I => \c0.data_out_frame2_19_2\
        );

    \I__1476\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16767\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__16767\,
            I => \c0.n17135\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__16764\,
            I => \c0.n17092_cascade_\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__16761\,
            I => \c0.n17_adj_2294_cascade_\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__16758\,
            I => \N__16755\
        );

    \I__1471\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16752\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__16752\,
            I => \N__16749\
        );

    \I__1469\ : Odrv12
    port map (
            O => \N__16749\,
            I => \c0.data_out_frame2_19_4\
        );

    \I__1468\ : InMux
    port map (
            O => \N__16746\,
            I => \N__16743\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__16743\,
            I => \c0.n12\
        );

    \I__1466\ : InMux
    port map (
            O => \N__16740\,
            I => \N__16735\
        );

    \I__1465\ : InMux
    port map (
            O => \N__16739\,
            I => \N__16730\
        );

    \I__1464\ : InMux
    port map (
            O => \N__16738\,
            I => \N__16730\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__16735\,
            I => \N__16727\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__16730\,
            I => data_out_frame2_14_0
        );

    \I__1461\ : Odrv12
    port map (
            O => \N__16727\,
            I => data_out_frame2_14_0
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__16722\,
            I => \c0.n17237_cascade_\
        );

    \I__1459\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16716\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__16716\,
            I => \c0.n16_adj_2293\
        );

    \I__1457\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16710\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__16710\,
            I => \N__16707\
        );

    \I__1455\ : Span4Mux_h
    port map (
            O => \N__16707\,
            I => \N__16704\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__16704\,
            I => \c0.data_out_frame2_20_4\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__16701\,
            I => \c0.n18277_cascade_\
        );

    \I__1452\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16695\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__16695\,
            I => \c0.n22_adj_2367\
        );

    \I__1450\ : InMux
    port map (
            O => \N__16692\,
            I => \N__16689\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__16689\,
            I => \c0.n18034\
        );

    \I__1448\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16683\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__16683\,
            I => \N__16679\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__16682\,
            I => \N__16676\
        );

    \I__1445\ : Span4Mux_h
    port map (
            O => \N__16679\,
            I => \N__16673\
        );

    \I__1444\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16670\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__16673\,
            I => \c0.n17225\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__16670\,
            I => \c0.n17225\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__16665\,
            I => \c0.n17135_cascade_\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__16662\,
            I => \c0.n21_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16656\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__16656\,
            I => \c0.n20_adj_2223\
        );

    \I__1437\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16650\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__16650\,
            I => \c0.n19_adj_2224\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__16647\,
            I => \c0.n14_adj_2308_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16641\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__16641\,
            I => \c0.n18022\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__16638\,
            I => \c0.n5_adj_2353_cascade_\
        );

    \I__1431\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16632\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__16632\,
            I => \N__16629\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__16629\,
            I => \c0.n6\
        );

    \I__1428\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16623\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__16623\,
            I => \N__16620\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__16620\,
            I => \c0.n6_adj_2138\
        );

    \I__1425\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16614\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__16614\,
            I => \N__16611\
        );

    \I__1423\ : Span4Mux_h
    port map (
            O => \N__16611\,
            I => \N__16608\
        );

    \I__1422\ : Span4Mux_v
    port map (
            O => \N__16608\,
            I => \N__16605\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__16605\,
            I => \c0.n17440\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__16602\,
            I => \c0.n18037_cascade_\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__16599\,
            I => \c0.n18274_cascade_\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__16596\,
            I => \c0.n5_adj_2315_cascade_\
        );

    \I__1417\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16586\
        );

    \I__1416\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16586\
        );

    \I__1415\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16583\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__16586\,
            I => data_out_frame2_13_7
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__16583\,
            I => data_out_frame2_13_7
        );

    \I__1412\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16574\
        );

    \I__1411\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16571\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__16574\,
            I => \N__16568\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__16571\,
            I => data_out_frame2_18_5
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__16568\,
            I => data_out_frame2_18_5
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__16563\,
            I => \c0.n24_cascade_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16557\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__16557\,
            I => \c0.n22\
        );

    \I__1404\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__16551\,
            I => \c0.n17174\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__16548\,
            I => \c0.n17174_cascade_\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__16545\,
            I => \c0.n10356_cascade_\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__16542\,
            I => \N__16539\
        );

    \I__1399\ : InMux
    port map (
            O => \N__16539\,
            I => \N__16536\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__16536\,
            I => \N__16533\
        );

    \I__1397\ : Odrv12
    port map (
            O => \N__16533\,
            I => \c0.n18139\
        );

    \I__1396\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16527\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__16527\,
            I => \N__16524\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__16524\,
            I => \c0.n14\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__16521\,
            I => \c0.n15_cascade_\
        );

    \I__1392\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16515\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__16515\,
            I => \c0.data_out_frame2_20_5\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__16512\,
            I => \c0.n17306_cascade_\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__16509\,
            I => \c0.n18094_cascade_\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__16506\,
            I => \c0.n18097_cascade_\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__16503\,
            I => \c0.n18262_cascade_\
        );

    \I__1386\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16497\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__16497\,
            I => \c0.n22_adj_2365\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__16494\,
            I => \c0.n18265_cascade_\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__16491\,
            I => \c0.n10468_cascade_\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__16488\,
            I => \c0.n17610_cascade_\
        );

    \I__1381\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16482\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__16482\,
            I => \c0.n18214\
        );

    \I__1379\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16476\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__16476\,
            I => \c0.n18217\
        );

    \I__1377\ : IoInMux
    port map (
            O => \N__16473\,
            I => \N__16470\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__16470\,
            I => \N__16467\
        );

    \I__1375\ : IoSpan4Mux
    port map (
            O => \N__16467\,
            I => \N__16464\
        );

    \I__1374\ : IoSpan4Mux
    port map (
            O => \N__16464\,
            I => \N__16461\
        );

    \I__1373\ : IoSpan4Mux
    port map (
            O => \N__16461\,
            I => \N__16458\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__16458\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_10_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16017,
            carryinitout => \bfn_10_26_0_\
        );

    \IN_MUX_bfv_10_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16025,
            carryinitout => \bfn_10_27_0_\
        );

    \IN_MUX_bfv_10_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16033,
            carryinitout => \bfn_10_28_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_5_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15986,
            carryinitout => \bfn_5_24_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n15994,
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16002,
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_24_0_\
        );

    \IN_MUX_bfv_6_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n16139\,
            carryinitout => \bfn_6_25_0_\
        );

    \IN_MUX_bfv_16_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_28_0_\
        );

    \IN_MUX_bfv_16_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n16124\,
            carryinitout => \bfn_16_29_0_\
        );

    \IN_MUX_bfv_4_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_32_0_\
        );

    \IN_MUX_bfv_12_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_31_0_\
        );

    \IN_MUX_bfv_12_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16073\,
            carryinitout => \bfn_12_32_0_\
        );

    \IN_MUX_bfv_4_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_27_0_\
        );

    \IN_MUX_bfv_4_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16086\,
            carryinitout => \bfn_4_28_0_\
        );

    \IN_MUX_bfv_4_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16094\,
            carryinitout => \bfn_4_29_0_\
        );

    \IN_MUX_bfv_4_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n16102\,
            carryinitout => \bfn_4_30_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_14_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_30_0_\
        );

    \IN_MUX_bfv_9_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_29_0_\
        );

    \IN_MUX_bfv_9_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16048,
            carryinitout => \bfn_9_30_0_\
        );

    \IN_MUX_bfv_9_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16056,
            carryinitout => \bfn_9_31_0_\
        );

    \IN_MUX_bfv_9_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n16064,
            carryinitout => \bfn_9_32_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16473\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_695_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24937\,
            in1 => \N__17460\,
            in2 => \_gnd_net_\,
            in3 => \N__18732\,
            lcout => \c0.n10440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18022_bdd_4_lut_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__28699\,
            in1 => \N__16644\,
            in2 => \N__17673\,
            in3 => \N__18086\,
            lcout => \c0.n18025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15153_3_lut_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__34724\,
            in1 => \N__28969\,
            in2 => \_gnd_net_\,
            in3 => \N__28700\,
            lcout => OPEN,
            ltout => \c0.n17610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18214_bdd_4_lut_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__16626\,
            in1 => \N__16485\,
            in2 => \N__16488\,
            in3 => \N__32463\,
            lcout => \c0.n18217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15410_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23412\,
            in1 => \N__32458\,
            in2 => \N__16542\,
            in3 => \N__32171\,
            lcout => \c0.n18214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__16479\,
            in1 => \N__32459\,
            in2 => \N__17049\,
            in3 => \N__32289\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49627\,
            ce => \N__24272\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15306_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__28652\,
            in1 => \N__16578\,
            in2 => \N__19677\,
            in3 => \N__29048\,
            lcout => OPEN,
            ltout => \c0.n18094_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18094_bdd_4_lut_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__17331\,
            in1 => \N__28653\,
            in2 => \N__16509\,
            in3 => \N__20561\,
            lcout => OPEN,
            ltout => \c0.n18097_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32172\,
            in1 => \N__16518\,
            in2 => \N__16506\,
            in3 => \N__21210\,
            lcout => \c0.n22_adj_2365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__17556\,
            in1 => \N__32460\,
            in2 => \N__16863\,
            in3 => \N__32173\,
            lcout => OPEN,
            ltout => \c0.n18262_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18262_bdd_4_lut_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32461\,
            in1 => \N__18015\,
            in2 => \N__16503\,
            in3 => \N__16635\,
            lcout => OPEN,
            ltout => \c0.n18265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__16500\,
            in1 => \N__32462\,
            in2 => \N__16494\,
            in3 => \N__32287\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49628\,
            ce => \N__24269\,
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_747_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37582\,
            in1 => \N__37637\,
            in2 => \N__18426\,
            in3 => \N__17274\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_477_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17670\,
            in2 => \_gnd_net_\,
            in3 => \N__18626\,
            lcout => OPEN,
            ltout => \c0.n10468_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_430_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24396\,
            in1 => \N__18140\,
            in2 => \N__16491\,
            in3 => \N__16845\,
            lcout => OPEN,
            ltout => \c0.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i166_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16530\,
            in1 => \N__24705\,
            in2 => \N__16521\,
            in3 => \N__20145\,
            lcout => \c0.data_out_frame2_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49631\,
            ce => \N__26610\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_431_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37581\,
            lcout => OPEN,
            ltout => \c0.n17306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i165_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24942\,
            in1 => \N__16746\,
            in2 => \N__16512\,
            in3 => \N__21870\,
            lcout => \c0.data_out_frame2_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49631\,
            ce => \N__26610\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_599_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23150\,
            lcout => \c0.n10437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15288_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__28684\,
            in1 => \N__29006\,
            in2 => \N__20396\,
            in3 => \N__24032\,
            lcout => \c0.n18064\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_721_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26054\,
            in1 => \N__24528\,
            in2 => \N__20439\,
            in3 => \N__20562\,
            lcout => \c0.n17225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18425\,
            in1 => \N__29007\,
            in2 => \_gnd_net_\,
            in3 => \N__17529\,
            lcout => \c0.n5_adj_2337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i105_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17940\,
            in1 => \N__30921\,
            in2 => \_gnd_net_\,
            in3 => \N__26589\,
            lcout => data_out_frame2_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i74_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26588\,
            in1 => \N__30843\,
            in2 => \_gnd_net_\,
            in3 => \N__17663\,
            lcout => data_out_frame2_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_586_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23303\,
            lcout => \c0.n17187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i150_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26587\,
            in1 => \N__30054\,
            in2 => \_gnd_net_\,
            in3 => \N__16577\,
            lcout => data_out_frame2_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__29008\,
            in1 => \N__19819\,
            in2 => \N__16914\,
            in3 => \N__28685\,
            lcout => \c0.n6_adj_2161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_422_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24653\,
            in1 => \N__37203\,
            in2 => \N__16899\,
            in3 => \N__16560\,
            lcout => OPEN,
            ltout => \c0.n24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i168_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18030\,
            in1 => \N__19638\,
            in2 => \N__16563\,
            in3 => \N__16811\,
            lcout => \c0.data_out_frame2_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49641\,
            ce => \N__26611\,
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17312\,
            in1 => \N__16554\,
            in2 => \N__16682\,
            in3 => \N__23453\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_648_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20087\,
            in1 => \N__18210\,
            in2 => \_gnd_net_\,
            in3 => \N__21828\,
            lcout => \c0.n17174\,
            ltout => \c0.n17174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_494_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19763\,
            in1 => \N__20525\,
            in2 => \N__16548\,
            in3 => \N__24327\,
            lcout => \c0.n10356\,
            ltout => \c0.n10356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_496_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18463\,
            in2 => \N__16545\,
            in3 => \N__24652\,
            lcout => \c0.n17184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18136_bdd_4_lut_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__16592\,
            in1 => \N__28694\,
            in2 => \N__20438\,
            in3 => \N__16791\,
            lcout => \c0.n18139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i126_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30599\,
            in1 => \N__16890\,
            in2 => \_gnd_net_\,
            in3 => \N__26597\,
            lcout => data_out_frame2_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i47_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31458\,
            in1 => \N__19817\,
            in2 => \_gnd_net_\,
            in3 => \N__26598\,
            lcout => data_out_frame2_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19762\,
            in1 => \N__29058\,
            in2 => \_gnd_net_\,
            in3 => \N__18792\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14663_4_lut_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__29059\,
            in1 => \N__28695\,
            in2 => \N__16596\,
            in3 => \N__21795\,
            lcout => \c0.n17440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_564_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23820\,
            in2 => \_gnd_net_\,
            in3 => \N__18080\,
            lcout => \c0.n17132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i112_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31400\,
            in1 => \N__16593\,
            in2 => \_gnd_net_\,
            in3 => \N__26596\,
            lcout => data_out_frame2_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i64_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30466\,
            in1 => \N__17104\,
            in2 => \_gnd_net_\,
            in3 => \N__26600\,
            lcout => data_out_frame2_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_478_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16591\,
            in1 => \N__17540\,
            in2 => \_gnd_net_\,
            in3 => \N__24482\,
            lcout => \c0.n17285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i78_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17577\,
            in1 => \N__31514\,
            in2 => \_gnd_net_\,
            in3 => \N__26601\,
            lcout => data_out_frame2_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_683_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17103\,
            in1 => \N__23296\,
            in2 => \N__23449\,
            in3 => \N__17576\,
            lcout => \c0.n10349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i128_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30465\,
            in1 => \N__24582\,
            in2 => \_gnd_net_\,
            in3 => \N__26599\,
            lcout => data_out_frame2_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i15_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19275\,
            in2 => \_gnd_net_\,
            in3 => \N__33220\,
            lcout => \c0.FRAME_MATCHER_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49661\,
            ce => 'H',
            sr => \N__20856\
        );

    \c0.FRAME_MATCHER_i_i20_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19236\,
            in2 => \_gnd_net_\,
            in3 => \N__33247\,
            lcout => \c0.FRAME_MATCHER_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49669\,
            ce => 'H',
            sr => \N__20757\
        );

    \c0.FRAME_MATCHER_i_i8_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19188\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33148\,
            lcout => \c0.FRAME_MATCHER_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49681\,
            ce => 'H',
            sr => \N__20907\
        );

    \c0.FRAME_MATCHER_i_i14_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19287\,
            in2 => \_gnd_net_\,
            in3 => \N__33149\,
            lcout => \c0.FRAME_MATCHER_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49692\,
            ce => 'H',
            sr => \N__27957\
        );

    \c0.FRAME_MATCHER_i_i4_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19008\,
            in2 => \_gnd_net_\,
            in3 => \N__33150\,
            lcout => \c0.FRAME_MATCHER_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49703\,
            ce => 'H',
            sr => \N__19131\
        );

    \c0.FRAME_MATCHER_i_i11_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19167\,
            in2 => \_gnd_net_\,
            in3 => \N__33151\,
            lcout => \c0.FRAME_MATCHER_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49717\,
            ce => 'H',
            sr => \N__20841\
        );

    \c0.FRAME_MATCHER_i_i23_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19386\,
            in2 => \_gnd_net_\,
            in3 => \N__33152\,
            lcout => \c0.FRAME_MATCHER_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49728\,
            ce => 'H',
            sr => \N__20967\
        );

    \c0.data_out_5__0__2216_LC_1_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__48166\,
            in1 => \N__30873\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_6__1__N_537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49738\,
            ce => \N__50589\,
            sr => \N__42807\
        );

    \c0.data_out_5__7__2209_LC_1_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48165\,
            in2 => \_gnd_net_\,
            in3 => \N__31344\,
            lcout => \c0.data_out_7__3__N_441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49738\,
            ce => \N__50589\,
            sr => \N__42807\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15356_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__28961\,
            in1 => \N__18726\,
            in2 => \N__28675\,
            in3 => \N__16740\,
            lcout => \c0.n18154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15250_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21572\,
            in1 => \N__28631\,
            in2 => \N__20088\,
            in3 => \N__28962\,
            lcout => \c0.n18022\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28967\,
            in1 => \N__18303\,
            in2 => \_gnd_net_\,
            in3 => \N__21958\,
            lcout => OPEN,
            ltout => \c0.n5_adj_2353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__18468\,
            in1 => \N__28638\,
            in2 => \N__16638\,
            in3 => \N__28968\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__17085\,
            in1 => \N__28637\,
            in2 => \N__18564\,
            in3 => \N__28966\,
            lcout => \c0.n6_adj_2138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18034_bdd_4_lut_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__32442\,
            in1 => \N__16617\,
            in2 => \N__19701\,
            in3 => \N__16692\,
            lcout => OPEN,
            ltout => \c0.n18037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__16698\,
            in1 => \N__32443\,
            in2 => \N__16602\,
            in3 => \N__32288\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49629\,
            ce => \N__24270\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18486\,
            in1 => \N__28639\,
            in2 => \N__16758\,
            in3 => \N__29047\,
            lcout => OPEN,
            ltout => \c0.n18274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18274_bdd_4_lut_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__28640\,
            in1 => \N__18384\,
            in2 => \N__16599\,
            in3 => \N__20123\,
            lcout => OPEN,
            ltout => \c0.n18277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32175\,
            in1 => \N__16713\,
            in2 => \N__16701\,
            in3 => \N__21212\,
            lcout => \c0.n22_adj_2367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15371_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__19848\,
            in1 => \N__32441\,
            in2 => \N__17346\,
            in3 => \N__32174\,
            lcout => \c0.n18034\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_667_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23389\,
            in1 => \N__23190\,
            in2 => \N__20187\,
            in3 => \N__20030\,
            lcout => \c0.n17135\,
            ltout => \c0.n17135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_521_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18000\,
            in1 => \N__16686\,
            in2 => \N__16665\,
            in3 => \N__17421\,
            lcout => OPEN,
            ltout => \c0.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i159_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16659\,
            in2 => \N__16662\,
            in3 => \N__16653\,
            lcout => \c0.data_out_frame2_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49632\,
            ce => \N__26564\,
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_518_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24105\,
            in1 => \N__24381\,
            in2 => \N__19941\,
            in3 => \N__20208\,
            lcout => \c0.n20_adj_2223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_520_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17671\,
            in1 => \N__16992\,
            in2 => \N__17739\,
            in3 => \N__23859\,
            lcout => \c0.n19_adj_2224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_571_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23207\,
            in1 => \N__21665\,
            in2 => \_gnd_net_\,
            in3 => \N__16980\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i155_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17481\,
            in1 => \N__21537\,
            in2 => \N__16647\,
            in3 => \N__16821\,
            lcout => \c0.data_out_frame2_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49636\,
            ce => \N__26608\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_538_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21525\,
            in2 => \_gnd_net_\,
            in3 => \N__23917\,
            lcout => OPEN,
            ltout => \c0.n17092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_535_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17156\,
            in1 => \N__16770\,
            in2 => \N__16764\,
            in3 => \N__41156\,
            lcout => OPEN,
            ltout => \c0.n17_adj_2294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i157_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23208\,
            in1 => \N__17292\,
            in2 => \N__16761\,
            in3 => \N__16719\,
            lcout => \c0.data_out_frame2_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49636\,
            ce => \N__26608\,
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23694\,
            in1 => \N__17402\,
            in2 => \N__20026\,
            in3 => \N__18231\,
            lcout => \c0.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i113_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30413\,
            in1 => \N__16739\,
            in2 => \_gnd_net_\,
            in3 => \N__26555\,
            lcout => data_out_frame2_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i52_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26554\,
            in1 => \N__31209\,
            in2 => \_gnd_net_\,
            in3 => \N__17533\,
            lcout => data_out_frame2_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_608_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17817\,
            in1 => \N__23024\,
            in2 => \_gnd_net_\,
            in3 => \N__16738\,
            lcout => \c0.n17237\,
            ltout => \c0.n17237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_456_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24098\,
            in1 => \N__16959\,
            in2 => \N__16722\,
            in3 => \N__18957\,
            lcout => \c0.n17165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i135_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17818\,
            in1 => \N__29993\,
            in2 => \_gnd_net_\,
            in3 => \N__26556\,
            lcout => data_out_frame2_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_534_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18753\,
            in1 => \N__24782\,
            in2 => \N__23151\,
            in3 => \N__16960\,
            lcout => \c0.n16_adj_2293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i66_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__30278\,
            in1 => \_gnd_net_\,
            in2 => \N__18085\,
            in3 => \N__26557\,
            lcout => data_out_frame2_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15341_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__24583\,
            in1 => \N__22095\,
            in2 => \N__28683\,
            in3 => \N__29024\,
            lcout => \c0.n18136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_650_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18791\,
            in1 => \N__24852\,
            in2 => \N__21369\,
            in3 => \N__20241\,
            lcout => \c0.n17228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15259_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__28655\,
            in1 => \N__20580\,
            in2 => \N__16785\,
            in3 => \N__29023\,
            lcout => \c0.n18028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_685_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23815\,
            in1 => \N__18061\,
            in2 => \_gnd_net_\,
            in3 => \N__21467\,
            lcout => \c0.n10371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_553_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21364\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20240\,
            lcout => \c0.n10462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i57_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29874\,
            in1 => \N__16961\,
            in2 => \_gnd_net_\,
            in3 => \N__26538\,
            lcout => data_out_frame2_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18556\,
            in1 => \N__18835\,
            in2 => \_gnd_net_\,
            in3 => \N__17588\,
            lcout => \c0.n17138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i116_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31208\,
            in1 => \N__17271\,
            in2 => \_gnd_net_\,
            in3 => \N__26561\,
            lcout => data_out_frame2_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_614_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19880\,
            in1 => \N__21457\,
            in2 => \N__16938\,
            in3 => \N__17105\,
            lcout => \c0.n10424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_530_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23725\,
            in2 => \_gnd_net_\,
            in3 => \N__21753\,
            lcout => OPEN,
            ltout => \c0.n10520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_484_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18664\,
            in1 => \N__23396\,
            in2 => \N__16848\,
            in3 => \N__16937\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_592_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17352\,
            in1 => \N__16841\,
            in2 => \N__20397\,
            in3 => \N__21824\,
            lcout => \c0.n17216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_524_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20124\,
            lcout => \c0.n10572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_578_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17502\,
            in1 => \N__24879\,
            in2 => \N__40842\,
            in3 => \N__16830\,
            lcout => \c0.n15_adj_2312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_483_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27595\,
            in1 => \N__17609\,
            in2 => \N__16812\,
            in3 => \N__18260\,
            lcout => \c0.n27_adj_2204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_492_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17909\,
            in1 => \N__18421\,
            in2 => \N__18952\,
            in3 => \N__18837\,
            lcout => \c0.n10_adj_2207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i80_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31392\,
            in1 => \N__23448\,
            in2 => \_gnd_net_\,
            in3 => \N__26562\,
            lcout => data_out_frame2_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_476_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23960\,
            in2 => \_gnd_net_\,
            in3 => \N__21956\,
            lcout => \c0.n10346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_516_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16891\,
            in2 => \_gnd_net_\,
            in3 => \N__22921\,
            lcout => \c0.n10530\,
            ltout => \c0.n10530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_692_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19818\,
            in1 => \N__19905\,
            in2 => \N__16983\,
            in3 => \N__16979\,
            lcout => \c0.n17303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16962\,
            in1 => \N__16932\,
            in2 => \_gnd_net_\,
            in3 => \N__29050\,
            lcout => \c0.n5_adj_2217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i49_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16933\,
            in1 => \N__30405\,
            in2 => \_gnd_net_\,
            in3 => \N__26563\,
            lcout => data_out_frame2_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29049\,
            in1 => \N__40892\,
            in2 => \_gnd_net_\,
            in3 => \N__18836\,
            lcout => \c0.n5_adj_2343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15311_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__28659\,
            in1 => \N__16898\,
            in2 => \N__29073\,
            in3 => \N__17869\,
            lcout => OPEN,
            ltout => \c0.n18100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18100_bdd_4_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__20166\,
            in1 => \N__23723\,
            in2 => \N__16866\,
            in3 => \N__28660\,
            lcout => \c0.n18103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i28_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41556\,
            in2 => \_gnd_net_\,
            in3 => \N__35200\,
            lcout => \c0.FRAME_MATCHER_state_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49682\,
            ce => 'H',
            sr => \N__33600\
        );

    \c0.FRAME_MATCHER_i_i19_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19251\,
            in2 => \_gnd_net_\,
            in3 => \N__33221\,
            lcout => \c0.FRAME_MATCHER_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49693\,
            ce => 'H',
            sr => \N__20826\
        );

    \c0.FRAME_MATCHER_i_i13_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19143\,
            lcout => \c0.FRAME_MATCHER_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49704\,
            ce => 'H',
            sr => \N__17718\
        );

    \c0.FRAME_MATCHER_i_i1_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19107\,
            in2 => \_gnd_net_\,
            in3 => \N__33225\,
            lcout => \c0.FRAME_MATCHER_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49718\,
            ce => 'H',
            sr => \N__25392\
        );

    \c0.FRAME_MATCHER_i_i28_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19359\,
            in2 => \_gnd_net_\,
            in3 => \N__33252\,
            lcout => \c0.FRAME_MATCHER_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49729\,
            ce => 'H',
            sr => \N__22464\
        );

    \c0.FRAME_MATCHER_state_i16_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45036\,
            in1 => \N__44817\,
            in2 => \N__37793\,
            in3 => \N__44611\,
            lcout => \c0.FRAME_MATCHER_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49739\,
            ce => 'H',
            sr => \N__33582\
        );

    \c0.data_out_7__3__2197_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__48426\,
            in1 => \N__50337\,
            in2 => \N__31995\,
            in3 => \N__46476\,
            lcout => \c0.data_out_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49750\,
            ce => \N__46935\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__17121\,
            in1 => \N__32424\,
            in2 => \N__17010\,
            in3 => \N__32275\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49633\,
            ce => \N__24273\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15240_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__29057\,
            in1 => \N__18249\,
            in2 => \N__28676\,
            in3 => \N__19587\,
            lcout => OPEN,
            ltout => \c0.n18010_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18010_bdd_4_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__19926\,
            in1 => \N__18627\,
            in2 => \N__17016\,
            in3 => \N__28636\,
            lcout => OPEN,
            ltout => \c0.n18013_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__21199\,
            in1 => \N__32153\,
            in2 => \N__17013\,
            in3 => \N__17973\,
            lcout => \c0.n22_adj_2375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15425_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__17001\,
            in1 => \N__32446\,
            in2 => \N__32170\,
            in3 => \N__23577\,
            lcout => OPEN,
            ltout => \c0.n18238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18238_bdd_4_lut_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32447\,
            in1 => \N__23061\,
            in2 => \N__17124\,
            in3 => \N__23349\,
            lcout => \c0.n18241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18665\,
            in1 => \_gnd_net_\,
            in2 => \N__29022\,
            in3 => \N__17115\,
            lcout => \c0.n5_adj_2137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18154_bdd_4_lut_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__17076\,
            in1 => \N__26053\,
            in2 => \N__17959\,
            in3 => \N__28632\,
            lcout => \c0.n18157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15336_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__28549\,
            in1 => \N__22005\,
            in2 => \N__17238\,
            in3 => \N__29056\,
            lcout => OPEN,
            ltout => \c0.n18130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18130_bdd_4_lut_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__18363\,
            in1 => \N__27655\,
            in2 => \N__17070\,
            in3 => \N__28550\,
            lcout => OPEN,
            ltout => \c0.n18133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17067\,
            in1 => \N__21203\,
            in2 => \N__17052\,
            in3 => \N__32169\,
            lcout => \c0.n22_adj_2363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18028_bdd_4_lut_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__28548\,
            in1 => \N__17037\,
            in2 => \N__21984\,
            in3 => \N__20339\,
            lcout => \c0.n18031\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15264_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__28546\,
            in1 => \N__21666\,
            in2 => \N__20625\,
            in3 => \N__29055\,
            lcout => OPEN,
            ltout => \c0.n18040_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18040_bdd_4_lut_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__17456\,
            in1 => \N__23916\,
            in2 => \N__17019\,
            in3 => \N__28547\,
            lcout => \c0.n18043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_502_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17184\,
            in1 => \N__40273\,
            in2 => \N__23046\,
            in3 => \N__17178\,
            lcout => \c0.n10263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_500_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37587\,
            in2 => \_gnd_net_\,
            in3 => \N__40103\,
            lcout => \c0.n6_adj_2215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_525_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17882\,
            in2 => \_gnd_net_\,
            in3 => \N__23259\,
            lcout => \c0.n17141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_499_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34326\,
            lcout => \c0.n17219\,
            ltout => \c0.n17219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18956\,
            in1 => \N__17172\,
            in2 => \N__17163\,
            in3 => \N__20340\,
            lcout => OPEN,
            ltout => \c0.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i167_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18312\,
            in1 => \N__24698\,
            in2 => \N__17160\,
            in3 => \N__17388\,
            lcout => \c0.data_out_frame2_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49637\,
            ce => \N__26609\,
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_505_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18560\,
            in1 => \N__23654\,
            in2 => \N__40680\,
            in3 => \N__22937\,
            lcout => \c0.n30_adj_2218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_503_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20284\,
            in2 => \_gnd_net_\,
            in3 => \N__17958\,
            lcout => OPEN,
            ltout => \c0.n17246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_508_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17157\,
            in1 => \N__17477\,
            in2 => \N__17139\,
            in3 => \N__17136\,
            lcout => OPEN,
            ltout => \c0.n33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i160_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17217\,
            in1 => \N__23676\,
            in2 => \N__17241\,
            in3 => \N__18123\,
            lcout => \c0.data_out_frame2_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49643\,
            ce => \N__26607\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_504_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23019\,
            in2 => \_gnd_net_\,
            in3 => \N__21957\,
            lcout => OPEN,
            ltout => \c0.n17300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_507_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17226\,
            in1 => \N__19829\,
            in2 => \N__17220\,
            in3 => \N__23186\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_664_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20332\,
            in1 => \N__24426\,
            in2 => \_gnd_net_\,
            in3 => \N__20619\,
            lcout => \c0.n17291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15269_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__29004\,
            in1 => \N__20230\,
            in2 => \N__28654\,
            in3 => \N__18201\,
            lcout => \c0.n18046\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18202\,
            in1 => \N__24498\,
            in2 => \N__17211\,
            in3 => \N__21820\,
            lcout => \c0.n14_adj_2346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15279_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__29005\,
            in1 => \N__17272\,
            in2 => \N__24433\,
            in3 => \N__28596\,
            lcout => \c0.n18058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_450_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18893\,
            in1 => \N__20460\,
            in2 => \N__17199\,
            in3 => \N__17628\,
            lcout => \c0.n15_adj_2185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i101_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30110\,
            in1 => \N__20012\,
            in2 => \_gnd_net_\,
            in3 => \N__26459\,
            lcout => data_out_frame2_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18076_bdd_4_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__20011\,
            in1 => \N__28589\,
            in2 => \N__41157\,
            in3 => \N__17598\,
            lcout => \c0.n17569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i142_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30598\,
            in1 => \N__17327\,
            in2 => \_gnd_net_\,
            in3 => \N__26460\,
            lcout => data_out_frame2_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_438_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18230\,
            in1 => \N__24551\,
            in2 => \N__17313\,
            in3 => \N__17613\,
            lcout => \c0.n12_adj_2178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_706_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23484\,
            in1 => \N__24483\,
            in2 => \_gnd_net_\,
            in3 => \N__24434\,
            lcout => \c0.n17312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_527_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24367\,
            in2 => \_gnd_net_\,
            in3 => \N__18299\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_528_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24176\,
            in1 => \N__18323\,
            in2 => \N__17295\,
            in3 => \N__17285\,
            lcout => \c0.n17116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_513_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__24748\,
            in1 => \N__22973\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_722_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40863\,
            in1 => \N__21300\,
            in2 => \N__40934\,
            in3 => \N__20517\,
            lcout => \c0.n17309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_545_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18177\,
            in1 => \N__17265\,
            in2 => \N__18084\,
            in3 => \N__40929\,
            lcout => \c0.n12_adj_2298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_682_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26052\,
            in1 => \N__23239\,
            in2 => \_gnd_net_\,
            in3 => \N__21573\,
            lcout => \c0.n17194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_684_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17442\,
            in1 => \N__24905\,
            in2 => \N__18730\,
            in3 => \N__17828\,
            lcout => \c0.n17267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_549_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17441\,
            lcout => \c0.n17168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i107_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17443\,
            in1 => \N__31675\,
            in2 => \_gnd_net_\,
            in3 => \N__26583\,
            lcout => data_out_frame2_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_481_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17414\,
            in1 => \N__17403\,
            in2 => \N__41055\,
            in3 => \N__17381\,
            lcout => OPEN,
            ltout => \c0.n28_adj_2200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17370\,
            in1 => \N__18570\,
            in2 => \N__17364\,
            in3 => \N__17361\,
            lcout => \c0.n10223\,
            ltout => \c0.n10223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_729_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18722\,
            in1 => \N__18464\,
            in2 => \N__17355\,
            in3 => \N__23666\,
            lcout => \c0.n14_adj_2206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_591_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18288\,
            in2 => \_gnd_net_\,
            in3 => \N__20557\,
            lcout => \c0.n6_adj_2318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i75_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26580\,
            in1 => \N__31676\,
            in2 => \_gnd_net_\,
            in3 => \N__18950\,
            lcout => data_out_frame2_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i111_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31453\,
            in1 => \N__22927\,
            in2 => \_gnd_net_\,
            in3 => \N__26581\,
            lcout => data_out_frame2_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_556_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18619\,
            in2 => \_gnd_net_\,
            in3 => \N__23958\,
            lcout => \c0.n10533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_734_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18618\,
            in1 => \N__17672\,
            in2 => \N__18517\,
            in3 => \N__17624\,
            lcout => \c0.n17231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15301_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__24783\,
            in1 => \N__28662\,
            in2 => \N__20526\,
            in3 => \N__29054\,
            lcout => \c0.n18076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18106_bdd_4_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__28663\,
            in1 => \N__20352\,
            in2 => \N__40938\,
            in3 => \N__17587\,
            lcout => \c0.n18109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27648\,
            in1 => \N__24079\,
            in2 => \_gnd_net_\,
            in3 => \N__27596\,
            lcout => \c0.n10_adj_2297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i118_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31089\,
            in1 => \N__17875\,
            in2 => \_gnd_net_\,
            in3 => \N__26582\,
            lcout => data_out_frame2_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_699_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21522\,
            in1 => \N__23903\,
            in2 => \_gnd_net_\,
            in3 => \N__20019\,
            lcout => \c0.n10334\,
            ltout => \c0.n10334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_542_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18743\,
            in1 => \N__17541\,
            in2 => \N__17505\,
            in3 => \N__17501\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_544_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18519\,
            in1 => \N__17490\,
            in2 => \N__17484\,
            in3 => \N__23447\,
            lcout => \c0.n17171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i121_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26559\,
            in1 => \N__29872\,
            in2 => \_gnd_net_\,
            in3 => \N__18712\,
            lcout => data_out_frame2_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i102_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30049\,
            in1 => \N__20167\,
            in2 => \_gnd_net_\,
            in3 => \N__26560\,
            lcout => data_out_frame2_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i110_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26558\,
            in1 => \N__31506\,
            in2 => \_gnd_net_\,
            in3 => \N__23724\,
            lcout => data_out_frame2_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i3_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19056\,
            in2 => \_gnd_net_\,
            in3 => \N__33246\,
            lcout => \c0.FRAME_MATCHER_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49694\,
            ce => 'H',
            sr => \N__18843\
        );

    \c0.FRAME_MATCHER_i_i7_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19197\,
            in2 => \_gnd_net_\,
            in3 => \N__33219\,
            lcout => \c0.FRAME_MATCHER_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49705\,
            ce => 'H',
            sr => \N__17724\
        );

    \c0.i18_4_lut_adj_674_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27081\,
            in1 => \N__25867\,
            in2 => \N__27206\,
            in3 => \N__19326\,
            lcout => \c0.n43_adj_2380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i29_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19311\,
            in2 => \_gnd_net_\,
            in3 => \N__33222\,
            lcout => \c0.FRAME_MATCHER_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49719\,
            ce => 'H',
            sr => \N__17682\
        );

    \c0.select_219_Select_29_i3_2_lut_3_lut_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41906\,
            in1 => \N__27840\,
            in2 => \_gnd_net_\,
            in3 => \N__19328\,
            lcout => \c0.n3_adj_2232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10659_2_lut_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19327\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41903\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_7_i3_2_lut_3_lut_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27842\,
            in1 => \N__27082\,
            in2 => \_gnd_net_\,
            in3 => \N__41907\,
            lcout => \c0.n3_adj_2278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_13_i3_2_lut_3_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__41905\,
            in1 => \N__27198\,
            in2 => \_gnd_net_\,
            in3 => \N__27841\,
            lcout => \c0.n3_adj_2266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10676_2_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41904\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i22_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19209\,
            in2 => \_gnd_net_\,
            in3 => \N__33224\,
            lcout => \c0.FRAME_MATCHER_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49730\,
            ce => 'H',
            sr => \N__25362\
        );

    \c0.FRAME_MATCHER_i_i31_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19569\,
            in2 => \_gnd_net_\,
            in3 => \N__33251\,
            lcout => \c0.FRAME_MATCHER_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49740\,
            ce => 'H',
            sr => \N__22344\
        );

    \c0.FRAME_MATCHER_i_i30_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19299\,
            in2 => \_gnd_net_\,
            in3 => \N__33248\,
            lcout => \c0.FRAME_MATCHER_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49751\,
            ce => 'H',
            sr => \N__22452\
        );

    \c0.FRAME_MATCHER_i_i21_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19221\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33249\,
            lcout => \c0.FRAME_MATCHER_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49763\,
            ce => 'H',
            sr => \N__20769\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15321_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__28970\,
            in1 => \N__17756\,
            in2 => \N__17709\,
            in3 => \N__28598\,
            lcout => \c0.n18112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__17835\,
            in1 => \N__32423\,
            in2 => \N__17766\,
            in3 => \N__32261\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49638\,
            ce => \N__24271\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i143_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30533\,
            in1 => \N__17792\,
            in2 => \_gnd_net_\,
            in3 => \N__26545\,
            lcout => data_out_frame2_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15400_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21429\,
            in1 => \N__32444\,
            in2 => \N__22905\,
            in3 => \N__32147\,
            lcout => OPEN,
            ltout => \c0.n18178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18178_bdd_4_lut_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32445\,
            in1 => \N__22806\,
            in2 => \N__17853\,
            in3 => \N__17850\,
            lcout => \c0.n18181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18112_bdd_4_lut_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__17829\,
            in1 => \N__17799\,
            in2 => \N__17793\,
            in3 => \N__28651\,
            lcout => OPEN,
            ltout => \c0.n18115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32148\,
            in1 => \N__17781\,
            in2 => \N__17769\,
            in3 => \N__21213\,
            lcout => \c0.n22_adj_2364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i151_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29992\,
            in1 => \N__17757\,
            in2 => \_gnd_net_\,
            in3 => \N__26546\,
            lcout => data_out_frame2_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__17745\,
            in1 => \N__21195\,
            in2 => \N__19773\,
            in3 => \N__32146\,
            lcout => \c0.n22_adj_2372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_515_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23564\,
            in2 => \_gnd_net_\,
            in3 => \N__23523\,
            lcout => \c0.n10548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_655_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23565\,
            in1 => \N__20395\,
            in2 => \_gnd_net_\,
            in3 => \N__23622\,
            lcout => \c0.n17249\,
            ltout => \c0.n17249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i156_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18117\,
            in1 => \N__18666\,
            in2 => \N__18102\,
            in3 => \N__18099\,
            lcout => \c0.data_out_frame2_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49639\,
            ce => \N__26543\,
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23025\,
            in1 => \N__18087\,
            in2 => \N__34325\,
            in3 => \N__21963\,
            lcout => \c0.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15151_3_lut_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__29052\,
            in1 => \_gnd_net_\,
            in2 => \N__28597\,
            in3 => \N__34318\,
            lcout => \c0.n17678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15004_2_lut_3_lut_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__40104\,
            in1 => \N__28483\,
            in2 => \_gnd_net_\,
            in3 => \N__29051\,
            lcout => \c0.n17586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i162_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17999\,
            in1 => \N__17961\,
            in2 => \N__20292\,
            in3 => \N__18867\,
            lcout => \c0.data_out_frame2_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49644\,
            ce => \N__26518\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_615_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17960\,
            in1 => \N__17916\,
            in2 => \N__23772\,
            in3 => \N__23261\,
            lcout => OPEN,
            ltout => \c0.n15_adj_2341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i153_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17898\,
            in1 => \N__18588\,
            in2 => \N__17886\,
            in3 => \N__23045\,
            lcout => \c0.data_out_frame2_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49644\,
            ce => \N__26518\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_717_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17883\,
            in1 => \N__21571\,
            in2 => \_gnd_net_\,
            in3 => \N__23260\,
            lcout => \c0.n17234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_596_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34725\,
            in1 => \N__23612\,
            in2 => \N__24003\,
            in3 => \N__23771\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i154_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18675\,
            in1 => \N__24798\,
            in2 => \N__18270\,
            in3 => \N__18267\,
            lcout => \c0.data_out_frame2_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49644\,
            ce => \N__26518\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i83_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31272\,
            in1 => \N__20234\,
            in2 => \_gnd_net_\,
            in3 => \N__26386\,
            lcout => data_out_frame2_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18058_bdd_4_lut_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__18240\,
            in1 => \N__18518\,
            in2 => \N__23563\,
            in3 => \N__28590\,
            lcout => \c0.n18061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_433_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40093\,
            in2 => \_gnd_net_\,
            in3 => \N__20453\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_434_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23851\,
            in1 => \N__21664\,
            in2 => \N__18234\,
            in3 => \N__21896\,
            lcout => \c0.n17258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_472_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18197\,
            in2 => \_gnd_net_\,
            in3 => \N__23185\,
            lcout => \c0.n17156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i91_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26385\,
            in1 => \_gnd_net_\,
            in2 => \N__18206\,
            in3 => \N__30783\,
            lcout => data_out_frame2_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19662\,
            in1 => \N__18176\,
            in2 => \N__18159\,
            in3 => \N__18144\,
            lcout => \c0.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i61_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26349\,
            in1 => \N__30657\,
            in2 => \_gnd_net_\,
            in3 => \N__19752\,
            lcout => data_out_frame2_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i149_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30109\,
            in1 => \N__18482\,
            in2 => \_gnd_net_\,
            in3 => \N__26351\,
            lcout => data_out_frame2_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i46_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26347\,
            in1 => \N__31515\,
            in2 => \_gnd_net_\,
            in3 => \N__18453\,
            lcout => data_out_frame2_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i60_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18411\,
            in1 => \N__30709\,
            in2 => \_gnd_net_\,
            in3 => \N__26352\,
            lcout => data_out_frame2_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i55_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26348\,
            in1 => \N__31030\,
            in2 => \_gnd_net_\,
            in3 => \N__40864\,
            lcout => data_out_frame2_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i141_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30656\,
            in1 => \N__18377\,
            in2 => \_gnd_net_\,
            in3 => \N__26350\,
            lcout => data_out_frame2_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i144_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26346\,
            in1 => \N__30467\,
            in2 => \_gnd_net_\,
            in3 => \N__18359\,
            lcout => data_out_frame2_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18345\,
            in1 => \N__21359\,
            in2 => \N__18333\,
            in3 => \N__21962\,
            lcout => \c0.n16_adj_2170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i54_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26378\,
            in1 => \N__31090\,
            in2 => \_gnd_net_\,
            in3 => \N__18295\,
            lcout => data_out_frame2_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i53_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31150\,
            in1 => \N__18787\,
            in2 => \_gnd_net_\,
            in3 => \N__26382\,
            lcout => data_out_frame2_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i56_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26379\,
            in1 => \N__30970\,
            in2 => \_gnd_net_\,
            in3 => \N__18649\,
            lcout => data_out_frame2_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i67_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30210\,
            in1 => \N__37238\,
            in2 => \_gnd_net_\,
            in3 => \N__26384\,
            lcout => data_out_frame2_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i51_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26377\,
            in1 => \N__31263\,
            in2 => \_gnd_net_\,
            in3 => \N__23814\,
            lcout => data_out_frame2_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i130_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30257\,
            in1 => \N__18617\,
            in2 => \_gnd_net_\,
            in3 => \N__26381\,
            lcout => data_out_frame2_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i99_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26380\,
            in1 => \N__30211\,
            in2 => \_gnd_net_\,
            in3 => \N__23902\,
            lcout => data_out_frame2_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i63_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30534\,
            in1 => \N__18828\,
            in2 => \_gnd_net_\,
            in3 => \N__26383\,
            lcout => data_out_frame2_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_610_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21353\,
            in1 => \N__18759\,
            in2 => \N__37252\,
            in3 => \N__20207\,
            lcout => \c0.n17153\,
            ltout => \c0.n17153_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18537\,
            in1 => \N__18579\,
            in2 => \N__18573\,
            in3 => \N__24282\,
            lcout => \c0.n26_adj_2203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i48_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26571\,
            in1 => \N__31399\,
            in2 => \_gnd_net_\,
            in3 => \N__18538\,
            lcout => data_out_frame2_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i108_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31618\,
            in1 => \N__18516\,
            in2 => \_gnd_net_\,
            in3 => \N__26573\,
            lcout => data_out_frame2_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_621_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18818\,
            in1 => \N__18780\,
            in2 => \_gnd_net_\,
            in3 => \N__24846\,
            lcout => \c0.n6_adj_2339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i79_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31449\,
            in1 => \N__21456\,
            in2 => \_gnd_net_\,
            in3 => \N__26575\,
            lcout => data_out_frame2_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i96_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26572\,
            in1 => \N__30447\,
            in2 => \_gnd_net_\,
            in3 => \N__23240\,
            lcout => data_out_frame2_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i77_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19884\,
            in1 => \N__31565\,
            in2 => \_gnd_net_\,
            in3 => \N__26574\,
            lcout => data_out_frame2_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i41_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26577\,
            in1 => \_gnd_net_\,
            in2 => \N__21304\,
            in3 => \N__30915\,
            lcout => data_out_frame2_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i122_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29810\,
            in1 => \N__23959\,
            in2 => \_gnd_net_\,
            in3 => \N__26579\,
            lcout => data_out_frame2_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i50_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26578\,
            in1 => \_gnd_net_\,
            in2 => \N__30351\,
            in3 => \N__23295\,
            lcout => data_out_frame2_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_665_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20620\,
            in1 => \N__21293\,
            in2 => \N__37254\,
            in3 => \N__20323\,
            lcout => \c0.n10507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_590_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23667\,
            in2 => \_gnd_net_\,
            in3 => \N__18731\,
            lcout => \c0.n17273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18046_bdd_4_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__28701\,
            in1 => \N__37245\,
            in2 => \N__18951\,
            in3 => \N__18912\,
            lcout => \c0.n18049\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i129_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26576\,
            in1 => \N__29459\,
            in2 => \_gnd_net_\,
            in3 => \N__24915\,
            lcout => data_out_frame2_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_459_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21794\,
            in1 => \N__18900\,
            in2 => \N__18882\,
            in3 => \N__18873\,
            lcout => \c0.n10_adj_2190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i0_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19119\,
            in2 => \_gnd_net_\,
            in3 => \N__33160\,
            lcout => \c0.FRAME_MATCHER_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49695\,
            ce => 'H',
            sr => \N__22437\
        );

    \c0.i1_2_lut_3_lut_adj_663_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18983\,
            in1 => \N__27835\,
            in2 => \_gnd_net_\,
            in3 => \N__41863\,
            lcout => \c0.n3_adj_2282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i5_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18966\,
            in2 => \_gnd_net_\,
            in3 => \N__33197\,
            lcout => \c0.FRAME_MATCHER_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49706\,
            ce => 'H',
            sr => \N__18855\
        );

    \c0.i2_3_lut_adj_656_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18981\,
            in1 => \N__19038\,
            in2 => \_gnd_net_\,
            in3 => \N__19074\,
            lcout => \c0.n15164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_552_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18982\,
            lcout => \c0.n43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_3_i3_2_lut_3_lut_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27839\,
            in1 => \N__19075\,
            in2 => \_gnd_net_\,
            in3 => \N__41864\,
            lcout => \c0.n3_adj_2227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_4_i3_2_lut_3_lut_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__41865\,
            in1 => \_gnd_net_\,
            in2 => \N__27843\,
            in3 => \N__19040\,
            lcout => \c0.n3_adj_2179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_407_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19039\,
            in2 => \_gnd_net_\,
            in3 => \N__41860\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_750_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__41862\,
            in1 => \N__19079\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_2_lut_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27048\,
            in1 => \N__37155\,
            in2 => \N__19545\,
            in3 => \N__19110\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_0\,
            ltout => OPEN,
            carryin => \bfn_4_27_0_\,
            carryout => \c0.n16079\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_3_lut_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__25377\,
            in1 => \N__19494\,
            in2 => \N__32872\,
            in3 => \N__19095\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_1\,
            ltout => OPEN,
            carryin => \c0.n16079\,
            carryout => \c0.n16080\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_4_lut_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22332\,
            in1 => \N__37088\,
            in2 => \N__19546\,
            in3 => \N__19092\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_2\,
            ltout => OPEN,
            carryin => \c0.n16080\,
            carryout => \c0.n16081\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_5_lut_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19089\,
            in1 => \N__19498\,
            in2 => \N__19083\,
            in3 => \N__19050\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_3\,
            ltout => OPEN,
            carryin => \c0.n16081\,
            carryout => \c0.n16082\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_6_lut_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__19047\,
            in1 => \N__19041\,
            in2 => \N__19547\,
            in3 => \N__18996\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_4\,
            ltout => OPEN,
            carryin => \c0.n16082\,
            carryout => \c0.n16083\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_7_lut_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__18993\,
            in1 => \N__19502\,
            in2 => \N__18987\,
            in3 => \N__18960\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_5\,
            ltout => OPEN,
            carryin => \c0.n16083\,
            carryout => \c0.n16084\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_8_lut_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20862\,
            in1 => \N__20880\,
            in2 => \N__19548\,
            in3 => \N__19200\,
            lcout => \c0.n3\,
            ltout => OPEN,
            carryin => \c0.n16084\,
            carryout => \c0.n16085\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_9_lut_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__27063\,
            in1 => \N__19506\,
            in2 => \N__27095\,
            in3 => \N__19191\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_7\,
            ltout => OPEN,
            carryin => \c0.n16085\,
            carryout => \c0.n16086\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_10_lut_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20892\,
            in1 => \N__19507\,
            in2 => \N__22192\,
            in3 => \N__19176\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_8\,
            ltout => OPEN,
            carryin => \bfn_4_28_0_\,
            carryout => \c0.n16087\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_11_lut_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20886\,
            in1 => \N__22632\,
            in2 => \N__19549\,
            in3 => \N__19173\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_9\,
            ltout => OPEN,
            carryin => \c0.n16087\,
            carryout => \c0.n16088\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_12_lut_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__27969\,
            in1 => \N__19511\,
            in2 => \N__28005\,
            in3 => \N__19170\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_10\,
            ltout => OPEN,
            carryin => \c0.n16088\,
            carryout => \c0.n16089\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_13_lut_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27114\,
            in1 => \N__27158\,
            in2 => \N__19550\,
            in3 => \N__19155\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_11\,
            ltout => OPEN,
            carryin => \c0.n16089\,
            carryout => \c0.n16090\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_14_lut_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19152\,
            in1 => \N__19515\,
            in2 => \N__25872\,
            in3 => \N__19146\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_12\,
            ltout => OPEN,
            carryin => \c0.n16090\,
            carryout => \c0.n16091\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_15_lut_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27174\,
            in1 => \N__27202\,
            in2 => \N__19551\,
            in3 => \N__19134\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_13\,
            ltout => OPEN,
            carryin => \c0.n16091\,
            carryout => \c0.n16092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_16_lut_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__27900\,
            in1 => \N__19519\,
            in2 => \N__27941\,
            in3 => \N__19278\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_14\,
            ltout => OPEN,
            carryin => \c0.n16092\,
            carryout => \c0.n16093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_17_lut_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27222\,
            in1 => \N__27263\,
            in2 => \N__19552\,
            in3 => \N__19263\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_15\,
            ltout => OPEN,
            carryin => \c0.n16093\,
            carryout => \c0.n16094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_18_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24954\,
            in1 => \N__27891\,
            in2 => \N__19553\,
            in3 => \N__19260\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_16\,
            ltout => OPEN,
            carryin => \bfn_4_29_0_\,
            carryout => \c0.n16095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_19_lut_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20781\,
            in1 => \N__20799\,
            in2 => \N__19557\,
            in3 => \N__19257\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_17\,
            ltout => OPEN,
            carryin => \c0.n16095\,
            carryout => \c0.n16096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_20_lut_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25404\,
            in1 => \N__25432\,
            in2 => \N__19554\,
            in3 => \N__19254\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_18\,
            ltout => OPEN,
            carryin => \c0.n16096\,
            carryout => \c0.n16097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_21_lut_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__24969\,
            in1 => \N__19529\,
            in2 => \N__25008\,
            in3 => \N__19239\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_19\,
            ltout => OPEN,
            carryin => \c0.n16097\,
            carryout => \c0.n16098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_22_lut_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25020\,
            in1 => \N__25059\,
            in2 => \N__19555\,
            in3 => \N__19224\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_20\,
            ltout => OPEN,
            carryin => \c0.n16098\,
            carryout => \c0.n16099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_23_lut_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20919\,
            in1 => \N__19533\,
            in2 => \N__20952\,
            in3 => \N__19212\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_21\,
            ltout => OPEN,
            carryin => \c0.n16099\,
            carryout => \c0.n16100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_24_lut_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25311\,
            in1 => \N__25327\,
            in2 => \N__19556\,
            in3 => \N__19203\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_22\,
            ltout => OPEN,
            carryin => \c0.n16100\,
            carryout => \c0.n16101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_25_lut_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__25074\,
            in1 => \N__19537\,
            in2 => \N__25124\,
            in3 => \N__19374\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_23\,
            ltout => OPEN,
            carryin => \c0.n16101\,
            carryout => \c0.n16102\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_26_lut_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25140\,
            in1 => \N__25170\,
            in2 => \N__19541\,
            in3 => \N__19371\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_24\,
            ltout => OPEN,
            carryin => \bfn_4_30_0_\,
            carryout => \c0.n16103\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_27_lut_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__25182\,
            in1 => \N__19478\,
            in2 => \N__25221\,
            in3 => \N__19368\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_25\,
            ltout => OPEN,
            carryin => \c0.n16103\,
            carryout => \c0.n16104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_28_lut_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25233\,
            in1 => \N__25281\,
            in2 => \N__19542\,
            in3 => \N__19365\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_26\,
            ltout => OPEN,
            carryin => \c0.n16104\,
            carryout => \c0.n16105\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_29_lut_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__20913\,
            in1 => \N__19482\,
            in2 => \N__22698\,
            in3 => \N__19362\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_27\,
            ltout => OPEN,
            carryin => \c0.n16105\,
            carryout => \c0.n16106\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_30_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__26997\,
            in1 => \N__27024\,
            in2 => \N__19543\,
            in3 => \N__19350\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_28\,
            ltout => OPEN,
            carryin => \c0.n16106\,
            carryout => \c0.n16107\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_31_lut_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19347\,
            in1 => \N__19486\,
            in2 => \N__19335\,
            in3 => \N__19302\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_29\,
            ltout => OPEN,
            carryin => \c0.n16107\,
            carryout => \c0.n16108\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_32_lut_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__33618\,
            in1 => \N__33651\,
            in2 => \N__19544\,
            in3 => \N__19293\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_30\,
            ltout => OPEN,
            carryin => \c0.n16108\,
            carryout => \c0.n16109\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_977_33_lut_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__29542\,
            in1 => \N__19490\,
            in2 => \N__21039\,
            in3 => \N__19290\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1278_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__37852\,
            in1 => \N__25624\,
            in2 => \_gnd_net_\,
            in3 => \N__21119\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2593_2_lut_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37851\,
            in2 => \_gnd_net_\,
            in3 => \N__37933\,
            lcout => n5244,
            ltout => \n5244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14631_3_lut_4_lut_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100101010"
        )
    port map (
            in0 => \N__25544\,
            in1 => \N__37902\,
            in2 => \N__19563\,
            in3 => \N__25623\,
            lcout => n11018,
            ltout => \n11018_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000001000000"
        )
    port map (
            in0 => \N__25625\,
            in1 => \N__37853\,
            in2 => \N__19560\,
            in3 => \N__37934\,
            lcout => \r_Bit_Index_1_adj_2436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15231_1_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39016\,
            lcout => \c0.n18008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15224_2_lut_3_lut_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__25484\,
            in1 => \N__25545\,
            in2 => \_gnd_net_\,
            in3 => \N__31851\,
            lcout => \c0.rx.n17058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111111"
        )
    port map (
            in0 => \N__21131\,
            in1 => \N__37903\,
            in2 => \N__25602\,
            in3 => \N__25485\,
            lcout => OPEN,
            ltout => \n13692_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__31852\,
            in1 => \N__25546\,
            in2 => \N__19392\,
            in3 => \N__21009\,
            lcout => \c0.rx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22559\,
            in2 => \_gnd_net_\,
            in3 => \N__19389\,
            lcout => \c0.rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_4_32_0_\,
            carryout => \c0.rx.n16125\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i1_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20991\,
            in2 => \_gnd_net_\,
            in3 => \N__19608\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.rx.n16125\,
            carryout => \c0.rx.n16126\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i2_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22574\,
            in2 => \_gnd_net_\,
            in3 => \N__19605\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.rx.n16126\,
            carryout => \c0.rx.n16127\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i3_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22541\,
            in2 => \_gnd_net_\,
            in3 => \N__19602\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.rx.n16127\,
            carryout => \c0.rx.n16128\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i4_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21003\,
            in2 => \_gnd_net_\,
            in3 => \N__19599\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.rx.n16128\,
            carryout => \c0.rx.n16129\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i5_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31933\,
            in2 => \_gnd_net_\,
            in3 => \N__19596\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.rx.n16129\,
            carryout => \c0.rx.n16130\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i6_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31726\,
            in2 => \_gnd_net_\,
            in3 => \N__19593\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.rx.n16130\,
            carryout => \c0.rx.n16131\,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.rx.r_Clock_Count__i7_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31767\,
            in2 => \_gnd_net_\,
            in3 => \N__19590\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49776\,
            ce => \N__20979\,
            sr => \N__21018\
        );

    \c0.data_out_frame2_0___i146_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30264\,
            in1 => \N__19586\,
            in2 => \_gnd_net_\,
            in3 => \N__26517\,
            lcout => data_out_frame2_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i7_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__26664\,
            in1 => \N__39702\,
            in2 => \N__34477\,
            in3 => \N__42095\,
            lcout => \c0.byte_transmit_counter2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49645\,
            ce => 'H',
            sr => \N__32043\
        );

    \c0.i5_3_lut_4_lut_adj_690_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19830\,
            in1 => \N__21524\,
            in2 => \N__19971\,
            in3 => \N__19904\,
            lcout => OPEN,
            ltout => \c0.n14_adj_2188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i163_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20043\,
            in1 => \N__19722\,
            in2 => \N__19791\,
            in3 => \N__19788\,
            lcout => \c0.data_out_frame2_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49634\,
            ce => \N__26544\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_447_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40290\,
            in2 => \_gnd_net_\,
            in3 => \N__23999\,
            lcout => \c0.n17294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_470_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19764\,
            lcout => \c0.n17240\,
            ltout => \c0.n17240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i161_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20478\,
            in1 => \N__20265\,
            in2 => \N__19716\,
            in3 => \N__19713\,
            lcout => \c0.data_out_frame2_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49634\,
            ce => \N__26544\,
            sr => \_gnd_net_\
        );

    \c0.i15015_3_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__28648\,
            in1 => \N__40672\,
            in2 => \_gnd_net_\,
            in3 => \N__28972\,
            lcout => \c0.n17603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14662_3_lut_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001000100"
        )
    port map (
            in0 => \N__28971\,
            in1 => \N__37636\,
            in2 => \_gnd_net_\,
            in3 => \N__28647\,
            lcout => \c0.n17439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i158_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19977\,
            in1 => \N__19614\,
            in2 => \N__19686\,
            in3 => \N__20138\,
            lcout => \c0.data_out_frame2_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49646\,
            ce => \N__26542\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_531_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19836\,
            in1 => \N__19661\,
            in2 => \N__19631\,
            in3 => \N__24845\,
            lcout => \c0.n15_adj_2291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_710_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24080\,
            in1 => \N__26645\,
            in2 => \N__23922\,
            in3 => \N__41107\,
            lcout => \c0.n17288\,
            ltout => \c0.n17288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_671_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23381\,
            in1 => \N__20034\,
            in2 => \N__19980\,
            in3 => \N__26055\,
            lcout => \c0.n14_adj_2292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_523_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26646\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24081\,
            lcout => OPEN,
            ltout => \c0.n10428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i164_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19970\,
            in1 => \N__20624\,
            in2 => \N__19956\,
            in3 => \N__19953\,
            lcout => \c0.data_out_frame2_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49646\,
            ce => \N__26542\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_522_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23918\,
            lcout => \c0.n10504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i90_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26415\,
            in2 => \N__20080\,
            in3 => \N__29812\,
            lcout => data_out_frame2_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i138_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__29811\,
            in1 => \N__19922\,
            in2 => \N__26547\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18208_bdd_4_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__28649\,
            in1 => \N__24380\,
            in2 => \N__19903\,
            in3 => \N__21687\,
            lcout => \c0.n17568\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_529_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21311\,
            in2 => \_gnd_net_\,
            in3 => \N__20521\,
            lcout => \c0.n10554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_486_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20288\,
            in1 => \N__20183\,
            in2 => \N__24555\,
            in3 => \N__20431\,
            lcout => \c0.n15_adj_2205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__20256\,
            in1 => \N__28650\,
            in2 => \N__23522\,
            in3 => \N__29053\,
            lcout => \c0.n6_adj_2139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_609_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23602\,
            in1 => \N__20106\,
            in2 => \_gnd_net_\,
            in3 => \N__20229\,
            lcout => \c0.n10492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_714_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20182\,
            in1 => \N__23744\,
            in2 => \_gnd_net_\,
            in3 => \N__21752\,
            lcout => \c0.n17255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i133_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30105\,
            in1 => \N__26363\,
            in2 => \_gnd_net_\,
            in3 => \N__20113\,
            lcout => data_out_frame2_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i98_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26361\,
            in1 => \_gnd_net_\,
            in2 => \N__30274\,
            in3 => \N__23613\,
            lcout => data_out_frame2_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i94_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30594\,
            in1 => \N__26364\,
            in2 => \_gnd_net_\,
            in3 => \N__21866\,
            lcout => data_out_frame2_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i93_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26360\,
            in1 => \N__30646\,
            in2 => \_gnd_net_\,
            in3 => \N__21897\,
            lcout => data_out_frame2_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_445_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20064\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24744\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_446_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21745\,
            in1 => \N__20474\,
            in2 => \N__20463\,
            in3 => \N__24036\,
            lcout => \c0.n10229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i103_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29991\,
            in1 => \N__26362\,
            in2 => \_gnd_net_\,
            in3 => \N__22962\,
            lcout => data_out_frame2_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i68_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26359\,
            in1 => \N__30158\,
            in2 => \_gnd_net_\,
            in3 => \N__24832\,
            lcout => data_out_frame2_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i76_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24636\,
            in1 => \N__31623\,
            in2 => \_gnd_net_\,
            in3 => \N__26337\,
            lcout => data_out_frame2_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_4_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40248\,
            in1 => \N__36092\,
            in2 => \N__33687\,
            in3 => \N__39758\,
            lcout => n10725,
            ltout => \n10725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i104_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29916\,
            in2 => \N__20442\,
            in3 => \N__20424\,
            lcout => data_out_frame2_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i84_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26335\,
            in1 => \N__31194\,
            in2 => \_gnd_net_\,
            in3 => \N__20379\,
            lcout => data_out_frame2_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15316_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__28641\,
            in1 => \N__28959\,
            in2 => \N__24073\,
            in3 => \N__21868\,
            lcout => \c0.n18106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i131_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26334\,
            in1 => \N__30215\,
            in2 => \_gnd_net_\,
            in3 => \N__20322\,
            lcout => data_out_frame2_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i123_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30780\,
            in1 => \N__20612\,
            in2 => \_gnd_net_\,
            in3 => \N__26336\,
            lcout => data_out_frame2_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i124_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26333\,
            in1 => \N__30708\,
            in2 => \_gnd_net_\,
            in3 => \N__24422\,
            lcout => data_out_frame2_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i137_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29861\,
            in1 => \N__26343\,
            in2 => \_gnd_net_\,
            in3 => \N__21713\,
            lcout => data_out_frame2_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i147_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26340\,
            in1 => \N__30209\,
            in2 => \_gnd_net_\,
            in3 => \N__20576\,
            lcout => data_out_frame2_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i89_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29862\,
            in1 => \N__26345\,
            in2 => \_gnd_net_\,
            in3 => \N__24743\,
            lcout => data_out_frame2_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i134_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26339\,
            in1 => \N__30039\,
            in2 => \_gnd_net_\,
            in3 => \N__20547\,
            lcout => data_out_frame2_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i81_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30406\,
            in1 => \N__26344\,
            in2 => \_gnd_net_\,
            in3 => \N__21360\,
            lcout => data_out_frame2_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i125_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26338\,
            in1 => \N__30645\,
            in2 => \_gnd_net_\,
            in3 => \N__20513\,
            lcout => data_out_frame2_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i120_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30960\,
            in1 => \N__26342\,
            in2 => \_gnd_net_\,
            in3 => \N__22094\,
            lcout => data_out_frame2_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i71_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26341\,
            in1 => \N__29966\,
            in2 => \_gnd_net_\,
            in3 => \N__21509\,
            lcout => data_out_frame2_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i0_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29431\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => rand_data_0,
            ltout => OPEN,
            carryin => \bfn_5_23_0_\,
            carryout => n15979,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i1_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30250\,
            in2 => \_gnd_net_\,
            in3 => \N__20649\,
            lcout => rand_data_1,
            ltout => OPEN,
            carryin => n15979,
            carryout => n15980,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i2_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30205\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => rand_data_2,
            ltout => OPEN,
            carryin => n15980,
            carryout => n15981,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i3_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30143\,
            in2 => \_gnd_net_\,
            in3 => \N__20643\,
            lcout => rand_data_3,
            ltout => OPEN,
            carryin => n15981,
            carryout => n15982,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i4_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30088\,
            in2 => \_gnd_net_\,
            in3 => \N__20640\,
            lcout => rand_data_4,
            ltout => OPEN,
            carryin => n15982,
            carryout => n15983,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i5_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30031\,
            in2 => \_gnd_net_\,
            in3 => \N__20637\,
            lcout => rand_data_5,
            ltout => OPEN,
            carryin => n15983,
            carryout => n15984,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i6_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29965\,
            in2 => \_gnd_net_\,
            in3 => \N__20634\,
            lcout => rand_data_6,
            ltout => OPEN,
            carryin => n15984,
            carryout => n15985,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i7_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29903\,
            in2 => \_gnd_net_\,
            in3 => \N__20631\,
            lcout => rand_data_7,
            ltout => OPEN,
            carryin => n15985,
            carryout => n15986,
            clk => \N__49685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i8_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29846\,
            in2 => \_gnd_net_\,
            in3 => \N__20628\,
            lcout => rand_data_8,
            ltout => OPEN,
            carryin => \bfn_5_24_0_\,
            carryout => n15987,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i9_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29783\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => rand_data_9,
            ltout => OPEN,
            carryin => n15987,
            carryout => n15988,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i10_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30751\,
            in2 => \_gnd_net_\,
            in3 => \N__20676\,
            lcout => rand_data_10,
            ltout => OPEN,
            carryin => n15988,
            carryout => n15989,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i11_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30681\,
            in2 => \_gnd_net_\,
            in3 => \N__20673\,
            lcout => rand_data_11,
            ltout => OPEN,
            carryin => n15989,
            carryout => n15990,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i12_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30629\,
            in2 => \_gnd_net_\,
            in3 => \N__20670\,
            lcout => rand_data_12,
            ltout => OPEN,
            carryin => n15990,
            carryout => n15991,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i13_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30574\,
            in2 => \_gnd_net_\,
            in3 => \N__20667\,
            lcout => rand_data_13,
            ltout => OPEN,
            carryin => n15991,
            carryout => n15992,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i14_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30502\,
            in2 => \_gnd_net_\,
            in3 => \N__20664\,
            lcout => rand_data_14,
            ltout => OPEN,
            carryin => n15992,
            carryout => n15993,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i15_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30446\,
            in2 => \_gnd_net_\,
            in3 => \N__20661\,
            lcout => rand_data_15,
            ltout => OPEN,
            carryin => n15993,
            carryout => n15994,
            clk => \N__49696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i16_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30392\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => rand_data_16,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => n15995,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i17_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30329\,
            in2 => \_gnd_net_\,
            in3 => \N__20655\,
            lcout => rand_data_17,
            ltout => OPEN,
            carryin => n15995,
            carryout => n15996,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i18_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31238\,
            in2 => \_gnd_net_\,
            in3 => \N__20706\,
            lcout => rand_data_18,
            ltout => OPEN,
            carryin => n15996,
            carryout => n15997,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i19_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31181\,
            in2 => \_gnd_net_\,
            in3 => \N__20703\,
            lcout => rand_data_19,
            ltout => OPEN,
            carryin => n15997,
            carryout => n15998,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i20_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31127\,
            in2 => \_gnd_net_\,
            in3 => \N__20700\,
            lcout => rand_data_20,
            ltout => OPEN,
            carryin => n15998,
            carryout => n15999,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i21_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31064\,
            in2 => \_gnd_net_\,
            in3 => \N__20697\,
            lcout => rand_data_21,
            ltout => OPEN,
            carryin => n15999,
            carryout => n16000,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i22_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31002\,
            in2 => \_gnd_net_\,
            in3 => \N__20694\,
            lcout => rand_data_22,
            ltout => OPEN,
            carryin => n16000,
            carryout => n16001,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i23_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30948\,
            in2 => \_gnd_net_\,
            in3 => \N__20691\,
            lcout => rand_data_23,
            ltout => OPEN,
            carryin => n16001,
            carryout => n16002,
            clk => \N__49707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i24_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30899\,
            in2 => \_gnd_net_\,
            in3 => \N__20688\,
            lcout => rand_data_24,
            ltout => OPEN,
            carryin => \bfn_5_26_0_\,
            carryout => n16003,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i25_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30810\,
            in2 => \_gnd_net_\,
            in3 => \N__20685\,
            lcout => rand_data_25,
            ltout => OPEN,
            carryin => n16003,
            carryout => n16004,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i26_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31655\,
            in2 => \_gnd_net_\,
            in3 => \N__20682\,
            lcout => rand_data_26,
            ltout => OPEN,
            carryin => n16004,
            carryout => n16005,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i27_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31596\,
            in2 => \_gnd_net_\,
            in3 => \N__20742\,
            lcout => rand_data_27,
            ltout => OPEN,
            carryin => n16005,
            carryout => n16006,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i28_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31544\,
            in2 => \_gnd_net_\,
            in3 => \N__20739\,
            lcout => rand_data_28,
            ltout => OPEN,
            carryin => n16006,
            carryout => n16007,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i29_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31482\,
            in2 => \_gnd_net_\,
            in3 => \N__20736\,
            lcout => rand_data_29,
            ltout => OPEN,
            carryin => n16007,
            carryout => n16008,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i30_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31430\,
            in2 => \_gnd_net_\,
            in3 => \N__20733\,
            lcout => rand_data_30,
            ltout => OPEN,
            carryin => n16008,
            carryout => n16009,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_2358__i31_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31376\,
            in2 => \_gnd_net_\,
            in3 => \N__20730\,
            lcout => rand_data_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i6_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20727\,
            in2 => \_gnd_net_\,
            in3 => \N__33218\,
            lcout => \c0.FRAME_MATCHER_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49731\,
            ce => 'H',
            sr => \N__20718\
        );

    \c0.i1_2_lut_adj_659_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25288\,
            in2 => \_gnd_net_\,
            in3 => \N__20877\,
            lcout => OPEN,
            ltout => \c0.n26_adj_2373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_669_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24993\,
            in1 => \N__27147\,
            in2 => \N__20721\,
            in3 => \N__27258\,
            lcout => \c0.n44_adj_2378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_652_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__41883\,
            in1 => \_gnd_net_\,
            in2 => \N__27830\,
            in3 => \N__20879\,
            lcout => \c0.n3_adj_2280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_579_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41882\,
            lcout => \c0.n41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_15_i3_2_lut_3_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__41885\,
            in1 => \_gnd_net_\,
            in2 => \N__27831\,
            in3 => \N__27259\,
            lcout => \c0.n3_adj_2261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_11_i3_2_lut_3_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__27151\,
            in1 => \N__27786\,
            in2 => \_gnd_net_\,
            in3 => \N__41884\,
            lcout => \c0.n3_adj_2270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_19_i3_2_lut_3_lut_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__41886\,
            in1 => \_gnd_net_\,
            in2 => \N__27832\,
            in3 => \N__24994\,
            lcout => \c0.n3_adj_2252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_660_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25054\,
            in1 => \N__20946\,
            in2 => \N__25119\,
            in3 => \N__20796\,
            lcout => \c0.n42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i17_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20814\,
            in2 => \_gnd_net_\,
            in3 => \N__33235\,
            lcout => \c0.FRAME_MATCHER_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49741\,
            ce => 'H',
            sr => \N__20808\
        );

    \c0.select_219_Select_17_i3_2_lut_3_lut_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41878\,
            in1 => \N__27796\,
            in2 => \_gnd_net_\,
            in3 => \N__20798\,
            lcout => \c0.n3_adj_2257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10671_2_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41877\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_21_i3_2_lut_3_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41880\,
            in1 => \N__27795\,
            in2 => \_gnd_net_\,
            in3 => \N__20948\,
            lcout => \c0.n3_adj_2248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_20_i3_2_lut_3_lut_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27793\,
            in1 => \N__25055\,
            in2 => \_gnd_net_\,
            in3 => \N__41879\,
            lcout => \c0.n3_adj_2250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_23_i3_2_lut_3_lut_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41881\,
            in1 => \_gnd_net_\,
            in2 => \N__25120\,
            in3 => \N__27794\,
            lcout => \c0.n3_adj_2244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10667_2_lut_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20947\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41876\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i6_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45019\,
            in1 => \N__44811\,
            in2 => \N__27395\,
            in3 => \N__44542\,
            lcout => \c0.FRAME_MATCHER_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49752\,
            ce => 'H',
            sr => \N__27363\
        );

    \c0.select_219_Select_27_i3_2_lut_3_lut_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41870\,
            in1 => \_gnd_net_\,
            in2 => \N__22693\,
            in3 => \N__27781\,
            lcout => \c0.n3_adj_2236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_686_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22683\,
            in2 => \_gnd_net_\,
            in3 => \N__41866\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_8_i3_2_lut_3_lut_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41871\,
            in1 => \N__27780\,
            in2 => \_gnd_net_\,
            in3 => \N__22194\,
            lcout => \c0.n3_adj_2276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10680_2_lut_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22193\,
            in2 => \_gnd_net_\,
            in3 => \N__41869\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_9_i3_2_lut_3_lut_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__41872\,
            in1 => \N__22631\,
            in2 => \_gnd_net_\,
            in3 => \N__27782\,
            lcout => \c0.n3_adj_2274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10679_2_lut_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41868\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10657_2_lut_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29564\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i25_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21030\,
            in2 => \_gnd_net_\,
            in3 => \N__33236\,
            lcout => \c0.FRAME_MATCHER_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49765\,
            ce => 'H',
            sr => \N__22476\
        );

    \c0.FRAME_MATCHER_i_i26_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21024\,
            in2 => \_gnd_net_\,
            in3 => \N__33250\,
            lcout => \c0.FRAME_MATCHER_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49777\,
            ce => 'H',
            sr => \N__25257\
        );

    \c0.rx.i1_4_lut_adj_396_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__31866\,
            in1 => \N__22587\,
            in2 => \N__25560\,
            in3 => \N__22512\,
            lcout => \c0.rx.n10845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__25551\,
            in1 => \N__31868\,
            in2 => \N__39059\,
            in3 => \N__25638\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__25487\,
            in1 => \N__45267\,
            in2 => \_gnd_net_\,
            in3 => \N__22854\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21002\,
            in2 => \_gnd_net_\,
            in3 => \N__20990\,
            lcout => \c0.rx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15215_4_lut_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__25486\,
            in1 => \N__25550\,
            in2 => \N__31869\,
            in3 => \N__22839\,
            lcout => \c0.rx.n10656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15089_2_lut_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25488\,
            in2 => \_gnd_net_\,
            in3 => \N__25598\,
            lcout => OPEN,
            ltout => \n17708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000010101"
        )
    port map (
            in0 => \N__31867\,
            in1 => \N__25552\,
            in2 => \N__21135\,
            in3 => \N__22581\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010000000000"
        )
    port map (
            in0 => \N__25626\,
            in1 => \N__21132\,
            in2 => \N__37907\,
            in3 => \N__21120\,
            lcout => \r_Bit_Index_2_adj_2435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6489_2_lut_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28585\,
            in2 => \_gnd_net_\,
            in3 => \N__28932\,
            lcout => \c0.n9157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__21108\,
            in2 => \N__21699\,
            in3 => \N__21211\,
            lcout => \c0.n22_adj_2387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__23787\,
            in1 => \N__28613\,
            in2 => \N__24177\,
            in3 => \N__29003\,
            lcout => \c0.n6_adj_2140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15435_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21102\,
            in1 => \N__32369\,
            in2 => \N__21087\,
            in3 => \N__32141\,
            lcout => OPEN,
            ltout => \c0.n18244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18244_bdd_4_lut_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32370\,
            in1 => \N__21072\,
            in2 => \N__21060\,
            in3 => \N__21057\,
            lcout => \c0.n18247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__21582\,
            in1 => \N__22812\,
            in2 => \N__25794\,
            in3 => \N__25736\,
            lcout => OPEN,
            ltout => \c0.tx2.n18232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n18232_bdd_4_lut_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__21399\,
            in1 => \N__21051\,
            in2 => \N__21042\,
            in3 => \N__25791\,
            lcout => \c0.tx2.n18235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__21375\,
            in1 => \N__32414\,
            in2 => \N__32276\,
            in3 => \N__21405\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49640\,
            ce => \N__24265\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15420_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__21393\,
            in1 => \N__32412\,
            in2 => \N__21321\,
            in3 => \N__32149\,
            lcout => OPEN,
            ltout => \c0.n18226_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18226_bdd_4_lut_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32413\,
            in1 => \N__21384\,
            in2 => \N__21378\,
            in3 => \N__21246\,
            lcout => \c0.n18229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15351_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__21368\,
            in1 => \N__28891\,
            in2 => \N__28661\,
            in3 => \N__24750\,
            lcout => OPEN,
            ltout => \c0.n18148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18148_bdd_4_lut_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__41108\,
            in1 => \N__24323\,
            in2 => \N__21324\,
            in3 => \N__28610\,
            lcout => \c0.n18151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__28611\,
            in1 => \N__21312\,
            in2 => \N__21267\,
            in3 => \N__28892\,
            lcout => \c0.n6_adj_2143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15274_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21416\,
            in1 => \N__28614\,
            in2 => \N__21240\,
            in3 => \N__28938\,
            lcout => OPEN,
            ltout => \c0.n18052_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18052_bdd_4_lut_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__28615\,
            in1 => \N__21681\,
            in2 => \N__21228\,
            in3 => \N__24481\,
            lcout => OPEN,
            ltout => \c0.n18055_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32167\,
            in1 => \N__21225\,
            in2 => \N__21216\,
            in3 => \N__21194\,
            lcout => \c0.n22_adj_2371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_15440_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23322\,
            in1 => \N__32415\,
            in2 => \N__21615\,
            in3 => \N__32168\,
            lcout => OPEN,
            ltout => \c0.n18256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18256_bdd_4_lut_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32416\,
            in1 => \N__28716\,
            in2 => \N__21600\,
            in3 => \N__21597\,
            lcout => OPEN,
            ltout => \c0.n18259_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__21591\,
            in1 => \N__32417\,
            in2 => \N__21585\,
            in3 => \N__32277\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49652\,
            ce => \N__24254\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i82_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26514\,
            in1 => \N__30363\,
            in2 => \_gnd_net_\,
            in3 => \N__21564\,
            lcout => data_out_frame2_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i42_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23397\,
            in1 => \N__30842\,
            in2 => \_gnd_net_\,
            in3 => \N__26516\,
            lcout => data_out_frame2_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_680_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23137\,
            in1 => \N__21860\,
            in2 => \_gnd_net_\,
            in3 => \N__21895\,
            lcout => \c0.n17203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18124_bdd_4_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__21523\,
            in1 => \N__23103\,
            in2 => \N__21474\,
            in3 => \N__28505\,
            lcout => \c0.n18127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i148_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26513\,
            in1 => \N__30169\,
            in2 => \_gnd_net_\,
            in3 => \N__21417\,
            lcout => data_out_frame2_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i136_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29931\,
            in1 => \N__27635\,
            in2 => \_gnd_net_\,
            in3 => \N__26515\,
            lcout => data_out_frame2_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18160_bdd_4_lut_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__28506\,
            in1 => \N__23073\,
            in2 => \N__21717\,
            in3 => \N__24941\,
            lcout => \c0.n18163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15450_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__21894\,
            in1 => \N__28504\,
            in2 => \N__24138\,
            in3 => \N__28999\,
            lcout => \c0.n18208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i140_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30717\,
            in1 => \N__21680\,
            in2 => \_gnd_net_\,
            in3 => \N__26370\,
            lcout => data_out_frame2_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i127_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26366\,
            in1 => \N__30536\,
            in2 => \_gnd_net_\,
            in3 => \N__23012\,
            lcout => data_out_frame2_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i145_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23085\,
            in1 => \N__29454\,
            in2 => \_gnd_net_\,
            in3 => \N__26371\,
            lcout => data_out_frame2_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i87_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26368\,
            in1 => \N__31026\,
            in2 => \_gnd_net_\,
            in3 => \N__23184\,
            lcout => data_out_frame2_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i106_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30834\,
            in1 => \N__23652\,
            in2 => \_gnd_net_\,
            in3 => \N__26369\,
            lcout => data_out_frame2_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i115_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26365\,
            in1 => \N__31264\,
            in2 => \_gnd_net_\,
            in3 => \N__21660\,
            lcout => data_out_frame2_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_724_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41098\,
            in1 => \N__41149\,
            in2 => \N__21787\,
            in3 => \N__21630\,
            lcout => \c0.n17095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i59_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26367\,
            in1 => \N__30782\,
            in2 => \_gnd_net_\,
            in3 => \N__23844\,
            lcout => data_out_frame2_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i43_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26353\,
            in1 => \N__31674\,
            in2 => \_gnd_net_\,
            in3 => \N__24163\,
            lcout => data_out_frame2_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i119_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24526\,
            in1 => \_gnd_net_\,
            in2 => \N__31032\,
            in3 => \N__26356\,
            lcout => data_out_frame2_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i85_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26355\,
            in1 => \N__31149\,
            in2 => \_gnd_net_\,
            in3 => \N__24133\,
            lcout => data_out_frame2_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_672_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23123\,
            in1 => \N__21893\,
            in2 => \N__21867\,
            in3 => \N__24024\,
            lcout => \c0.n10359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i45_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26354\,
            in1 => \N__31564\,
            in2 => \_gnd_net_\,
            in3 => \N__21783\,
            lcout => data_out_frame2_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i95_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__23124\,
            in1 => \_gnd_net_\,
            in2 => \N__30537\,
            in3 => \N__26358\,
            lcout => data_out_frame2_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15346_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__23255\,
            in1 => \N__21740\,
            in2 => \N__28599\,
            in3 => \N__28960\,
            lcout => \c0.n18142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i88_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21741\,
            in1 => \N__30975\,
            in2 => \_gnd_net_\,
            in3 => \N__26357\,
            lcout => data_out_frame2_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i11067_2_lut_4_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__22145\,
            in1 => \N__26839\,
            in2 => \N__22287\,
            in3 => \N__22044\,
            lcout => OPEN,
            ltout => \c0.tx2.n13748_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__26742\,
            in1 => \N__25941\,
            in2 => \N__22008\,
            in3 => \N__22068\,
            lcout => \c0.tx2.n17322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i73_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__26374\,
            in1 => \N__30919\,
            in2 => \N__41105\,
            in3 => \_gnd_net_\,
            lcout => data_out_frame2_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i152_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29912\,
            in1 => \N__22001\,
            in2 => \_gnd_net_\,
            in3 => \N__26376\,
            lcout => data_out_frame2_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i139_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26372\,
            in1 => \N__30781\,
            in2 => \_gnd_net_\,
            in3 => \N__21977\,
            lcout => data_out_frame2_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_4_lut_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__22043\,
            in1 => \N__22067\,
            in2 => \N__22146\,
            in3 => \N__22283\,
            lcout => \r_SM_Main_2_N_2031_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i70_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26373\,
            in1 => \N__30032\,
            in2 => \_gnd_net_\,
            in3 => \N__40925\,
            lcout => data_out_frame2_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i109_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31563\,
            in1 => \N__41144\,
            in2 => \_gnd_net_\,
            in3 => \N__26375\,
            lcout => data_out_frame2_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i62_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21955\,
            in1 => \N__30584\,
            in2 => \_gnd_net_\,
            in3 => \N__26566\,
            lcout => data_out_frame2_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49697\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i69_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26565\,
            in1 => \N__30104\,
            in2 => \_gnd_net_\,
            in3 => \N__24358\,
            lcout => data_out_frame2_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49697\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i4_4_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22058\,
            in1 => \N__22323\,
            in2 => \N__22305\,
            in3 => \N__22022\,
            lcout => \c0.tx2.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22114\,
            in1 => \N__25672\,
            in2 => \_gnd_net_\,
            in3 => \N__22719\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49697\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i65_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29453\,
            in1 => \N__24316\,
            in2 => \_gnd_net_\,
            in3 => \N__26567\,
            lcout => data_out_frame2_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49697\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_613_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24596\,
            in2 => \_gnd_net_\,
            in3 => \N__22093\,
            lcout => \c0.n10563\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15218_2_lut_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22074\,
            in2 => \_gnd_net_\,
            in3 => \N__26852\,
            lcout => \c0.tx2.n10852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22230\,
            in1 => \N__22262\,
            in2 => \_gnd_net_\,
            in3 => \N__22247\,
            lcout => \c0.tx2.n17018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22059\,
            in2 => \_gnd_net_\,
            in3 => \N__22047\,
            lcout => \c0.tx2.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_6_24_0_\,
            carryout => \c0.tx2.n16132\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i1_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22042\,
            in2 => \_gnd_net_\,
            in3 => \N__22026\,
            lcout => \c0.tx2.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.tx2.n16132\,
            carryout => \c0.tx2.n16133\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i2_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22023\,
            in2 => \_gnd_net_\,
            in3 => \N__22011\,
            lcout => \c0.tx2.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.tx2.n16133\,
            carryout => \c0.tx2.n16134\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i3_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22322\,
            in2 => \_gnd_net_\,
            in3 => \N__22308\,
            lcout => \c0.tx2.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.tx2.n16134\,
            carryout => \c0.tx2.n16135\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i4_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22304\,
            in2 => \_gnd_net_\,
            in3 => \N__22290\,
            lcout => \c0.tx2.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.tx2.n16135\,
            carryout => \c0.tx2.n16136\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i5_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22282\,
            in2 => \_gnd_net_\,
            in3 => \N__22266\,
            lcout => \c0.tx2.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.tx2.n16136\,
            carryout => \c0.tx2.n16137\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i6_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22263\,
            in2 => \_gnd_net_\,
            in3 => \N__22251\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.tx2.n16137\,
            carryout => \c0.tx2.n16138\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i7_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22248\,
            in2 => \_gnd_net_\,
            in3 => \N__22236\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \c0.tx2.n16138\,
            carryout => \c0.tx2.n16139\,
            clk => \N__49708\,
            ce => \N__25676\,
            sr => \N__22215\
        );

    \c0.tx2.r_Clock_Count__i8_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22229\,
            in2 => \_gnd_net_\,
            in3 => \N__22233\,
            lcout => \c0.tx2.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49721\,
            ce => \N__25677\,
            sr => \N__22214\
        );

    \c0.i14_4_lut_adj_668_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22694\,
            in1 => \N__25431\,
            in2 => \N__25342\,
            in3 => \N__27996\,
            lcout => \c0.n39_adj_2377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_639_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37077\,
            in2 => \_gnd_net_\,
            in3 => \N__22373\,
            lcout => \c0.n10161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_666_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22626\,
            in1 => \N__27928\,
            in2 => \N__27890\,
            in3 => \N__22182\,
            lcout => OPEN,
            ltout => \c0.n41_adj_2376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22416\,
            in1 => \N__22506\,
            in2 => \N__22407\,
            in3 => \N__22404\,
            lcout => OPEN,
            ltout => \c0.n48_adj_2379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_675_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22398\,
            in1 => \N__32791\,
            in2 => \N__22386\,
            in3 => \N__22383\,
            lcout => \c0.n9995\,
            ltout => \c0.n9995_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10584_4_lut_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__29560\,
            in1 => \N__32865\,
            in2 => \N__22377\,
            in3 => \N__32640\,
            lcout => n3779,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10579_2_lut_3_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__37079\,
            in1 => \N__29558\,
            in2 => \_gnd_net_\,
            in3 => \N__22374\,
            lcout => n4408,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i2_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22362\,
            in2 => \_gnd_net_\,
            in3 => \N__33185\,
            lcout => \c0.FRAME_MATCHER_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49742\,
            ce => 'H',
            sr => \N__22353\
        );

    \c0.select_219_Select_2_i3_2_lut_3_lut_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__37081\,
            in1 => \_gnd_net_\,
            in2 => \N__27833\,
            in3 => \N__41874\,
            lcout => \c0.n3_adj_2286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_31_i3_2_lut_3_lut_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41875\,
            in1 => \N__27801\,
            in2 => \_gnd_net_\,
            in3 => \N__29559\,
            lcout => \c0.n3_adj_2226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10686_2_lut_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41873\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_658_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37156\,
            in2 => \_gnd_net_\,
            in3 => \N__37078\,
            lcout => \c0.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_661_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25218\,
            in1 => \N__27025\,
            in2 => \N__33657\,
            in3 => \N__25158\,
            lcout => \c0.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i24_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22497\,
            lcout => \c0.FRAME_MATCHER_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49753\,
            ce => 'H',
            sr => \N__22485\
        );

    \c0.select_219_Select_24_i3_2_lut_3_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41889\,
            in1 => \N__27800\,
            in2 => \_gnd_net_\,
            in3 => \N__25159\,
            lcout => \c0.n3_adj_2242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_25_i3_2_lut_3_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27797\,
            in1 => \N__25219\,
            in2 => \_gnd_net_\,
            in3 => \N__41890\,
            lcout => \c0.n3_adj_2240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_28_i3_2_lut_3_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41888\,
            in1 => \N__27799\,
            in2 => \_gnd_net_\,
            in3 => \N__27026\,
            lcout => \c0.n3_adj_2234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_30_i3_2_lut_3_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27798\,
            in1 => \N__33655\,
            in2 => \_gnd_net_\,
            in3 => \N__41891\,
            lcout => \c0.n3_adj_2230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_4_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__35492\,
            in1 => \N__33444\,
            in2 => \N__35766\,
            in3 => \N__35832\,
            lcout => \c0.n10009\,
            ltout => \c0.n10009_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_588_LC_6_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__37185\,
            in1 => \_gnd_net_\,
            in2 => \N__22440\,
            in3 => \N__41887\,
            lcout => \c0.n3_adj_2181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i18_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22425\,
            in2 => \_gnd_net_\,
            in3 => \N__33187\,
            lcout => \c0.FRAME_MATCHER_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49766\,
            ce => 'H',
            sr => \N__25449\
        );

    \c0.FRAME_MATCHER_i_i27_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22707\,
            lcout => \c0.FRAME_MATCHER_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49778\,
            ce => 'H',
            sr => \N__22659\
        );

    \c0.FRAME_MATCHER_i_i9_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33234\,
            in2 => \_gnd_net_\,
            in3 => \N__22644\,
            lcout => \c0.FRAME_MATCHER_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49788\,
            ce => 'H',
            sr => \N__22599\
        );

    \c0.rx.i15081_4_lut_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__31891\,
            in1 => \N__31853\,
            in2 => \N__31695\,
            in3 => \N__31939\,
            lcout => \c0.rx.n17636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15113_3_lut_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__22853\,
            in1 => \N__25508\,
            in2 => \_gnd_net_\,
            in3 => \N__45263\,
            lcout => n17707,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22575\,
            in1 => \N__22560\,
            in2 => \N__22545\,
            in3 => \N__22527\,
            lcout => \c0.rx.n17022\,
            ltout => \c0.rx.n17022_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_4_lut_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__31719\,
            in1 => \N__31937\,
            in2 => \N__22521\,
            in3 => \N__31774\,
            lcout => \c0.rx.r_SM_Main_2_N_2094_0\,
            ltout => \c0.rx.r_SM_Main_2_N_2094_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14604_2_lut_3_lut_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__31938\,
            in1 => \_gnd_net_\,
            in2 => \N__22518\,
            in3 => \N__45261\,
            lcout => OPEN,
            ltout => \c0.rx.n17380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15000_4_lut_LC_6_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010101"
        )
    port map (
            in0 => \N__25507\,
            in1 => \N__31691\,
            in2 => \N__22515\,
            in3 => \N__31890\,
            lcout => \c0.rx.n17635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_adj_395_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45262\,
            in2 => \_gnd_net_\,
            in3 => \N__22852\,
            lcout => \c0.rx.n6_adj_2130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__6__2279_LC_6_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39030\,
            in1 => \N__29679\,
            in2 => \_gnd_net_\,
            in3 => \N__26973\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__22833\,
            in1 => \N__32388\,
            in2 => \N__22827\,
            in3 => \N__32260\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49659\,
            ce => \N__24264\,
            sr => \_gnd_net_\
        );

    \c0.i15080_3_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__39264\,
            in1 => \N__28612\,
            in2 => \_gnd_net_\,
            in3 => \N__28901\,
            lcout => \c0.n17620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_15415_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__22794\,
            in1 => \N__25729\,
            in2 => \N__22782\,
            in3 => \N__25771\,
            lcout => OPEN,
            ltout => \c0.tx2.n18082_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n18082_bdd_4_lut_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__25772\,
            in1 => \N__22764\,
            in2 => \N__22749\,
            in3 => \N__22746\,
            lcout => OPEN,
            ltout => \c0.tx2.n18085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i11130210_i1_3_lut_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22868\,
            in1 => \_gnd_net_\,
            in2 => \N__22731\,
            in3 => \N__22728\,
            lcout => OPEN,
            ltout => \c0.tx2.o_Tx_Serial_N_2062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26751\,
            in2 => \N__22722\,
            in3 => \N__25936\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25730\,
            in1 => \N__22867\,
            in2 => \_gnd_net_\,
            in3 => \N__25773\,
            lcout => \c0.tx2.n13614\,
            ltout => \c0.tx2.n13614_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5661_4_lut_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26752\,
            in1 => \N__35610\,
            in2 => \N__23064\,
            in3 => \N__25983\,
            lcout => n8191,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__25734\,
            in1 => \N__24673\,
            in2 => \_gnd_net_\,
            in3 => \N__22880\,
            lcout => \r_Bit_Index_0_adj_2442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15074_3_lut_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__28934\,
            in1 => \N__28448\,
            in2 => \_gnd_net_\,
            in3 => \N__40286\,
            lcout => \c0.n17587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__25735\,
            in1 => \N__24674\,
            in2 => \N__25792\,
            in3 => \N__22881\,
            lcout => \r_Bit_Index_1_adj_2441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_612_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39259\,
            in2 => \_gnd_net_\,
            in3 => \N__34710\,
            lcout => \c0.n17107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15326_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__28447\,
            in1 => \N__24527\,
            in2 => \N__23023\,
            in3 => \N__28933\,
            lcout => OPEN,
            ltout => \c0.n18118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18118_bdd_4_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__28449\,
            in2 => \N__22941\,
            in3 => \N__22938\,
            lcout => \c0.n18121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i14643_3_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__26746\,
            in1 => \N__22890\,
            in2 => \_gnd_net_\,
            in3 => \N__24672\,
            lcout => n10976,
            ltout => \n10976_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000000100000"
        )
    port map (
            in0 => \N__25701\,
            in1 => \N__24675\,
            in2 => \N__22872\,
            in3 => \N__22869\,
            lcout => \r_Bit_Index_2_adj_2440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__28925\,
            in1 => \N__23268\,
            in2 => \N__23388\,
            in3 => \N__28497\,
            lcout => \c0.n6_adj_2142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18064_bdd_4_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__28498\,
            in1 => \N__23337\,
            in2 => \N__24654\,
            in3 => \N__24850\,
            lcout => \c0.n18067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001110"
        )
    port map (
            in0 => \N__23316\,
            in1 => \N__25939\,
            in2 => \N__26848\,
            in3 => \N__25984\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__28924\,
            in1 => \_gnd_net_\,
            in2 => \N__26639\,
            in3 => \N__23307\,
            lcout => \c0.n5_adj_2289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_593_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__26032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23262\,
            lcout => OPEN,
            ltout => \c0.n10413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_653_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24137\,
            in1 => \N__23554\,
            in2 => \N__23211\,
            in3 => \N__23621\,
            lcout => \c0.n17282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15331_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__23180\,
            in1 => \N__28923\,
            in2 => \N__28600\,
            in3 => \N__23136\,
            lcout => \c0.n18124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i100_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30171\,
            in1 => \N__23547\,
            in2 => \_gnd_net_\,
            in3 => \N__26585\,
            lcout => data_out_frame2_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15395_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__28998\,
            in1 => \N__23097\,
            in2 => \N__28601\,
            in3 => \N__23084\,
            lcout => \c0.n18160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_509_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40896\,
            in1 => \N__23762\,
            in2 => \N__23748\,
            in3 => \N__23687\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18016_bdd_4_lut_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__28503\,
            in1 => \N__23931\,
            in2 => \N__23653\,
            in3 => \N__23614\,
            lcout => \c0.n18019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_735_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23503\,
            in1 => \N__23546\,
            in2 => \_gnd_net_\,
            in3 => \N__23475\,
            lcout => \c0.n6_adj_2197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i72_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__26584\,
            in1 => \_gnd_net_\,
            in2 => \N__23483\,
            in3 => \N__29929\,
            lcout => data_out_frame2_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i44_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23504\,
            in1 => \N__31622\,
            in2 => \_gnd_net_\,
            in3 => \N__26586\,
            lcout => data_out_frame2_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18142_bdd_4_lut_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__28499\,
            in1 => \N__23490\,
            in2 => \N__23482\,
            in3 => \N__23454\,
            lcout => \c0.n18145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i114_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30359\,
            in1 => \N__23992\,
            in2 => \_gnd_net_\,
            in3 => \N__26511\,
            lcout => data_out_frame2_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i15179_4_lut_4_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__25934\,
            in1 => \N__26750\,
            in2 => \N__35605\,
            in3 => \N__25968\,
            lcout => n4_adj_2484,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_3_lut_4_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__35595\,
            in1 => \N__26847\,
            in2 => \N__26754\,
            in3 => \N__25935\,
            lcout => \c0.tx2.n9269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i132_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26509\,
            in1 => \N__30170\,
            in2 => \_gnd_net_\,
            in3 => \N__24464\,
            lcout => data_out_frame2_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_511_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24129\,
            lcout => \c0.n10456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i86_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26510\,
            in1 => \N__31095\,
            in2 => \_gnd_net_\,
            in3 => \N__24063\,
            lcout => data_out_frame2_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i92_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30716\,
            in1 => \N__24031\,
            in2 => \_gnd_net_\,
            in3 => \N__26512\,
            lcout => data_out_frame2_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i117_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__26508\,
            in1 => \_gnd_net_\,
            in2 => \N__31155\,
            in3 => \N__24778\,
            lcout => data_out_frame2_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_15245_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__23985\,
            in1 => \N__28493\,
            in2 => \N__29066\,
            in3 => \N__23964\,
            lcout => \c0.n18016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_681_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24315\,
            in1 => \N__23910\,
            in2 => \_gnd_net_\,
            in3 => \N__24357\,
            lcout => \c0.n17098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28997\,
            in1 => \N__23852\,
            in2 => \_gnd_net_\,
            in3 => \N__23819\,
            lcout => \c0.n5_adj_2290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_429_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24774\,
            in2 => \_gnd_net_\,
            in3 => \N__24749\,
            lcout => \c0.n17276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i14635_3_lut_4_lut_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__25940\,
            in1 => \N__26840\,
            in2 => \N__26753\,
            in3 => \N__25962\,
            lcout => n17412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_474_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24651\,
            in1 => \N__24609\,
            in2 => \N__27657\,
            in3 => \N__24597\,
            lcout => \c0.n17123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_606_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26042\,
            in2 => \_gnd_net_\,
            in3 => \N__24525\,
            lcout => \c0.n10434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_533_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24471\,
            in2 => \_gnd_net_\,
            in3 => \N__24435\,
            lcout => \c0.n10482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_584_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24308\,
            lcout => \c0.n10513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_514_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42192\,
            in1 => \N__45495\,
            in2 => \N__46647\,
            in3 => \N__48883\,
            lcout => \c0.n17110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_12_i3_2_lut_3_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27834\,
            in1 => \N__25866\,
            in2 => \_gnd_net_\,
            in3 => \N__41765\,
            lcout => \c0.n3_adj_2268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__2__2267_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39221\,
            in1 => \N__36881\,
            in2 => \_gnd_net_\,
            in3 => \N__38967\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_597_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27579\,
            in1 => \N__24936\,
            in2 => \N__24869\,
            in3 => \N__24851\,
            lcout => \c0.n17_adj_2321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__6__2271_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39220\,
            in1 => \N__35094\,
            in2 => \_gnd_net_\,
            in3 => \N__26962\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i19_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44990\,
            in1 => \N__44777\,
            in2 => \N__27430\,
            in3 => \N__44602\,
            lcout => \c0.FRAME_MATCHER_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49722\,
            ce => 'H',
            sr => \N__27408\
        );

    \c0.FRAME_MATCHER_state_i12_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__27347\,
            in1 => \N__44991\,
            in2 => \N__44618\,
            in3 => \N__44799\,
            lcout => \c0.FRAME_MATCHER_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49732\,
            ce => 'H',
            sr => \N__27333\
        );

    \c0.i1_2_lut_adj_410_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33322\,
            in2 => \_gnd_net_\,
            in3 => \N__27346\,
            lcout => OPEN,
            ltout => \c0.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29609\,
            in1 => \N__27323\,
            in2 => \N__24786\,
            in3 => \N__27391\,
            lcout => \c0.n51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15142_3_lut_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__48421\,
            in1 => \N__42492\,
            in2 => \_gnd_net_\,
            in3 => \N__44287\,
            lcout => \c0.n17574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15001_3_lut_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__48419\,
            in1 => \N__47133\,
            in2 => \_gnd_net_\,
            in3 => \N__49109\,
            lcout => \c0.n17643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15002_3_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__49110\,
            in1 => \N__48420\,
            in2 => \_gnd_net_\,
            in3 => \N__44286\,
            lcout => \c0.n17647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i8_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44992\,
            in1 => \N__44800\,
            in2 => \N__33332\,
            in3 => \N__44610\,
            lcout => \c0.FRAME_MATCHER_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49743\,
            ce => 'H',
            sr => \N__33306\
        );

    \c0.i10662_2_lut_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25299\,
            in2 => \_gnd_net_\,
            in3 => \N__41836\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10663_2_lut_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25220\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10664_2_lut_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25169\,
            in2 => \_gnd_net_\,
            in3 => \N__41838\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10665_2_lut_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25125\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10668_2_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41840\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10669_2_lut_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25007\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10672_2_lut_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27889\,
            in2 => \_gnd_net_\,
            in3 => \N__41842\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i5_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45020\,
            in1 => \N__44801\,
            in2 => \N__33469\,
            in3 => \N__44606\,
            lcout => \c0.FRAME_MATCHER_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49754\,
            ce => 'H',
            sr => \N__29475\
        );

    \c0.select_219_Select_18_i3_2_lut_3_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41851\,
            in1 => \_gnd_net_\,
            in2 => \N__25437\,
            in3 => \N__27819\,
            lcout => \c0.n3_adj_2254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10670_2_lut_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25433\,
            in2 => \_gnd_net_\,
            in3 => \N__41849\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_1_i3_2_lut_3_lut_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41852\,
            in1 => \_gnd_net_\,
            in2 => \N__32884\,
            in3 => \N__27817\,
            lcout => \c0.n3_adj_2288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10687_2_lut_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32873\,
            in2 => \_gnd_net_\,
            in3 => \N__41850\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_22_i3_2_lut_3_lut_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41853\,
            in1 => \_gnd_net_\,
            in2 => \N__25347\,
            in3 => \N__27818\,
            lcout => \c0.n3_adj_2246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10666_2_lut_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25343\,
            in2 => \_gnd_net_\,
            in3 => \N__41848\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_26_i3_2_lut_3_lut_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41854\,
            in1 => \N__27816\,
            in2 => \_gnd_net_\,
            in3 => \N__25298\,
            lcout => \c0.n3_adj_2238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i10_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25242\,
            in2 => \_gnd_net_\,
            in3 => \N__33184\,
            lcout => \c0.FRAME_MATCHER_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49767\,
            ce => 'H',
            sr => \N__28017\
        );

    \c0.FRAME_MATCHER_state_i14_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45021\,
            in1 => \N__44812\,
            in2 => \N__27322\,
            in3 => \N__44615\,
            lcout => \c0.FRAME_MATCHER_state_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49779\,
            ce => 'H',
            sr => \N__27297\
        );

    \c0.tx2.i2615_2_lut_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25793\,
            in2 => \_gnd_net_\,
            in3 => \N__25740\,
            lcout => n5266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43880\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_1_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26853\,
            lcout => n10674,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__1__2199_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__25647\,
            in1 => \N__48089\,
            in2 => \N__50321\,
            in3 => \N__29757\,
            lcout => \c0.data_out_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49789\,
            ce => \N__46933\,
            sr => \_gnd_net_\
        );

    \c0.i15053_2_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48088\,
            lcout => \c0.n17626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i13_4_lut_4_lut_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__31850\,
            in1 => \N__25584\,
            in2 => \N__25509\,
            in3 => \N__25563\,
            lcout => \c0.rx.n10620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i14585_4_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__25561\,
            in1 => \N__25503\,
            in2 => \N__25591\,
            in3 => \N__31849\,
            lcout => n17361,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_3_lut_4_lut_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__31775\,
            in1 => \N__31735\,
            in2 => \N__31952\,
            in3 => \N__31895\,
            lcout => \c0.rx.r_SM_Main_2_N_2088_2\,
            ltout => \c0.rx.r_SM_Main_2_N_2088_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_4_lut_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__25562\,
            in1 => \N__31848\,
            in2 => \N__25512\,
            in3 => \N__25502\,
            lcout => \c0.rx.n10158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i12_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25884\,
            in2 => \_gnd_net_\,
            in3 => \N__33232\,
            lcout => \c0.FRAME_MATCHER_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49799\,
            ce => 'H',
            sr => \N__25833\
        );

    \c0.FRAME_MATCHER_state_i20_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__45032\,
            in1 => \N__44813\,
            in2 => \N__44619\,
            in3 => \N__29608\,
            lcout => \c0.FRAME_MATCHER_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \N__29586\
        );

    \c0.byte_transmit_counter2_i4_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__25806\,
            in1 => \N__32234\,
            in2 => \N__39683\,
            in3 => \N__42086\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49676\,
            ce => 'H',
            sr => \N__26922\
        );

    \c0.add_2510_2_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34110\,
            in1 => \N__28783\,
            in2 => \_gnd_net_\,
            in3 => \N__25818\,
            lcout => \c0.n17659\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \c0.n15972\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_3_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34112\,
            in1 => \N__28465\,
            in2 => \_gnd_net_\,
            in3 => \N__25815\,
            lcout => \c0.n17589\,
            ltout => OPEN,
            carryin => \c0.n15972\,
            carryout => \c0.n15973\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_4_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34108\,
            in1 => \N__32109\,
            in2 => \_gnd_net_\,
            in3 => \N__25812\,
            lcout => \c0.n17710\,
            ltout => OPEN,
            carryin => \c0.n15973\,
            carryout => \c0.n15974\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_5_lut_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34113\,
            in1 => \N__32334\,
            in2 => \_gnd_net_\,
            in3 => \N__25809\,
            lcout => \c0.n17711\,
            ltout => OPEN,
            carryin => \c0.n15974\,
            carryout => \c0.n15975\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_6_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34109\,
            in1 => \N__32225\,
            in2 => \_gnd_net_\,
            in3 => \N__25800\,
            lcout => \c0.n17606\,
            ltout => OPEN,
            carryin => \c0.n15975\,
            carryout => \c0.n15976\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_7_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34111\,
            in1 => \N__39623\,
            in2 => \_gnd_net_\,
            in3 => \N__25797\,
            lcout => \c0.n17712\,
            ltout => OPEN,
            carryin => \c0.n15976\,
            carryout => \c0.n15977\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_8_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34106\,
            in1 => \N__34446\,
            in2 => \_gnd_net_\,
            in3 => \N__26670\,
            lcout => \c0.n17713\,
            ltout => OPEN,
            carryin => \c0.n15977\,
            carryout => \c0.n15978\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2510_9_lut_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__34485\,
            in1 => \N__34107\,
            in2 => \_gnd_net_\,
            in3 => \N__26667\,
            lcout => \c0.n17714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i1_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__26652\,
            in1 => \N__28362\,
            in2 => \N__39679\,
            in3 => \N__42084\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49677\,
            ce => 'H',
            sr => \N__28263\
        );

    \c0.i1_2_lut_adj_415_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37186\,
            in2 => \_gnd_net_\,
            in3 => \N__37105\,
            lcout => \c0.n15179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i58_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29817\,
            in1 => \N__26632\,
            in2 => \_gnd_net_\,
            in3 => \N__26612\,
            lcout => data_out_frame2_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__0__2277_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39207\,
            in1 => \N__29140\,
            in2 => \_gnd_net_\,
            in3 => \N__34934\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__25985\,
            in1 => \N__25937\,
            in2 => \N__26741\,
            in3 => \N__26818\,
            lcout => \r_SM_Main_1_adj_2439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i97_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29458\,
            in1 => \N__26022\,
            in2 => \_gnd_net_\,
            in3 => \N__26613\,
            lcout => data_out_frame2_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__25986\,
            in1 => \N__25938\,
            in2 => \N__26740\,
            in3 => \N__26819\,
            lcout => \r_SM_Main_2_adj_2438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_3_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__48425\,
            in1 => \N__48167\,
            in2 => \_gnd_net_\,
            in3 => \N__50315\,
            lcout => n10705,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14597_3_lut_4_lut_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__32514\,
            in1 => \N__34773\,
            in2 => \N__35127\,
            in3 => \N__37398\,
            lcout => \c0.n17373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i50_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39479\,
            in1 => \N__34673\,
            in2 => \_gnd_net_\,
            in3 => \N__32562\,
            lcout => data_in_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110100"
        )
    port map (
            in0 => \N__26826\,
            in1 => \N__26769\,
            in2 => \N__34395\,
            in3 => \N__26720\,
            lcout => tx2_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32563\,
            in1 => \N__39553\,
            in2 => \_gnd_net_\,
            in3 => \N__36992\,
            lcout => data_in_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34550\,
            in1 => \N__36801\,
            in2 => \_gnd_net_\,
            in3 => \N__32561\,
            lcout => data_in_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__2__2283_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39206\,
            in1 => \N__28048\,
            in2 => \_gnd_net_\,
            in3 => \N__38940\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__5__2272_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29180\,
            in1 => \N__29651\,
            in2 => \_gnd_net_\,
            in3 => \N__39211\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__3__2290_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26868\,
            in1 => \N__39095\,
            in2 => \_gnd_net_\,
            in3 => \N__26901\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_657_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26900\,
            in1 => \N__29176\,
            in2 => \N__29154\,
            in3 => \N__29280\,
            lcout => \c0.n17_adj_2370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10774_2_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29328\,
            in2 => \_gnd_net_\,
            in3 => \N__26899\,
            lcout => \c0.n13450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__7__2286_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29329\,
            in1 => \N__39212\,
            in2 => \_gnd_net_\,
            in3 => \N__26880\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__3__2274_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39210\,
            in1 => \N__29213\,
            in2 => \_gnd_net_\,
            in3 => \N__35241\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__3__2282_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29214\,
            in1 => \N__39213\,
            in2 => \_gnd_net_\,
            in3 => \N__26867\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__0__2285_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39209\,
            in1 => \N__29153\,
            in2 => \_gnd_net_\,
            in3 => \N__35051\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_627_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27531\,
            in1 => \N__26943\,
            in2 => \N__35009\,
            in3 => \N__26979\,
            lcout => \c0.n10133\,
            ltout => \c0.n10133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_631_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26889\,
            in3 => \N__27277\,
            lcout => OPEN,
            ltout => \c0.n6_adj_2356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_632_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__26907\,
            in1 => \N__29211\,
            in2 => \N__26886\,
            in3 => \N__29232\,
            lcout => \c0.n10027\,
            ltout => \c0.n10027_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_642_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__35377\,
            in1 => \N__28029\,
            in2 => \N__26883\,
            in3 => \N__29253\,
            lcout => n63_adj_2418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14556_2_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26879\,
            in2 => \_gnd_net_\,
            in3 => \N__26866\,
            lcout => OPEN,
            ltout => \c0.n17331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14633_4_lut_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35050\,
            in1 => \N__27546\,
            in2 => \N__26982\,
            in3 => \N__27516\,
            lcout => \c0.n17410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__4__2281_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39184\,
            in1 => \N__26937\,
            in2 => \_gnd_net_\,
            in3 => \N__29233\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_625_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26963\,
            in1 => \N__35237\,
            in2 => \N__35405\,
            in3 => \N__26935\,
            lcout => \c0.n12_adj_2355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__4__2273_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26936\,
            in1 => \N__39186\,
            in2 => \_gnd_net_\,
            in3 => \N__29733\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14650_4_lut_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000110000"
        )
    port map (
            in0 => \N__36245\,
            in1 => \N__36275\,
            in2 => \N__36174\,
            in3 => \N__36203\,
            lcout => n17427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_414_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32247\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33537\,
            lcout => \c0.n4_adj_2150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__1__2276_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__35401\,
            in1 => \_gnd_net_\,
            in2 => \N__39218\,
            in3 => \N__35010\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_646_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__29731\,
            in1 => \N__26913\,
            in2 => \N__27282\,
            in3 => \N__27566\,
            lcout => \c0.n17_adj_2362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14629_4_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38977\,
            in1 => \N__29730\,
            in2 => \N__27567\,
            in3 => \N__34933\,
            lcout => \c0.n17406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__6__2287_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27281\,
            in1 => \N__39185\,
            in2 => \_gnd_net_\,
            in3 => \N__29712\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i9_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44931\,
            in1 => \N__44776\,
            in2 => \N__33290\,
            in3 => \N__44601\,
            lcout => \c0.FRAME_MATCHER_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49744\,
            ce => 'H',
            sr => \N__33264\
        );

    \c0.i10673_2_lut_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27264\,
            in2 => \_gnd_net_\,
            in3 => \N__41672\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10675_2_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27210\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10677_2_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27159\,
            in2 => \_gnd_net_\,
            in3 => \N__41674\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10681_2_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27099\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_405_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41670\,
            lcout => \c0.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_701_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41671\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27033\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15155_2_lut_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36297\,
            in2 => \_gnd_net_\,
            in3 => \N__47842\,
            lcout => \c0.n17701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27431\,
            in1 => \N__27482\,
            in2 => \N__38070\,
            in3 => \N__27451\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i13_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__27453\,
            in1 => \N__44932\,
            in2 => \N__44603\,
            in3 => \N__44768\,
            lcout => \c0.FRAME_MATCHER_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49755\,
            ce => 'H',
            sr => \N__27441\
        );

    \c0.i1_2_lut_adj_712_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27452\,
            in2 => \_gnd_net_\,
            in3 => \N__40796\,
            lcout => \c0.n8_adj_2332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_723_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27432\,
            lcout => \c0.n8_adj_2328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_705_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27396\,
            in2 => \_gnd_net_\,
            in3 => \N__40793\,
            lcout => \c0.n8_adj_2334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_709_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37299\,
            lcout => \c0.n8_adj_2333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_711_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27351\,
            in2 => \_gnd_net_\,
            in3 => \N__40795\,
            lcout => \c0.n16708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_713_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27324\,
            lcout => \c0.n8_adj_2331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_718_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__41332\,
            in1 => \N__27483\,
            in2 => \N__41427\,
            in3 => \N__41457\,
            lcout => \c0.n16716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_594_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27656\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27606\,
            lcout => \c0.n10459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_398_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__37868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37829\,
            lcout => n10010,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__5__2288_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27515\,
            in1 => \N__39131\,
            in2 => \_gnd_net_\,
            in3 => \N__27562\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__4__2289_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39129\,
            in1 => \N__29241\,
            in2 => \_gnd_net_\,
            in3 => \N__27545\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__2__2291_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28054\,
            in1 => \N__39130\,
            in2 => \_gnd_net_\,
            in3 => \N__27530\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__5__2280_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29181\,
            in1 => \N__39132\,
            in2 => \_gnd_net_\,
            in3 => \N__27514\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i16_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27498\,
            in2 => \_gnd_net_\,
            in3 => \N__33159\,
            lcout => \c0.FRAME_MATCHER_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49780\,
            ce => 'H',
            sr => \N__27687\
        );

    \c0.FRAME_MATCHER_state_i4_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__44986\,
            in1 => \N__44798\,
            in2 => \N__44616\,
            in3 => \N__27481\,
            lcout => \c0.FRAME_MATCHER_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49790\,
            ce => 'H',
            sr => \N__27462\
        );

    \c0.i2_3_lut_adj_628_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__28055\,
            in1 => \N__35092\,
            in2 => \_gnd_net_\,
            in3 => \N__35385\,
            lcout => \c0.n10141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14611_2_lut_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35093\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28056\,
            lcout => \c0.n17388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_10_i3_2_lut_3_lut_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41845\,
            in1 => \N__27821\,
            in2 => \_gnd_net_\,
            in3 => \N__28001\,
            lcout => \c0.n3_adj_2272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10678_2_lut_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28000\,
            in2 => \_gnd_net_\,
            in3 => \N__41844\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_14_i3_2_lut_3_lut_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41846\,
            in1 => \_gnd_net_\,
            in2 => \N__27942\,
            in3 => \N__27820\,
            lcout => \c0.n3_adj_2264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10674_2_lut_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27937\,
            in2 => \_gnd_net_\,
            in3 => \N__41843\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_219_Select_16_i3_2_lut_3_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__41847\,
            in1 => \N__27873\,
            in2 => \_gnd_net_\,
            in3 => \N__27822\,
            lcout => \c0.n3_adj_2259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i0_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27675\,
            in2 => \_gnd_net_\,
            in3 => \N__27669\,
            lcout => n26_adj_2423,
            ltout => OPEN,
            carryin => \bfn_9_29_0_\,
            carryout => n16041,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i1_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27666\,
            in2 => \_gnd_net_\,
            in3 => \N__27660\,
            lcout => n25_adj_2424,
            ltout => OPEN,
            carryin => n16041,
            carryout => n16042,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i2_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28137\,
            in2 => \_gnd_net_\,
            in3 => \N__28131\,
            lcout => n24,
            ltout => OPEN,
            carryin => n16042,
            carryout => n16043,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i3_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28128\,
            in2 => \_gnd_net_\,
            in3 => \N__28122\,
            lcout => n23_adj_2425,
            ltout => OPEN,
            carryin => n16043,
            carryout => n16044,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i4_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28119\,
            in2 => \_gnd_net_\,
            in3 => \N__28113\,
            lcout => n22_adj_2426,
            ltout => OPEN,
            carryin => n16044,
            carryout => n16045,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i5_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28110\,
            in2 => \_gnd_net_\,
            in3 => \N__28104\,
            lcout => n21,
            ltout => OPEN,
            carryin => n16045,
            carryout => n16046,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i6_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28101\,
            in2 => \_gnd_net_\,
            in3 => \N__28095\,
            lcout => n20,
            ltout => OPEN,
            carryin => n16046,
            carryout => n16047,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i7_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28092\,
            in2 => \_gnd_net_\,
            in3 => \N__28086\,
            lcout => n19,
            ltout => OPEN,
            carryin => n16047,
            carryout => n16048,
            clk => \N__49800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i8_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28083\,
            in2 => \_gnd_net_\,
            in3 => \N__28077\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_9_30_0_\,
            carryout => n16049,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i9_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28074\,
            in2 => \_gnd_net_\,
            in3 => \N__28068\,
            lcout => n17,
            ltout => OPEN,
            carryin => n16049,
            carryout => n16050,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i10_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28065\,
            in2 => \_gnd_net_\,
            in3 => \N__28059\,
            lcout => n16,
            ltout => OPEN,
            carryin => n16050,
            carryout => n16051,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i11_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28209\,
            in2 => \_gnd_net_\,
            in3 => \N__28203\,
            lcout => n15,
            ltout => OPEN,
            carryin => n16051,
            carryout => n16052,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i12_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28200\,
            in2 => \_gnd_net_\,
            in3 => \N__28194\,
            lcout => n14,
            ltout => OPEN,
            carryin => n16052,
            carryout => n16053,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i13_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28191\,
            in2 => \_gnd_net_\,
            in3 => \N__28185\,
            lcout => n13,
            ltout => OPEN,
            carryin => n16053,
            carryout => n16054,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i14_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28182\,
            in2 => \_gnd_net_\,
            in3 => \N__28176\,
            lcout => n12,
            ltout => OPEN,
            carryin => n16054,
            carryout => n16055,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i15_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28173\,
            in2 => \_gnd_net_\,
            in3 => \N__28167\,
            lcout => n11,
            ltout => OPEN,
            carryin => n16055,
            carryout => n16056,
            clk => \N__49807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i16_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28164\,
            in2 => \_gnd_net_\,
            in3 => \N__28158\,
            lcout => n10_adj_2420,
            ltout => OPEN,
            carryin => \bfn_9_31_0_\,
            carryout => n16057,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i17_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28155\,
            in2 => \_gnd_net_\,
            in3 => \N__28149\,
            lcout => n9_adj_2421,
            ltout => OPEN,
            carryin => n16057,
            carryout => n16058,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i18_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28146\,
            in2 => \_gnd_net_\,
            in3 => \N__28140\,
            lcout => n8_adj_2412,
            ltout => OPEN,
            carryin => n16058,
            carryout => n16059,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i19_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28248\,
            in2 => \_gnd_net_\,
            in3 => \N__28242\,
            lcout => n7,
            ltout => OPEN,
            carryin => n16059,
            carryout => n16060,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i20_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28239\,
            in2 => \_gnd_net_\,
            in3 => \N__28233\,
            lcout => n6_adj_2429,
            ltout => OPEN,
            carryin => n16060,
            carryout => n16061,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i21_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36154\,
            in2 => \_gnd_net_\,
            in3 => \N__28230\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n16061,
            carryout => n16062,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i22_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36190\,
            in2 => \_gnd_net_\,
            in3 => \N__28227\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n16062,
            carryout => n16063,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i23_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36226\,
            in2 => \_gnd_net_\,
            in3 => \N__28224\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n16063,
            carryout => n16064,
            clk => \N__49815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i24_LC_9_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36257\,
            in2 => \_gnd_net_\,
            in3 => \N__28221\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_9_32_0_\,
            carryout => n16065,
            clk => \N__49823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2360__i25_LC_9_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36005\,
            in2 => \_gnd_net_\,
            in3 => \N__28218\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i3_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__28215\,
            in1 => \N__32363\,
            in2 => \N__39678\,
            in3 => \N__42096\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49679\,
            ce => 'H',
            sr => \N__29079\
        );

    \c0.i10493_2_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35606\,
            in2 => \_gnd_net_\,
            in3 => \N__34398\,
            lcout => \c0.n11867\,
            ltout => \c0.n11867_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i0_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__29097\,
            in1 => \N__28818\,
            in2 => \N__29091\,
            in3 => \N__42093\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49668\,
            ce => 'H',
            sr => \N__29088\
        );

    \c0.i1_2_lut_adj_763_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33535\,
            lcout => \c0.n4_adj_2187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_412_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__33534\,
            in1 => \N__32362\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n4_adj_2152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15170_3_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__37580\,
            in1 => \N__28360\,
            in2 => \_gnd_net_\,
            in3 => \N__28816\,
            lcout => \c0.n17761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i47_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__40421\,
            in1 => \N__32492\,
            in2 => \N__39554\,
            in3 => \N__32706\,
            lcout => \c0.data_in_frame_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i31_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__28257\,
            in1 => \N__39545\,
            in2 => \N__40623\,
            in3 => \N__39394\,
            lcout => \c0.data_in_frame_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_408_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28361\,
            in2 => \_gnd_net_\,
            in3 => \N__33536\,
            lcout => \c0.n4_adj_2155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__40606\,
            in1 => \N__35276\,
            in2 => \N__38899\,
            in3 => \N__40422\,
            lcout => \c0.data_in_frame_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_562_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__28256\,
            in1 => \N__37010\,
            in2 => \N__29301\,
            in3 => \N__34832\,
            lcout => \c0.n19_adj_2303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__37983\,
            in1 => \N__45260\,
            in2 => \N__35297\,
            in3 => \N__36710\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35287\,
            in1 => \N__32936\,
            in2 => \_gnd_net_\,
            in3 => \N__32564\,
            lcout => data_in_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i32_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__40619\,
            in1 => \N__40504\,
            in2 => \N__37523\,
            in3 => \N__39386\,
            lcout => \c0.data_in_frame_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_574_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__29108\,
            in1 => \N__32765\,
            in2 => \N__39288\,
            in3 => \N__32619\,
            lcout => OPEN,
            ltout => \c0.n15_adj_2310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_595_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110111"
        )
    port map (
            in0 => \N__34161\,
            in1 => \N__36906\,
            in2 => \N__29112\,
            in3 => \N__37471\,
            lcout => \c0.n22_adj_2319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__5__2264_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36675\,
            in1 => \N__39208\,
            in2 => \_gnd_net_\,
            in3 => \N__29646\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i28_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__29109\,
            in1 => \N__35288\,
            in2 => \N__40626\,
            in3 => \N__39385\,
            lcout => \c0.data_in_frame_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__40600\,
            in1 => \N__34521\,
            in2 => \N__36689\,
            in3 => \N__40419\,
            lcout => \c0.data_in_frame_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i45_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__40418\,
            in1 => \N__38849\,
            in2 => \N__45133\,
            in3 => \N__32680\,
            lcout => \c0.data_in_frame_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36877\,
            in1 => \N__34343\,
            in2 => \_gnd_net_\,
            in3 => \N__32559\,
            lcout => data_in_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_696_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__34767\,
            in1 => \N__37397\,
            in2 => \_gnd_net_\,
            in3 => \N__34574\,
            lcout => \c0.n2137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i42_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__34655\,
            in1 => \N__39476\,
            in2 => \N__32695\,
            in3 => \N__40420\,
            lcout => \c0.data_in_frame_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32560\,
            in1 => \N__36680\,
            in2 => \_gnd_net_\,
            in3 => \N__34253\,
            lcout => data_in_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_616_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__37113\,
            in1 => \N__37187\,
            in2 => \_gnd_net_\,
            in3 => \N__39362\,
            lcout => n17075,
            ltout => \n17075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40505\,
            in1 => \_gnd_net_\,
            in2 => \N__29184\,
            in3 => \N__34974\,
            lcout => data_in_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__7__2270_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39217\,
            in1 => \N__29392\,
            in2 => \_gnd_net_\,
            in3 => \N__32921\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14623_3_lut_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__29391\,
            in1 => \N__29175\,
            in2 => \_gnd_net_\,
            in3 => \N__29278\,
            lcout => OPEN,
            ltout => \c0.n17400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_637_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__29149\,
            in1 => \N__38932\,
            in2 => \N__29124\,
            in3 => \N__32898\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_640_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__29647\,
            in1 => \N__29710\,
            in2 => \N__29121\,
            in3 => \N__29118\,
            lcout => \c0.n10136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__7__2278_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39216\,
            in1 => \N__29333\,
            in2 => \_gnd_net_\,
            in3 => \N__29393\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i29_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__40599\,
            in1 => \N__45134\,
            in2 => \N__29300\,
            in3 => \N__39361\,
            lcout => \c0.data_in_frame_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__7__2262_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40503\,
            in1 => \N__39215\,
            in2 => \_gnd_net_\,
            in3 => \N__32920\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__1__2292_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39214\,
            in1 => \N__35384\,
            in2 => \_gnd_net_\,
            in3 => \N__29279\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_3_lut_4_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__36091\,
            in1 => \N__44862\,
            in2 => \N__41976\,
            in3 => \N__41700\,
            lcout => OPEN,
            ltout => \c0.n7_adj_2384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i3_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33488\,
            in1 => \N__33669\,
            in2 => \N__29265\,
            in3 => \N__35757\,
            lcout => \c0.FRAME_MATCHER_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49724\,
            ce => 'H',
            sr => \N__29262\
        );

    \c0.i1_2_lut_adj_700_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33487\,
            in2 => \_gnd_net_\,
            in3 => \N__41297\,
            lcout => \c0.n6_adj_2336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33384\,
            in1 => \N__41606\,
            in2 => \N__33740\,
            in3 => \N__33359\,
            lcout => \c0.n9369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_645_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__29252\,
            in1 => \N__38978\,
            in2 => \N__29240\,
            in3 => \N__34935\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_647_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__29212\,
            in1 => \N__29375\,
            in2 => \N__29193\,
            in3 => \N__29190\,
            lcout => n63,
            ltout => \n63_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_793_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__36090\,
            in1 => \N__33383\,
            in2 => \N__29400\,
            in3 => \N__33732\,
            lcout => \FRAME_MATCHER_state_31_N_1406_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_649_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38939\,
            in1 => \N__29397\,
            in2 => \N__29376\,
            in3 => \N__29355\,
            lcout => OPEN,
            ltout => \c0.n16_adj_2366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_670_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__29622\,
            in1 => \N__29349\,
            in2 => \N__29337\,
            in3 => \N__29334\,
            lcout => n63_adj_2428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41268\,
            in1 => \N__33280\,
            in2 => \N__41235\,
            in3 => \N__37335\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_638_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33354\,
            in1 => \N__33728\,
            in2 => \_gnd_net_\,
            in3 => \N__33380\,
            lcout => n9378,
            ltout => \n9378_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_618_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33554\,
            in2 => \N__29310\,
            in3 => \N__33012\,
            lcout => \c0.n47_adj_2347\,
            ltout => \c0.n47_adj_2347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_762_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__35941\,
            in1 => \N__35892\,
            in2 => \N__29307\,
            in3 => \N__41669\,
            lcout => \c0.n17069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_673_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__33381\,
            in1 => \_gnd_net_\,
            in2 => \N__33739\,
            in3 => \N__33355\,
            lcout => \c0.n13146\,
            ltout => \c0.n13146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__35940\,
            in1 => \_gnd_net_\,
            in2 => \N__29304\,
            in3 => \N__35891\,
            lcout => \c0.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__4__2265_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45120\,
            in1 => \N__39190\,
            in2 => \_gnd_net_\,
            in3 => \N__29732\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14625_4_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29711\,
            in1 => \N__35034\,
            in2 => \N__29655\,
            in3 => \N__32922\,
            lcout => \c0.n17402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_725_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29616\,
            in2 => \_gnd_net_\,
            in3 => \N__40792\,
            lcout => \c0.n8_adj_2327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10589_4_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__32880\,
            in1 => \N__37174\,
            in2 => \N__29571\,
            in3 => \N__29508\,
            lcout => n2061,
            ltout => \n2061_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29496\,
            in3 => \N__41668\,
            lcout => \c0.n9334\,
            ltout => \c0.n9334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_739_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__41362\,
            in1 => \N__29493\,
            in2 => \N__29487\,
            in3 => \N__29484\,
            lcout => \c0.n15821\,
            ltout => \c0.n15821_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_704_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29478\,
            in3 => \N__33471\,
            lcout => \c0.n8_adj_2335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i0_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29460\,
            in2 => \N__38018\,
            in3 => \_gnd_net_\,
            lcout => rand_setpoint_0,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => n16010,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i1_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30279\,
            in2 => \N__36410\,
            in3 => \N__30219\,
            lcout => rand_setpoint_1,
            ltout => OPEN,
            carryin => n16010,
            carryout => n16011,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i2_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30216\,
            in2 => \N__33831\,
            in3 => \N__30174\,
            lcout => rand_setpoint_2,
            ltout => OPEN,
            carryin => n16011,
            carryout => n16012,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i3_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30162\,
            in2 => \N__33815\,
            in3 => \N__30114\,
            lcout => rand_setpoint_3,
            ltout => OPEN,
            carryin => n16012,
            carryout => n16013,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i4_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30111\,
            in2 => \N__36338\,
            in3 => \N__30057\,
            lcout => rand_setpoint_4,
            ltout => OPEN,
            carryin => n16013,
            carryout => n16014,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i5_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30053\,
            in2 => \N__43736\,
            in3 => \N__29997\,
            lcout => rand_setpoint_5,
            ltout => OPEN,
            carryin => n16014,
            carryout => n16015,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i6_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29994\,
            in2 => \N__36314\,
            in3 => \N__29934\,
            lcout => rand_setpoint_6,
            ltout => OPEN,
            carryin => n16015,
            carryout => n16016,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i7_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29930\,
            in2 => \N__38153\,
            in3 => \N__29877\,
            lcout => rand_setpoint_7,
            ltout => OPEN,
            carryin => n16016,
            carryout => n16017,
            clk => \N__49756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i8_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29873\,
            in2 => \N__42167\,
            in3 => \N__29820\,
            lcout => rand_setpoint_8,
            ltout => OPEN,
            carryin => \bfn_10_26_0_\,
            carryout => n16018,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i9_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29816\,
            in2 => \N__29753\,
            in3 => \N__29736\,
            lcout => rand_setpoint_9,
            ltout => OPEN,
            carryin => n16018,
            carryout => n16019,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i10_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30779\,
            in2 => \N__31973\,
            in3 => \N__30720\,
            lcout => rand_setpoint_10,
            ltout => OPEN,
            carryin => n16019,
            carryout => n16020,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i11_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30707\,
            in2 => \N__32012\,
            in3 => \N__30660\,
            lcout => rand_setpoint_11,
            ltout => OPEN,
            carryin => n16020,
            carryout => n16021,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i12_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30655\,
            in2 => \N__33983\,
            in3 => \N__30603\,
            lcout => rand_setpoint_12,
            ltout => OPEN,
            carryin => n16021,
            carryout => n16022,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i13_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30600\,
            in2 => \N__43646\,
            in3 => \N__30540\,
            lcout => rand_setpoint_13,
            ltout => OPEN,
            carryin => n16022,
            carryout => n16023,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i14_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30535\,
            in2 => \N__34067\,
            in3 => \N__30471\,
            lcout => rand_setpoint_14,
            ltout => OPEN,
            carryin => n16023,
            carryout => n16024,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i15_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30468\,
            in2 => \N__38099\,
            in3 => \N__30417\,
            lcout => rand_setpoint_15,
            ltout => OPEN,
            carryin => n16024,
            carryout => n16025,
            clk => \N__49769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i16_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30414\,
            in2 => \N__38120\,
            in3 => \N__30366\,
            lcout => rand_setpoint_16,
            ltout => OPEN,
            carryin => \bfn_10_27_0_\,
            carryout => n16026,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i17_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30355\,
            in2 => \N__30299\,
            in3 => \N__30282\,
            lcout => rand_setpoint_17,
            ltout => OPEN,
            carryin => n16026,
            carryout => n16027,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i18_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31268\,
            in2 => \N__33882\,
            in3 => \N__31212\,
            lcout => rand_setpoint_18,
            ltout => OPEN,
            carryin => n16027,
            carryout => n16028,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i19_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31201\,
            in2 => \N__33900\,
            in3 => \N__31158\,
            lcout => rand_setpoint_19,
            ltout => OPEN,
            carryin => n16028,
            carryout => n16029,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i20_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31154\,
            in2 => \N__33945\,
            in3 => \N__31098\,
            lcout => rand_setpoint_20,
            ltout => OPEN,
            carryin => n16029,
            carryout => n16030,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i21_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31094\,
            in2 => \N__33864\,
            in3 => \N__31035\,
            lcout => rand_setpoint_21,
            ltout => OPEN,
            carryin => n16030,
            carryout => n16031,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i22_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31031\,
            in2 => \N__33930\,
            in3 => \N__30978\,
            lcout => rand_setpoint_22,
            ltout => OPEN,
            carryin => n16031,
            carryout => n16032,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i23_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30974\,
            in2 => \N__33764\,
            in3 => \N__30924\,
            lcout => rand_setpoint_23,
            ltout => OPEN,
            carryin => n16032,
            carryout => n16033,
            clk => \N__49781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i24_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30920\,
            in2 => \N__30863\,
            in3 => \N__30846\,
            lcout => rand_setpoint_24,
            ltout => OPEN,
            carryin => \bfn_10_28_0_\,
            carryout => n16034,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i25_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30838\,
            in2 => \N__47894\,
            in3 => \N__30786\,
            lcout => rand_setpoint_25,
            ltout => OPEN,
            carryin => n16034,
            carryout => n16035,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i26_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31677\,
            in2 => \N__31319\,
            in3 => \N__31626\,
            lcout => rand_setpoint_26,
            ltout => OPEN,
            carryin => n16035,
            carryout => n16036,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i27_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31614\,
            in2 => \N__31287\,
            in3 => \N__31569\,
            lcout => rand_setpoint_27,
            ltout => OPEN,
            carryin => n16036,
            carryout => n16037,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i28_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31566\,
            in2 => \N__32031\,
            in3 => \N__31518\,
            lcout => rand_setpoint_28,
            ltout => OPEN,
            carryin => n16037,
            carryout => n16038,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i29_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31513\,
            in2 => \N__31302\,
            in3 => \N__31461\,
            lcout => rand_setpoint_29,
            ltout => OPEN,
            carryin => n16038,
            carryout => n16039,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i30_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31454\,
            in2 => \N__42293\,
            in3 => \N__31404\,
            lcout => rand_setpoint_30,
            ltout => OPEN,
            carryin => n16039,
            carryout => n16040,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_setpoint_2359__i31_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31401\,
            in1 => \N__31334\,
            in2 => \_gnd_net_\,
            in3 => \N__31347\,
            lcout => rand_setpoint_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__2__2214_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__48153\,
            in1 => \N__31320\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49801\,
            ce => \N__50575\,
            sr => \N__42806\
        );

    \c0.data_out_5__5__2211_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48152\,
            in2 => \_gnd_net_\,
            in3 => \N__31301\,
            lcout => \c0.data_out_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49801\,
            ce => \N__50575\,
            sr => \N__42806\
        );

    \c0.data_out_5__3__2213_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48151\,
            in2 => \_gnd_net_\,
            in3 => \N__31286\,
            lcout => \c0.data_out_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49801\,
            ce => \N__50575\,
            sr => \N__42806\
        );

    \c0.data_out_5__4__2212_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__48154\,
            in1 => \N__32030\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49801\,
            ce => \N__50575\,
            sr => \N__42806\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47156\,
            in1 => \N__46695\,
            in2 => \_gnd_net_\,
            in3 => \N__47819\,
            lcout => \c0.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14998_2_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32016\,
            in2 => \_gnd_net_\,
            in3 => \N__48130\,
            lcout => \c0.n17585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14993_2_lut_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31977\,
            lcout => OPEN,
            ltout => \c0.n17583_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__2__2198_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__50261\,
            in1 => \N__48409\,
            in2 => \N__31956\,
            in3 => \N__47321\,
            lcout => \c0.data_out_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49808\,
            ce => \N__46923\,
            sr => \_gnd_net_\
        );

    \c0.i15230_2_lut_3_lut_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__48131\,
            in1 => \N__48405\,
            in2 => \_gnd_net_\,
            in3 => \N__50260\,
            lcout => \c0.n10594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__31737\,
            in1 => \N__31953\,
            in2 => \N__31785\,
            in3 => \N__31899\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49816\,
            ce => 'H',
            sr => \N__31800\
        );

    \c0.rx.i1_2_lut_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31781\,
            in2 => \_gnd_net_\,
            in3 => \N__31736\,
            lcout => \c0.rx.n17080\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47818\,
            in1 => \N__34172\,
            in2 => \_gnd_net_\,
            in3 => \N__34214\,
            lcout => \c0.n2_adj_2145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15122_2_lut_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34226\,
            in2 => \_gnd_net_\,
            in3 => \N__47817\,
            lcout => \c0.n17622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10610_3_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__32333\,
            in1 => \N__32235\,
            in2 => \_gnd_net_\,
            in3 => \N__32069\,
            lcout => \c0.n13284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i2_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32071\,
            in1 => \N__32187\,
            in2 => \N__39693\,
            in3 => \N__42085\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49690\,
            ce => 'H',
            sr => \N__32049\
        );

    \c0.i1_2_lut_adj_411_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32070\,
            in2 => \_gnd_net_\,
            in3 => \N__33519\,
            lcout => \c0.n4_adj_2154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_605_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33521\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34441\,
            lcout => \c0.n4_adj_2325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_679_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34476\,
            in2 => \_gnd_net_\,
            in3 => \N__33522\,
            lcout => \c0.n4_adj_2345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_465_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39624\,
            lcout => \c0.n4_adj_2147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_585_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32474\,
            in1 => \N__38822\,
            in2 => \_gnd_net_\,
            in3 => \N__39994\,
            lcout => \c0.n16475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i48_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__32708\,
            in1 => \N__34628\,
            in2 => \N__40509\,
            in3 => \N__40429\,
            lcout => \c0.data_in_frame_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i46_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__32707\,
            in1 => \N__32601\,
            in2 => \N__36690\,
            in3 => \N__40428\,
            lcout => \c0.data_in_frame_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1010_2_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32751\,
            in2 => \_gnd_net_\,
            in3 => \N__34896\,
            lcout => \c0.n2122\,
            ltout => \c0.n2122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_464_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__32506\,
            in1 => \N__35324\,
            in2 => \N__32517\,
            in3 => \N__32766\,
            lcout => \c0.n20_adj_2195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__37736\,
            in1 => \N__36687\,
            in2 => \N__39396\,
            in3 => \N__32507\,
            lcout => \c0.data_in_frame_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__38823\,
            in1 => \N__36863\,
            in2 => \N__40625\,
            in3 => \N__40427\,
            lcout => \c0.data_in_frame_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i43_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__32702\,
            in1 => \N__40050\,
            in2 => \N__36882\,
            in3 => \N__40424\,
            lcout => \c0.data_in_frame_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_611_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011111111"
        )
    port map (
            in0 => \N__34528\,
            in1 => \N__34609\,
            in2 => \N__32493\,
            in3 => \N__34491\,
            lcout => \c0.n24_adj_2340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1012_2_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32749\,
            in2 => \_gnd_net_\,
            in3 => \N__34799\,
            lcout => \c0.n2124\,
            ltout => \c0.n2124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_498_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__34160\,
            in1 => \N__35120\,
            in2 => \N__32478\,
            in3 => \N__37472\,
            lcout => \c0.n17_adj_2214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i44_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__32475\,
            in1 => \N__35277\,
            in2 => \N__32709\,
            in3 => \N__40425\,
            lcout => \c0.data_in_frame_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_654_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__32607\,
            in1 => \N__34833\,
            in2 => \N__32532\,
            in3 => \N__34944\,
            lcout => \c0.n26_adj_2368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_634_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32600\,
            in1 => \N__38885\,
            in2 => \_gnd_net_\,
            in3 => \N__34608\,
            lcout => \c0.n16474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_589_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__35325\,
            in1 => \N__33416\,
            in2 => \N__32589\,
            in3 => \N__32574\,
            lcout => \c0.n24_adj_2317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37690\,
            in1 => \N__40408\,
            in2 => \N__35292\,
            in3 => \N__34895\,
            lcout => \c0.data_in_frame_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__40406\,
            in1 => \N__37692\,
            in2 => \N__36688\,
            in3 => \N__34800\,
            lcout => \c0.data_in_frame_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__40578\,
            in1 => \N__45131\,
            in2 => \N__34614\,
            in3 => \N__40409\,
            lcout => \c0.data_in_frame_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_730_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__32892\,
            in1 => \N__32810\,
            in2 => \N__39219\,
            in3 => \N__33039\,
            lcout => \c0.n17076\,
            ltout => \c0.n17076_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__37691\,
            in1 => \N__45132\,
            in2 => \N__32568\,
            in3 => \N__32750\,
            lcout => \c0.data_in_frame_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45130\,
            in1 => \N__32531\,
            in2 => \_gnd_net_\,
            in3 => \N__32565\,
            lcout => data_in_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__40577\,
            in1 => \N__40407\,
            in2 => \N__39998\,
            in3 => \N__39477\,
            lcout => \c0.data_in_frame_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_539_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34854\,
            in2 => \_gnd_net_\,
            in3 => \N__36947\,
            lcout => \c0.n10215\,
            ltout => \c0.n10215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_526_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32745\,
            in1 => \N__34890\,
            in2 => \N__32724\,
            in3 => \N__34796\,
            lcout => \c0.n17206\,
            ltout => \c0.n17206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1026_2_lut_3_lut_4_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37376\,
            in1 => \N__41030\,
            in2 => \N__32721\,
            in3 => \N__34763\,
            lcout => \c0.n2138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__37730\,
            in1 => \N__34772\,
            in2 => \N__40433\,
            in3 => \N__39552\,
            lcout => \c0.data_in_frame_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_495_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111011111"
        )
    port map (
            in0 => \N__34980\,
            in1 => \N__32718\,
            in2 => \N__34522\,
            in3 => \N__40021\,
            lcout => \c0.n26_adj_2210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i41_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__40410\,
            in1 => \N__36802\,
            in2 => \N__32696\,
            in3 => \N__34959\,
            lcout => \c0.data_in_frame_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__36876\,
            in1 => \N__40411\,
            in2 => \N__34865\,
            in3 => \N__37729\,
            lcout => \c0.data_in_frame_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__40022\,
            in1 => \N__36803\,
            in2 => \N__40434\,
            in3 => \N__40618\,
            lcout => \c0.data_in_frame_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_491_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111001111101"
        )
    port map (
            in0 => \N__37443\,
            in1 => \N__34820\,
            in2 => \N__33417\,
            in3 => \N__32618\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_480_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__37396\,
            in1 => \N__39993\,
            in2 => \N__40989\,
            in3 => \N__37464\,
            lcout => OPEN,
            ltout => \c0.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__38892\,
            in1 => \N__34613\,
            in2 => \N__32967\,
            in3 => \N__34806\,
            lcout => OPEN,
            ltout => \c0.n30_adj_2213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_517_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32964\,
            in1 => \N__32958\,
            in2 => \N__32952\,
            in3 => \N__32949\,
            lcout => n31_adj_2415,
            ltout => \n31_adj_2415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_3_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__35743\,
            in1 => \_gnd_net_\,
            in2 => \N__32940\,
            in3 => \N__33437\,
            lcout => n1_adj_2486,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_651_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40988\,
            in1 => \N__32937\,
            in2 => \N__34869\,
            in3 => \N__36949\,
            lcout => \c0.n16352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_635_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__32916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35026\,
            lcout => \c0.n6_adj_2358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i27_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__40610\,
            in1 => \N__34364\,
            in2 => \N__36862\,
            in3 => \N__39359\,
            lcout => \c0.data_in_frame_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_726_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__32888\,
            in1 => \N__39200\,
            in2 => \N__32811\,
            in3 => \N__33013\,
            lcout => \c0.n17072\,
            ltout => \c0.n17072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__37733\,
            in1 => \N__45135\,
            in2 => \N__32769\,
            in3 => \N__33412\,
            lcout => \c0.data_in_frame_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_620_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__36072\,
            in1 => \N__40197\,
            in2 => \N__35745\,
            in3 => \N__35532\,
            lcout => \FRAME_MATCHER_i_31__N_1273\,
            ltout => \FRAME_MATCHER_i_31__N_1273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_630_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35723\,
            in2 => \N__33390\,
            in3 => \N__35817\,
            lcout => n17086,
            ltout => \n17086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_626_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__35818\,
            in1 => \_gnd_net_\,
            in2 => \N__33387\,
            in3 => \N__35725\,
            lcout => \c0.n1034\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_641_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35724\,
            in2 => \_gnd_net_\,
            in3 => \N__35819\,
            lcout => \FRAME_MATCHER_i_31__N_1275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4980_2_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33382\,
            in2 => \_gnd_net_\,
            in3 => \N__33360\,
            lcout => n10088,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_707_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33336\,
            in2 => \_gnd_net_\,
            in3 => \N__40702\,
            lcout => \c0.n16666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_708_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40711\,
            in3 => \N__33291\,
            lcout => \c0.n16674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_644_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33553\,
            in2 => \_gnd_net_\,
            in3 => \N__33011\,
            lcout => n10140,
            ltout => \n10140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41592\,
            in2 => \N__32970\,
            in3 => \N__44414\,
            lcout => n17089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_629_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35820\,
            lcout => n44,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_753_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__35821\,
            in1 => \N__41445\,
            in2 => \N__35746\,
            in3 => \N__41296\,
            lcout => \c0.n8_adj_2385\,
            ltout => \c0.n8_adj_2385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_716_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33585\,
            in3 => \N__37809\,
            lcout => \c0.n16670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14591_2_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40198\,
            in2 => \_gnd_net_\,
            in3 => \N__35534\,
            lcout => OPEN,
            ltout => \c0.n17367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_418_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__42014\,
            in1 => \N__35702\,
            in2 => \N__33561\,
            in3 => \N__36061\,
            lcout => \c0.n10139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_751_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__36062\,
            in1 => \N__40199\,
            in2 => \_gnd_net_\,
            in3 => \N__35535\,
            lcout => n9,
            ltout => \n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_698_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__39753\,
            in1 => \N__35703\,
            in2 => \N__33558\,
            in3 => \N__33555\,
            lcout => \c0.n11833\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33489\,
            in1 => \N__33793\,
            in2 => \N__40761\,
            in3 => \N__33470\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_797_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__39754\,
            in1 => \N__33436\,
            in2 => \N__35744\,
            in3 => \N__35463\,
            lcout => OPEN,
            ltout => \n21_adj_2487_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i1_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__41389\,
            in1 => \N__33702\,
            in2 => \N__33747\,
            in3 => \N__33708\,
            lcout => \FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_798_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__35904\,
            in1 => \N__35462\,
            in2 => \N__35958\,
            in3 => \N__33744\,
            lcout => n6_adj_2410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i7_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44945\,
            in1 => \N__44772\,
            in2 => \N__33798\,
            in3 => \N__44564\,
            lcout => \c0.FRAME_MATCHER_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49770\,
            ce => 'H',
            sr => \N__33777\
        );

    \i14574_2_lut_3_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__35712\,
            in1 => \N__33698\,
            in2 => \_gnd_net_\,
            in3 => \N__35828\,
            lcout => n17349,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_428_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35711\,
            in2 => \_gnd_net_\,
            in3 => \N__35551\,
            lcout => \c0.n51_adj_2173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_420_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__35552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40239\,
            lcout => \c0.n10166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10658_2_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33656\,
            in2 => \_gnd_net_\,
            in3 => \N__41741\,
            lcout => \c0.FRAME_MATCHER_i_31_N_1310_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_765_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__35210\,
            in1 => \N__41472\,
            in2 => \N__41423\,
            in3 => \N__41333\,
            lcout => \c0.n16696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__47438\,
            in1 => \N__42912\,
            in2 => \N__42446\,
            in3 => \N__42367\,
            lcout => byte_transmit_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_745_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49170\,
            in1 => \N__47120\,
            in2 => \_gnd_net_\,
            in3 => \N__49099\,
            lcout => \c0.n17270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__42716\,
            in1 => \N__42945\,
            in2 => \N__42448\,
            in3 => \N__42369\,
            lcout => byte_transmit_counter_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__2__2190_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33830\,
            in1 => \_gnd_net_\,
            in2 => \N__49962\,
            in3 => \N__48718\,
            lcout => data_out_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__43050\,
            in1 => \N__46379\,
            in2 => \N__42447\,
            in3 => \N__42368\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__3__2189_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49930\,
            in1 => \N__33816\,
            in2 => \_gnd_net_\,
            in3 => \N__48825\,
            lcout => data_out_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13368_2_lut_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33794\,
            in2 => \_gnd_net_\,
            in3 => \N__40807\,
            lcout => \c0.n16141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__7__2201_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50150\,
            in1 => \N__33765\,
            in2 => \N__48157\,
            in3 => \N__42474\,
            lcout => \c0.data_out_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => \N__50588\,
            sr => \_gnd_net_\
        );

    \c0.data_out_1__1__2247_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__48381\,
            in1 => \N__48121\,
            in2 => \_gnd_net_\,
            in3 => \N__50151\,
            lcout => \c0.data_out_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => \N__50588\,
            sr => \_gnd_net_\
        );

    \c0.i15145_3_lut_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__45733\,
            in1 => \N__48380\,
            in2 => \_gnd_net_\,
            in3 => \N__47119\,
            lcout => OPEN,
            ltout => \c0.n17639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4__2204_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__48123\,
            in1 => \N__50153\,
            in2 => \N__33948\,
            in3 => \N__33944\,
            lcout => \c0.data_out_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => \N__50588\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__6__2202_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33929\,
            in1 => \N__48122\,
            in2 => \N__33915\,
            in3 => \N__50152\,
            lcout => \c0.data_out_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49792\,
            ce => \N__50588\,
            sr => \_gnd_net_\
        );

    \c0.i15088_2_lut_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45732\,
            in2 => \_gnd_net_\,
            in3 => \N__47700\,
            lcout => \c0.n17671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14999_3_lut_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__45728\,
            in1 => \_gnd_net_\,
            in2 => \N__48418\,
            in3 => \N__47877\,
            lcout => OPEN,
            ltout => \c0.n17631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__3__2205_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33899\,
            in1 => \N__48128\,
            in2 => \N__33885\,
            in3 => \N__50157\,
            lcout => \c0.data_out_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49802\,
            ce => \N__50566\,
            sr => \_gnd_net_\
        );

    \c0.i15033_3_lut_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__48392\,
            in1 => \N__43362\,
            in2 => \_gnd_net_\,
            in3 => \N__47876\,
            lcout => OPEN,
            ltout => \c0.n17627_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__2__2206_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33881\,
            in1 => \N__48127\,
            in2 => \N__33867\,
            in3 => \N__50156\,
            lcout => \c0.data_out_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49802\,
            ce => \N__50566\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__5__2203_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33863\,
            in1 => \N__48129\,
            in2 => \N__33849\,
            in3 => \N__50158\,
            lcout => \c0.data_out_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49802\,
            ce => \N__50566\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_720_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45727\,
            in1 => \N__43361\,
            in2 => \_gnd_net_\,
            in3 => \N__47875\,
            lcout => \c0.n10326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__33954\,
            in1 => \N__46252\,
            in2 => \N__33993\,
            in3 => \N__47482\,
            lcout => OPEN,
            ltout => \c0.n18268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18268_bdd_4_lut_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__46253\,
            in1 => \N__34035\,
            in2 => \N__33999\,
            in3 => \N__34080\,
            lcout => n18271,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_3_lut_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__42640\,
            in1 => \N__42583\,
            in2 => \_gnd_net_\,
            in3 => \N__36370\,
            lcout => OPEN,
            ltout => \c0.tx.n55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110111000000"
        )
    port map (
            in0 => \N__36371\,
            in1 => \N__44214\,
            in2 => \N__33996\,
            in3 => \N__42550\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48963\,
            in1 => \N__45646\,
            in2 => \_gnd_net_\,
            in3 => \N__47670\,
            lcout => \c0.n5_adj_2136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47669\,
            in1 => \N__48573\,
            in2 => \_gnd_net_\,
            in3 => \N__42129\,
            lcout => n8_adj_2447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__4__2196_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__48964\,
            in1 => \N__33984\,
            in2 => \N__43718\,
            in3 => \N__46905\,
            lcout => \c0.data_out_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15376_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__34050\,
            in1 => \N__46250\,
            in2 => \N__33966\,
            in3 => \N__47481\,
            lcout => OPEN,
            ltout => \c0.n18172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18172_bdd_4_lut_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__46251\,
            in1 => \N__36444\,
            in2 => \N__33957\,
            in3 => \N__34029\,
            lcout => n18175,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15173_2_lut_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49065\,
            lcout => \c0.n17764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15100_2_lut_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47675\,
            in2 => \_gnd_net_\,
            in3 => \N__34200\,
            lcout => \c0.n17676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__6__2194_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__47230\,
            in1 => \N__43693\,
            in2 => \N__34074\,
            in3 => \N__46918\,
            lcout => \c0.data_out_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15108_2_lut_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47672\,
            in2 => \_gnd_net_\,
            in3 => \N__47085\,
            lcout => \c0.n17703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__4__2244_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__34044\,
            in1 => \N__48388\,
            in2 => \N__50576\,
            in3 => \N__50266\,
            lcout => \c0.data_out_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15103_2_lut_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47674\,
            in2 => \_gnd_net_\,
            in3 => \N__34043\,
            lcout => \c0.n17675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15101_2_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34007\,
            lcout => \c0.n17697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_784_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__34020\,
            in1 => \N__46400\,
            in2 => \N__47352\,
            in3 => \N__46288\,
            lcout => OPEN,
            ltout => \n10_adj_2408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__44104\,
            in1 => \N__38249\,
            in2 => \N__34011\,
            in3 => \N__43841\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__3__2237_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__34008\,
            in1 => \N__50505\,
            in2 => \N__48417\,
            in3 => \N__50320\,
            lcout => \c0.data_out_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__0__2232_LC_11_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35858\,
            in1 => \N__50555\,
            in2 => \_gnd_net_\,
            in3 => \N__34184\,
            lcout => data_out_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__5__2251_LC_11_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34183\,
            in1 => \N__50552\,
            in2 => \_gnd_net_\,
            in3 => \N__34227\,
            lcout => data_out_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__2__2238_LC_11_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__50329\,
            in1 => \N__50554\,
            in2 => \_gnd_net_\,
            in3 => \N__34215\,
            lcout => data_out_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_1195_i1_3_lut_LC_11_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48384\,
            in1 => \N__48133\,
            in2 => \_gnd_net_\,
            in3 => \N__50328\,
            lcout => n2699,
            ltout => \n2699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__4__2228_LC_11_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50556\,
            in2 => \N__34203\,
            in3 => \N__34199\,
            lcout => data_out_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__2__2230_LC_11_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34185\,
            in1 => \N__50553\,
            in2 => \_gnd_net_\,
            in3 => \N__34173\,
            lcout => data_out_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__37745\,
            in1 => \N__34153\,
            in2 => \N__39555\,
            in3 => \N__39390\,
            lcout => \c0.data_in_frame_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i6_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__34131\,
            in1 => \N__34442\,
            in2 => \N__39701\,
            in3 => \N__42053\,
            lcout => \c0.byte_transmit_counter2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49701\,
            ce => 'H',
            sr => \N__34119\
        );

    \c0.i10953_1_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34409\,
            lcout => \c0.tx2_transmit_N_1996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_756_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__34410\,
            in1 => \N__34397\,
            in2 => \N__35765\,
            in3 => \N__35583\,
            lcout => \c0.n16261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_537_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34484\,
            in1 => \N__34437\,
            in2 => \N__39622\,
            in3 => \N__34416\,
            lcout => \c0.n13628\,
            ltout => \c0.n13628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_687_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35582\,
            in2 => \N__34401\,
            in3 => \N__34396\,
            lcout => n488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_601_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__34368\,
            in1 => \N__34238\,
            in2 => \N__35346\,
            in3 => \N__36921\,
            lcout => \c0.n21_adj_2323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_624_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41033\,
            in1 => \N__37045\,
            in2 => \N__34350\,
            in3 => \N__36954\,
            lcout => \c0.n16353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14698_4_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__40316\,
            in1 => \N__39825\,
            in2 => \N__34314\,
            in3 => \N__40144\,
            lcout => OPEN,
            ltout => \c0.n17475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i6_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__39826\,
            in1 => \N__39934\,
            in2 => \N__34329\,
            in3 => \N__39877\,
            lcout => \c0.data_out_frame2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_662_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111101"
        )
    port map (
            in0 => \N__34281\,
            in1 => \N__34269\,
            in2 => \N__34263\,
            in3 => \N__34239\,
            lcout => \c0.n28_adj_2374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14692_4_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__40315\,
            in1 => \N__39824\,
            in2 => \N__34714\,
            in3 => \N__40143\,
            lcout => OPEN,
            ltout => \c0.n17469_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i8_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__39827\,
            in1 => \N__39935\,
            in2 => \N__34728\,
            in3 => \N__39878\,
            lcout => \c0.data_out_frame2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_563_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37043\,
            in1 => \N__34529\,
            in2 => \N__34680\,
            in3 => \N__34562\,
            lcout => OPEN,
            ltout => \c0.n17114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_643_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__37378\,
            in1 => \N__34659\,
            in2 => \N__34641\,
            in3 => \N__40020\,
            lcout => \c0.n18_adj_2360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_623_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37044\,
            in1 => \N__40953\,
            in2 => \N__34638\,
            in3 => \N__34563\,
            lcout => \c0.n17214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_546_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40019\,
            in2 => \_gnd_net_\,
            in3 => \N__39983\,
            lcout => OPEN,
            ltout => \c0.n17101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_547_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34607\,
            in1 => \N__34771\,
            in2 => \N__34581\,
            in3 => \N__37377\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_554_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38828\,
            in1 => \N__38900\,
            in2 => \N__34578\,
            in3 => \N__34575\,
            lcout => \c0.n10407\,
            ltout => \c0.n10407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_604_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34554\,
            in1 => \N__40952\,
            in2 => \N__34533\,
            in3 => \N__34530\,
            lcout => \c0.n17215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__37379\,
            in1 => \N__37728\,
            in2 => \N__40502\,
            in3 => \N__40426\,
            lcout => \c0.data_in_frame_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1016_2_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34764\,
            in2 => \_gnd_net_\,
            in3 => \N__37380\,
            lcout => \c0.n2128\,
            ltout => \c0.n2128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_602_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__34973\,
            in1 => \N__34958\,
            in2 => \N__34947\,
            in3 => \N__37502\,
            lcout => \c0.n19_adj_2324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__0__2269_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36804\,
            in1 => \N__39194\,
            in2 => \_gnd_net_\,
            in3 => \N__34923\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1008_2_lut_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34894\,
            in2 => \_gnd_net_\,
            in3 => \N__34855\,
            lcout => \c0.n2120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_4_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111101101111"
        )
    port map (
            in0 => \N__34797\,
            in1 => \N__36898\,
            in2 => \N__37047\,
            in3 => \N__34765\,
            lcout => OPEN,
            ltout => \c0.n22_adj_2201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_482_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111011"
        )
    port map (
            in0 => \N__37417\,
            in1 => \N__38827\,
            in2 => \N__34809\,
            in3 => \N__36917\,
            lcout => \c0.n27_adj_2202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1014_2_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34766\,
            lcout => \c0.n2126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__37731\,
            in1 => \N__40423\,
            in2 => \N__39469\,
            in3 => \N__36953\,
            lcout => \c0.data_in_frame_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__37732\,
            in1 => \N__36798\,
            in2 => \N__35119\,
            in3 => \N__39360\,
            lcout => \c0.data_in_frame_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__37973\,
            in1 => \N__45258\,
            in2 => \N__36861\,
            in3 => \N__45156\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_677_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__35550\,
            in1 => \N__35750\,
            in2 => \N__36093\,
            in3 => \N__40235\,
            lcout => \c0.n5817\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__6__2263_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39541\,
            in1 => \N__39094\,
            in2 => \_gnd_net_\,
            in3 => \N__35074\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_691_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__40234\,
            in1 => \N__36086\,
            in2 => \N__35758\,
            in3 => \N__35549\,
            lcout => \c0.n5815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10706_2_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37327\,
            in2 => \_gnd_net_\,
            in3 => \N__40814\,
            lcout => \c0.n13381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__0__2293_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39093\,
            in1 => \N__35030\,
            in2 => \_gnd_net_\,
            in3 => \N__35055\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_794_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__35786\,
            in1 => \N__44424\,
            in2 => \N__41613\,
            in3 => \N__36109\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__1__2268_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39205\,
            in1 => \_gnd_net_\,
            in2 => \N__39478\,
            in3 => \N__34999\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__37734\,
            in1 => \N__36799\,
            in2 => \N__41034\,
            in3 => \N__40432\,
            lcout => \c0.data_in_frame_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__1__2284_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39204\,
            in1 => \N__35370\,
            in2 => \_gnd_net_\,
            in3 => \N__35409\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i25_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__37487\,
            in1 => \N__36800\,
            in2 => \N__40624\,
            in3 => \N__39372\,
            lcout => \c0.data_in_frame_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i30_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__39370\,
            in1 => \N__40614\,
            in2 => \N__35345\,
            in3 => \N__36679\,
            lcout => \c0.data_in_frame_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__37735\,
            in1 => \N__35317\,
            in2 => \N__35298\,
            in3 => \N__39371\,
            lcout => \c0.data_in_frame_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__3__2266_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35293\,
            in1 => \N__39142\,
            in2 => \_gnd_net_\,
            in3 => \N__35233\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43191\,
            in1 => \N__37285\,
            in2 => \N__43119\,
            in3 => \N__35214\,
            lcout => OPEN,
            ltout => \c0.n47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i27_4_lut_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35178\,
            in1 => \N__37773\,
            in2 => \N__35166\,
            in3 => \N__35163\,
            lcout => OPEN,
            ltout => \c0.n56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35157\,
            in1 => \N__40689\,
            in2 => \N__35145\,
            in3 => \N__35142\,
            lcout => \c0.n10018\,
            ltout => \c0.n10018_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__36071\,
            in1 => \N__35682\,
            in2 => \N__35130\,
            in3 => \N__40193\,
            lcout => \FRAME_MATCHER_i_31__N_1272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_636_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__40192\,
            in1 => \N__36070\,
            in2 => \_gnd_net_\,
            in3 => \N__35533\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i0_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101110101010"
        )
    port map (
            in0 => \N__35790\,
            in1 => \N__35775\,
            in2 => \N__40220\,
            in3 => \N__35445\,
            lcout => \FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_2261_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100100010"
        )
    port map (
            in0 => \N__35719\,
            in1 => \N__40219\,
            in2 => \N__35622\,
            in3 => \N__36069\,
            lcout => \c0.r_SM_Main_2_N_2034_0_adj_2167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49771\,
            ce => 'H',
            sr => \N__35553\
        );

    \i1_4_lut_adj_796_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__35438\,
            in1 => \N__35499\,
            in2 => \N__35493\,
            in3 => \N__35453\,
            lcout => n17063,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__35454\,
            in1 => \N__35439\,
            in2 => \N__35871\,
            in3 => \N__35421\,
            lcout => n17090,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41967\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42015\,
            lcout => n3_adj_2485,
            ltout => \n3_adj_2485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_795_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110101010"
        )
    port map (
            in0 => \N__35430\,
            in1 => \N__35420\,
            in2 => \N__35412\,
            in3 => \N__36120\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_689_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48713\,
            in1 => \N__42143\,
            in2 => \_gnd_net_\,
            in3 => \N__48815\,
            lcout => \c0.n10188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14651_4_lut_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010001100"
        )
    port map (
            in0 => \N__36279\,
            in1 => \N__36246\,
            in2 => \N__36210\,
            in3 => \N__36170\,
            lcout => n17428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_217_Select_2_i4_3_lut_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__36118\,
            in1 => \_gnd_net_\,
            in2 => \N__35957\,
            in3 => \N__35903\,
            lcout => OPEN,
            ltout => \n4_adj_2417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__36138\,
            in1 => \N__36129\,
            in2 => \N__36123\,
            in3 => \N__36119\,
            lcout => \FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14652_3_lut_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__36015\,
            in1 => \N__35994\,
            in2 => \_gnd_net_\,
            in3 => \N__35988\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_792_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35950\,
            in2 => \_gnd_net_\,
            in3 => \N__35902\,
            lcout => n6_adj_2488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37994\,
            in1 => \N__35862\,
            in2 => \_gnd_net_\,
            in3 => \N__47787\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_460_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43469\,
            in2 => \_gnd_net_\,
            in3 => \N__44285\,
            lcout => \c0.n17264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_782_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__35844\,
            in1 => \N__46375\,
            in2 => \N__42207\,
            in3 => \N__46290\,
            lcout => OPEN,
            ltout => \n10_adj_2409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43814\,
            in1 => \N__44105\,
            in2 => \N__36357\,
            in3 => \N__36392\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49169\,
            in1 => \N__48717\,
            in2 => \_gnd_net_\,
            in3 => \N__47794\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__47795\,
            in1 => \N__45465\,
            in2 => \N__36354\,
            in3 => \N__47458\,
            lcout => n10_adj_2450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__43813\,
            in1 => \N__42993\,
            in2 => \N__42452\,
            in3 => \N__42366\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15366_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__36351\,
            in1 => \N__46289\,
            in2 => \N__38274\,
            in3 => \N__47431\,
            lcout => \c0.n18166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15212_2_lut_3_lut_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__48276\,
            in1 => \N__48114\,
            in2 => \_gnd_net_\,
            in3 => \N__50135\,
            lcout => \data_out_10__7__N_110\,
            ltout => \data_out_10__7__N_110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__4__2188_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36345\,
            in1 => \_gnd_net_\,
            in2 => \N__36321\,
            in3 => \N__48472\,
            lcout => data_out_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i2_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101011010010"
        )
    port map (
            in0 => \N__50136\,
            in1 => \N__48278\,
            in2 => \N__48155\,
            in3 => \N__38343\,
            lcout => \UART_TRANSMITTER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__6__2186_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49929\,
            in1 => \N__36318\,
            in2 => \_gnd_net_\,
            in3 => \N__43386\,
            lcout => data_out_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__2__2246_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__50137\,
            in1 => \N__48277\,
            in2 => \N__50587\,
            in3 => \N__36293\,
            lcout => \c0.data_out_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15075_2_lut_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__47802\,
            in1 => \N__42768\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n17696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n18070_bdd_4_lut_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__42626\,
            in1 => \N__38694\,
            in2 => \N__36426\,
            in3 => \N__36378\,
            lcout => OPEN,
            ltout => \n18073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i33_3_lut_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42578\,
            in2 => \N__36432\,
            in3 => \N__38232\,
            lcout => \c0.tx.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__45927\,
            in1 => \N__44014\,
            in2 => \N__44212\,
            in3 => \N__43950\,
            lcout => \c0.tx.n10688\,
            ltout => \c0.tx.n10688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44203\,
            in2 => \N__36429\,
            in3 => \N__42579\,
            lcout => \c0.tx.r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__36425\,
            in1 => \N__42231\,
            in2 => \N__43842\,
            in3 => \N__44099\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__1__2191_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36414\,
            in1 => \_gnd_net_\,
            in2 => \N__49963\,
            in3 => \N__42136\,
            lcout => data_out_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_15385_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__42625\,
            in1 => \N__36393\,
            in2 => \N__43608\,
            in3 => \N__42546\,
            lcout => n18070,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011110000"
        )
    port map (
            in0 => \N__42584\,
            in1 => \N__44204\,
            in2 => \N__42641\,
            in3 => \N__36372\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__47677\,
            in1 => \N__42894\,
            in2 => \N__42461\,
            in3 => \N__42350\,
            lcout => byte_transmit_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_607_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__50719\,
            in1 => \N__38664\,
            in2 => \N__48099\,
            in3 => \N__38558\,
            lcout => n4_adj_2419,
            ltout => \n4_adj_2419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__50205\,
            in1 => \_gnd_net_\,
            in2 => \N__36465\,
            in3 => \_gnd_net_\,
            lcout => n5_adj_2407,
            ltout => \n5_adj_2407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_788_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48020\,
            in1 => \N__48298\,
            in2 => \N__36462\,
            in3 => \N__38214\,
            lcout => n10_adj_2444,
            ltout => \n10_adj_2444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__42456\,
            in1 => \N__42852\,
            in2 => \N__36459\,
            in3 => \N__46255\,
            lcout => byte_transmit_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i52_4_lut_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__36456\,
            in1 => \N__47497\,
            in2 => \N__48759\,
            in3 => \N__47676\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15147_4_lut_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010101000"
        )
    port map (
            in0 => \N__50206\,
            in1 => \N__36450\,
            in2 => \N__48371\,
            in3 => \N__38340\,
            lcout => n17765,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__44016\,
            in1 => \N__45894\,
            in2 => \N__44213\,
            in3 => \N__43956\,
            lcout => \c0.tx.r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10536_2_lut_3_lut_4_lut_LC_12_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__38564\,
            in1 => \N__38745\,
            in2 => \N__50742\,
            in3 => \N__38647\,
            lcout => \c0.n22_adj_2313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10543_2_lut_3_lut_4_lut_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__50718\,
            in1 => \N__38638\,
            in2 => \N__38415\,
            in3 => \N__38562\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10539_2_lut_3_lut_4_lut_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__38563\,
            in1 => \N__38493\,
            in2 => \N__50741\,
            in3 => \N__38646\,
            lcout => \c0.n25_adj_2386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_12_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43629\,
            in1 => \N__47653\,
            in2 => \_gnd_net_\,
            in3 => \N__48864\,
            lcout => \c0.n5_adj_2163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10535_2_lut_3_lut_4_lut_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__38565\,
            in1 => \N__38454\,
            in2 => \N__50743\,
            in3 => \N__38648\,
            lcout => \c0.n21_adj_2262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i0_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38304\,
            in2 => \N__38289\,
            in3 => \_gnd_net_\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_12_31_0_\,
            carryout => \c0.n16066\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i1_LC_12_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36495\,
            in2 => \_gnd_net_\,
            in3 => \N__36489\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \c0.n16066\,
            carryout => \c0.n16067\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i2_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38763\,
            in2 => \_gnd_net_\,
            in3 => \N__36486\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \c0.n16067\,
            carryout => \c0.n16068\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i3_LC_12_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36483\,
            in3 => \N__36474\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \c0.n16068\,
            carryout => \c0.n16069\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i4_LC_12_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38355\,
            in2 => \_gnd_net_\,
            in3 => \N__36471\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \c0.n16069\,
            carryout => \c0.n16070\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i5_LC_12_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38298\,
            in3 => \N__36468\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \c0.n16070\,
            carryout => \c0.n16071\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i6_LC_12_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36591\,
            in3 => \N__36582\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \c0.n16071\,
            carryout => \c0.n16072\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i7_LC_12_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36579\,
            in2 => \_gnd_net_\,
            in3 => \N__36573\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \c0.n16072\,
            carryout => \c0.n16073\,
            clk => \N__49831\,
            ce => \N__36551\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i8_LC_12_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38460\,
            in2 => \_gnd_net_\,
            in3 => \N__36570\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_12_32_0_\,
            carryout => \c0.n16074\,
            clk => \N__49836\,
            ce => \N__36552\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i9_LC_12_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38322\,
            in3 => \N__36567\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \c0.n16074\,
            carryout => \c0.n16075\,
            clk => \N__49836\,
            ce => \N__36552\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i10_LC_12_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38718\,
            in2 => \_gnd_net_\,
            in3 => \N__36564\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \c0.n16075\,
            carryout => \c0.n16076\,
            clk => \N__49836\,
            ce => \N__36552\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i11_LC_12_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38511\,
            in2 => \_gnd_net_\,
            in3 => \N__36561\,
            lcout => \c0.delay_counter_11\,
            ltout => OPEN,
            carryin => \c0.n16076\,
            carryout => \c0.n16077\,
            clk => \N__49836\,
            ce => \N__36552\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i12_LC_12_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38778\,
            in2 => \_gnd_net_\,
            in3 => \N__36558\,
            lcout => \c0.delay_counter_12\,
            ltout => OPEN,
            carryin => \c0.n16077\,
            carryout => \c0.n16078\,
            clk => \N__49836\,
            ce => \N__36552\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_2361__i13_LC_12_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38700\,
            in2 => \_gnd_net_\,
            in3 => \N__36555\,
            lcout => \c0.delay_counter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49836\,
            ce => \N__36552\,
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_678_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__36528\,
            in1 => \N__36522\,
            in2 => \N__36513\,
            in3 => \N__36501\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__37961\,
            in1 => \N__45216\,
            in2 => \N__36778\,
            in3 => \N__45175\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__39936\,
            in1 => \N__39875\,
            in2 => \N__39846\,
            in3 => \N__40632\,
            lcout => \c0.data_out_frame2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36738\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_561_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40243\,
            lcout => \c0.n26_adj_2174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__36720\,
            in1 => \N__39572\,
            in2 => \N__40501\,
            in3 => \N__45219\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__45217\,
            in1 => \N__37962\,
            in2 => \N__39446\,
            in3 => \N__36718\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__36719\,
            in1 => \N__36655\,
            in2 => \N__45294\,
            in3 => \N__45218\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_603_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36618\,
            in1 => \N__37341\,
            in2 => \N__36609\,
            in3 => \N__36597\,
            lcout => \c0.n4494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15063_3_lut_4_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__37568\,
            in1 => \N__41957\,
            in2 => \N__40146\,
            in3 => \N__40246\,
            lcout => \c0.n17688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_413_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37191\,
            in2 => \_gnd_net_\,
            in3 => \N__37112\,
            lcout => \c0.n15171\,
            ltout => \c0.n15171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__37046\,
            in1 => \N__39519\,
            in2 => \N__37050\,
            in3 => \N__40430\,
            lcout => \c0.data_in_frame_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_676_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111011111111"
        )
    port map (
            in0 => \N__38796\,
            in1 => \N__37017\,
            in2 => \N__36999\,
            in3 => \N__36978\,
            lcout => OPEN,
            ltout => \c0.n27_adj_2381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_702_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__40244\,
            in1 => \N__36972\,
            in2 => \N__36966\,
            in3 => \N__36963\,
            lcout => \c0.n12491\,
            ltout => \c0.n12491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15059_3_lut_4_lut_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__37622\,
            in1 => \N__41956\,
            in2 => \N__36957\,
            in3 => \N__40245\,
            lcout => \c0.n17686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_458_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41031\,
            in2 => \_gnd_net_\,
            in3 => \N__36948\,
            lcout => \c0.n10259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__37439\,
            in1 => \N__37740\,
            in2 => \N__39480\,
            in3 => \N__39388\,
            lcout => \c0.data_in_frame_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__39387\,
            in1 => \N__40500\,
            in2 => \N__37746\,
            in3 => \N__36902\,
            lcout => \c0.data_in_frame_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__36840\,
            in1 => \N__37741\,
            in2 => \N__37422\,
            in3 => \N__39389\,
            lcout => \c0.data_in_frame_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i5_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__37644\,
            in1 => \N__37623\,
            in2 => \N__39729\,
            in3 => \N__39946\,
            lcout => \c0.data_out_frame2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i4_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__39945\,
            in1 => \N__39725\,
            in2 => \N__37583\,
            in3 => \N__37593\,
            lcout => \c0.data_out_frame2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_587_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__37524\,
            in1 => \N__37503\,
            in2 => \N__37491\,
            in3 => \N__37473\,
            lcout => OPEN,
            ltout => \c0.n18_adj_2316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_600_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111011"
        )
    port map (
            in0 => \N__37438\,
            in1 => \N__37418\,
            in2 => \N__37401\,
            in3 => \N__37389\,
            lcout => \c0.n23_adj_2322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i23_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44982\,
            in1 => \N__44714\,
            in2 => \N__37334\,
            in3 => \N__44566\,
            lcout => \c0.FRAME_MATCHER_state_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49747\,
            ce => 'H',
            sr => \N__37308\
        );

    \c0.FRAME_MATCHER_state_i11_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44915\,
            in1 => \N__44676\,
            in2 => \N__37295\,
            in3 => \N__44512\,
            lcout => \c0.FRAME_MATCHER_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49759\,
            ce => 'H',
            sr => \N__37269\
        );

    \c0.i1_2_lut_adj_754_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41227\,
            in2 => \_gnd_net_\,
            in3 => \N__40718\,
            lcout => \c0.n16658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37253\,
            in2 => \_gnd_net_\,
            in3 => \N__39263\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_52_i4_2_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__37917\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37947\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_55_i4_2_lut_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__37948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37918\,
            lcout => n4_adj_2427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_56_i4_2_lut_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__37919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37949\,
            lcout => n4_adj_2416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i10445_2_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37950\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37920\,
            lcout => n13116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_397_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__37875\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37836\,
            lcout => n9999,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43158\,
            in1 => \N__37808\,
            in2 => \N__41192\,
            in3 => \N__37765\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i30_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37767\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41545\,
            lcout => \c0.FRAME_MATCHER_state_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49772\,
            ce => 'H',
            sr => \N__37755\
        );

    \c0.i1_2_lut_4_lut_adj_767_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__41322\,
            in1 => \N__41400\,
            in2 => \N__41492\,
            in3 => \N__37766\,
            lcout => \c0.n16698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_737_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__41188\,
            in1 => \N__41473\,
            in2 => \N__41417\,
            in3 => \N__41318\,
            lcout => \c0.n16710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_746_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__41263\,
            in1 => \N__41474\,
            in2 => \N__41418\,
            in3 => \N__41319\,
            lcout => \c0.n16704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_759_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__41320\,
            in1 => \N__41396\,
            in2 => \N__41491\,
            in3 => \N__43118\,
            lcout => \c0.n16688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_764_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__38069\,
            in1 => \N__41478\,
            in2 => \N__41419\,
            in3 => \N__41321\,
            lcout => \c0.n16718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i18_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44977\,
            in1 => \N__44677\,
            in2 => \N__40760\,
            in3 => \N__44599\,
            lcout => \c0.FRAME_MATCHER_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49784\,
            ce => 'H',
            sr => \N__40731\
        );

    \c0.FRAME_MATCHER_state_i27_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__44718\,
            in1 => \N__44565\,
            in2 => \N__45017\,
            in3 => \N__38065\,
            lcout => \c0.FRAME_MATCHER_state_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49794\,
            ce => 'H',
            sr => \N__38043\
        );

    \c0.data_out_8__0__2192_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38031\,
            in1 => \N__45406\,
            in2 => \_gnd_net_\,
            in3 => \N__49935\,
            lcout => \c0.data_out_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i53_4_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__47792\,
            in1 => \N__38001\,
            in2 => \N__38136\,
            in3 => \N__47454\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49006\,
            in1 => \N__48827\,
            in2 => \_gnd_net_\,
            in3 => \N__47793\,
            lcout => \c0.n3_adj_2193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__0__2240_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__50541\,
            in1 => \N__50154\,
            in2 => \_gnd_net_\,
            in3 => \N__37995\,
            lcout => data_out_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__7__2185_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__38157\,
            in1 => \_gnd_net_\,
            in2 => \N__45837\,
            in3 => \N__49934\,
            lcout => data_out_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__0__2256_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__38135\,
            in1 => \N__48150\,
            in2 => \N__50574\,
            in3 => \N__50155\,
            lcout => data_out_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__0__2208_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__38124\,
            in1 => \N__50542\,
            in2 => \N__43719\,
            in3 => \N__46817\,
            lcout => \c0.data_out_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_473_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45405\,
            in1 => \N__46507\,
            in2 => \N__45513\,
            in3 => \N__46759\,
            lcout => \c0.n17147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47796\,
            in1 => \N__43308\,
            in2 => \_gnd_net_\,
            in3 => \N__48925\,
            lcout => \c0.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__7__2193_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__43309\,
            in1 => \N__38103\,
            in2 => \N__43716\,
            in3 => \N__46922\,
            lcout => \c0.data_out_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_780_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__38166\,
            in1 => \N__46413\,
            in2 => \N__38082\,
            in3 => \N__46298\,
            lcout => OPEN,
            ltout => \n10_adj_2411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__44103\,
            in1 => \N__38265\,
            in2 => \N__38073\,
            in3 => \N__43815\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15044_4_lut_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__46784\,
            in1 => \N__42518\,
            in2 => \N__48404\,
            in3 => \N__44288\,
            lcout => \c0.n17653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_449_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42323\,
            in2 => \_gnd_net_\,
            in3 => \N__48465\,
            lcout => \c0.n10392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_697_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__50204\,
            in1 => \N__38349\,
            in2 => \N__48144\,
            in3 => \N__42655\,
            lcout => n4_adj_2414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i3_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110010"
        )
    port map (
            in0 => \N__48302\,
            in1 => \N__38220\,
            in2 => \N__43715\,
            in3 => \N__38280\,
            lcout => \UART_TRANSMITTER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43465\,
            in1 => \N__46997\,
            in2 => \_gnd_net_\,
            in3 => \N__47671\,
            lcout => \c0.n5_adj_2141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__43758\,
            in1 => \N__38264\,
            in2 => \N__42636\,
            in3 => \N__42555\,
            lcout => OPEN,
            ltout => \n18196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n18196_bdd_4_lut_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__43515\,
            in1 => \N__38253\,
            in2 => \N__38235\,
            in3 => \N__42624\,
            lcout => n18199,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i26_3_lut_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__44208\,
            in1 => \N__44015\,
            in2 => \_gnd_net_\,
            in3 => \N__38226\,
            lcout => \c0.tx.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15178_4_lut_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__50270\,
            in1 => \N__38341\,
            in2 => \N__48100\,
            in3 => \N__42656\,
            lcout => n17759,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15020_4_lut_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110011"
        )
    port map (
            in0 => \N__38424\,
            in1 => \N__42671\,
            in2 => \N__50721\,
            in3 => \N__43040\,
            lcout => n17664,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18166_bdd_4_lut_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__38205\,
            in1 => \N__38196\,
            in2 => \N__38184\,
            in3 => \N__46254\,
            lcout => n18169,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i149_3_lut_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__50688\,
            in1 => \N__42670\,
            in2 => \_gnd_net_\,
            in3 => \N__43039\,
            lcout => \c0.n453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14639_4_lut_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__50271\,
            in1 => \N__38342\,
            in2 => \N__48410\,
            in3 => \N__42657\,
            lcout => n17416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__42699\,
            in1 => \N__42351\,
            in2 => \N__42462\,
            in3 => \N__43076\,
            lcout => byte_transmit_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10532_2_lut_3_lut_4_lut_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__50733\,
            in1 => \N__38570\,
            in2 => \N__38397\,
            in3 => \N__38662\,
            lcout => \c0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_733_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42961\,
            in1 => \N__42934\,
            in2 => \N__42989\,
            in3 => \N__43075\,
            lcout => n9524,
            ltout => \n9524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_736_LC_13_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__43038\,
            in1 => \N__42844\,
            in2 => \N__38310\,
            in3 => \N__42876\,
            lcout => \c0.n16267\,
            ltout => \c0.n16267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15186_2_lut_3_lut_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__50780\,
            in1 => \_gnd_net_\,
            in2 => \N__38307\,
            in3 => \N__50817\,
            lcout => \c0.n445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10537_2_lut_3_lut_4_lut_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__38560\,
            in1 => \N__50698\,
            in2 => \N__38442\,
            in3 => \N__38636\,
            lcout => \c0.n23_adj_2314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10454_2_lut_3_lut_4_lut_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__38635\,
            in1 => \N__38757\,
            in2 => \N__50723\,
            in3 => \N__38559\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14615_2_lut_4_lut_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__38561\,
            in1 => \N__50699\,
            in2 => \N__48411\,
            in3 => \N__38637\,
            lcout => OPEN,
            ltout => \n17392_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i1_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111011"
        )
    port map (
            in0 => \N__38475\,
            in1 => \N__48032\,
            in2 => \N__38469\,
            in3 => \N__38466\,
            lcout => \UART_TRANSMITTER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10566_2_lut_LC_13_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48021\,
            in2 => \_gnd_net_\,
            in3 => \N__50259\,
            lcout => n2594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10533_2_lut_3_lut_4_lut_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__38568\,
            in1 => \N__50676\,
            in2 => \N__38660\,
            in3 => \N__38505\,
            lcout => \c0.n20_adj_2255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_741_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38675\,
            in1 => \N__38789\,
            in2 => \N__38370\,
            in3 => \N__38453\,
            lcout => OPEN,
            ltout => \c0.n24_adj_2389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_744_LC_13_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38438\,
            in1 => \N__38771\,
            in2 => \N__38427\,
            in3 => \N__38481\,
            lcout => \c0.n26_adj_2391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14552_2_lut_3_lut_LC_13_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__50248\,
            in1 => \N__42845\,
            in2 => \_gnd_net_\,
            in3 => \N__42874\,
            lcout => n17327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_748_LC_13_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38414\,
            in1 => \N__38733\,
            in2 => \N__38393\,
            in3 => \N__38376\,
            lcout => \c0.n9453\,
            ltout => \c0.n9453_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10538_2_lut_3_lut_4_lut_LC_13_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__38369\,
            in1 => \N__50684\,
            in2 => \N__38358\,
            in3 => \N__38567\,
            lcout => \c0.n24_adj_2342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10527_2_lut_3_lut_4_lut_LC_13_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__38569\,
            in1 => \N__50677\,
            in2 => \N__38661\,
            in3 => \N__38790\,
            lcout => \c0.n16_adj_2212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10541_2_lut_3_lut_4_lut_LC_13_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__38772\,
            in1 => \N__38639\,
            in2 => \N__50717\,
            in3 => \N__38566\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_743_LC_13_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38726\,
            in1 => \N__38756\,
            in2 => \N__38712\,
            in3 => \N__38744\,
            lcout => \c0.n22_adj_2390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10531_2_lut_3_lut_4_lut_LC_13_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__38727\,
            in1 => \N__38652\,
            in2 => \N__50744\,
            in3 => \N__38578\,
            lcout => \c0.n18_adj_2220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10522_2_lut_3_lut_4_lut_LC_13_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__38580\,
            in1 => \N__50740\,
            in2 => \N__38663\,
            in3 => \N__38711\,
            lcout => \c0.n15_adj_2211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_13_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__38690\,
            in1 => \N__43290\,
            in2 => \N__44106\,
            in3 => \N__43845\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10528_2_lut_3_lut_4_lut_LC_13_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101010"
        )
    port map (
            in0 => \N__38676\,
            in1 => \N__38653\,
            in2 => \N__50745\,
            in3 => \N__38579\,
            lcout => \c0.n17_adj_2219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_LC_13_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38504\,
            in2 => \_gnd_net_\,
            in3 => \N__38492\,
            lcout => \c0.n18_adj_2388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_i5_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__39711\,
            in1 => \N__39612\,
            in2 => \N__39697\,
            in3 => \N__42094\,
            lcout => \c0.byte_transmit_counter2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49711\,
            ce => 'H',
            sr => \N__39588\
        );

    \c0.rx.r_Rx_Byte_i6_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__45220\,
            in1 => \N__39576\,
            in2 => \N__39523\,
            in3 => \N__45177\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45054\,
            in1 => \N__45315\,
            in2 => \_gnd_net_\,
            in3 => \N__47846\,
            lcout => \c0.n1_adj_2160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i26_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__40567\,
            in1 => \N__39281\,
            in2 => \N__39462\,
            in3 => \N__39395\,
            lcout => \c0.data_in_frame_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14695_4_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011010000"
        )
    port map (
            in0 => \N__39835\,
            in1 => \N__40317\,
            in2 => \N__39258\,
            in3 => \N__40145\,
            lcout => OPEN,
            ltout => \c0.n17472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i7_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__39837\,
            in1 => \N__39951\,
            in2 => \N__39267\,
            in3 => \N__39879\,
            lcout => \c0.data_out_frame2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__2__2275_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39222\,
            in1 => \N__38985\,
            in2 => \_gnd_net_\,
            in3 => \N__38922\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_633_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__39957\,
            in1 => \N__38901\,
            in2 => \N__38853\,
            in3 => \N__38832\,
            lcout => \c0.n21_adj_2357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14713_4_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110000"
        )
    port map (
            in0 => \N__40313\,
            in1 => \N__39831\,
            in2 => \N__40663\,
            in3 => \N__40140\,
            lcout => \c0.n17490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__40598\,
            in1 => \N__40499\,
            in2 => \N__40984\,
            in3 => \N__40431\,
            lcout => \c0.data_in_frame_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14710_4_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010101100"
        )
    port map (
            in0 => \N__40141\,
            in1 => \N__40272\,
            in2 => \N__39844\,
            in3 => \N__40314\,
            lcout => OPEN,
            ltout => \c0.n17487_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i2_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__39836\,
            in1 => \N__39876\,
            in2 => \N__40293\,
            in3 => \N__39947\,
            lcout => \c0.data_out_frame2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15061_3_lut_4_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__41968\,
            in1 => \N__40247\,
            in2 => \N__40089\,
            in3 => \N__40142\,
            lcout => OPEN,
            ltout => \c0.n17690_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame2_0___i3_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__39944\,
            in1 => \N__40079\,
            in2 => \N__40107\,
            in3 => \N__39724\,
            lcout => \c0.data_out_frame2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_622_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40049\,
            in1 => \N__40026\,
            in2 => \_gnd_net_\,
            in3 => \N__39999\,
            lcout => \c0.n17102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n5817_bdd_4_lut_15430_4_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100011111000"
        )
    port map (
            in0 => \N__39943\,
            in1 => \N__39874\,
            in2 => \N__39845\,
            in3 => \N__39759\,
            lcout => \c0.n18202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i29_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41228\,
            in2 => \_gnd_net_\,
            in3 => \N__41552\,
            lcout => \c0.FRAME_MATCHER_state_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49760\,
            ce => 'H',
            sr => \N__41208\
        );

    \c0.FRAME_MATCHER_state_i10_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44975\,
            in1 => \N__44673\,
            in2 => \N__41193\,
            in3 => \N__44510\,
            lcout => \c0.FRAME_MATCHER_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49773\,
            ce => 'H',
            sr => \N__41169\
        );

    \c0.i1_2_lut_adj_488_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41109\,
            lcout => \c0.n17315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_543_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40978\,
            lcout => \c0.n17213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_551_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40933\,
            in2 => \_gnd_net_\,
            in3 => \N__40891\,
            lcout => \c0.n10472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_715_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40820\,
            lcout => \c0.n8_adj_2330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_719_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40759\,
            lcout => \c0.n8_adj_2329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_728_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43150\,
            in2 => \_gnd_net_\,
            in3 => \N__40719\,
            lcout => \c0.n16686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41524\,
            in1 => \N__43264\,
            in2 => \N__43230\,
            in3 => \N__44372\,
            lcout => \c0.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_732_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__41525\,
            in1 => \N__41493\,
            in2 => \N__41420\,
            in3 => \N__41334\,
            lcout => \c0.n16700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i260_2_lut_3_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__42040\,
            in1 => \N__41972\,
            in2 => \_gnd_net_\,
            in3 => \N__41858\,
            lcout => \c0.n276\,
            ltout => \c0.n276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_404_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__41859\,
            in1 => \N__41605\,
            in2 => \N__41559\,
            in3 => \N__44513\,
            lcout => \c0.n4_adj_2135\,
            ltout => \c0.n4_adj_2135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i31_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41529\,
            in3 => \N__41526\,
            lcout => \c0.FRAME_MATCHER_state_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49785\,
            ce => 'H',
            sr => \N__41511\
        );

    \c0.i1_2_lut_4_lut_adj_755_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__44373\,
            in1 => \N__41494\,
            in2 => \N__41421\,
            in3 => \N__41335\,
            lcout => \c0.n16714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_760_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__41336\,
            in1 => \N__41407\,
            in2 => \N__41499\,
            in3 => \N__43265\,
            lcout => \c0.n16690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_761_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__43229\,
            in1 => \N__41498\,
            in2 => \N__41422\,
            in3 => \N__41337\,
            lcout => \c0.n16702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i17_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44978\,
            in1 => \N__44674\,
            in2 => \N__41264\,
            in3 => \N__44600\,
            lcout => \c0.FRAME_MATCHER_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49795\,
            ce => 'H',
            sr => \N__42222\
        );

    \c0.data_out_9__3__2181_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43407\,
            in1 => \N__45620\,
            in2 => \N__46599\,
            in3 => \N__43533\,
            lcout => \c0.data_out_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49805\,
            ce => \N__49970\,
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_463_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__42216\,
            in1 => \N__47488\,
            in2 => \N__47847\,
            in3 => \N__45671\,
            lcout => n10_adj_2431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__3__2173_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__49005\,
            in1 => \N__42177\,
            in2 => \_gnd_net_\,
            in3 => \N__46626\,
            lcout => \c0.data_out_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49805\,
            ce => \N__49970\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_512_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45670\,
            in2 => \_gnd_net_\,
            in3 => \N__46696\,
            lcout => \c0.n6_adj_2221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_437_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42176\,
            in1 => \N__43431\,
            in2 => \N__45696\,
            in3 => \N__48500\,
            lcout => \c0.n15_adj_2177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__0__2200_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__48156\,
            in1 => \N__42168\,
            in2 => \N__50314\,
            in3 => \N__42150\,
            lcout => \c0.data_out_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49812\,
            ce => \N__46934\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_489_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__45398\,
            in1 => \N__42144\,
            in2 => \_gnd_net_\,
            in3 => \N__43313\,
            lcout => \c0.n10183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46506\,
            in1 => \N__47124\,
            in2 => \_gnd_net_\,
            in3 => \N__49111\,
            lcout => \c0.n17129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15405_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42276\,
            in1 => \N__46295\,
            in2 => \N__42309\,
            in3 => \N__47486\,
            lcout => OPEN,
            ltout => \c0.n18184_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18184_bdd_4_lut_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__46296\,
            in1 => \N__42108\,
            in2 => \N__42099\,
            in3 => \N__42270\,
            lcout => OPEN,
            ltout => \n18187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_773_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__46402\,
            in1 => \N__43908\,
            in2 => \N__42327\,
            in3 => \N__46297\,
            lcout => n10_adj_2443,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47256\,
            in1 => \N__42324\,
            in2 => \_gnd_net_\,
            in3 => \N__47812\,
            lcout => \c0.n5_adj_2159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_5__6__2210_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48164\,
            in2 => \_gnd_net_\,
            in3 => \N__42300\,
            lcout => \c0.data_out_7__2__N_447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49820\,
            ce => \N__50567\,
            sr => \N__42793\
        );

    \c0.i15149_2_lut_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47300\,
            in2 => \_gnd_net_\,
            in3 => \N__47811\,
            lcout => \c0.n17698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15119_2_lut_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43284\,
            lcout => \c0.n17612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_452_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45836\,
            in2 => \_gnd_net_\,
            in3 => \N__47873\,
            lcout => \c0.n10395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1__2207_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111011"
        )
    port map (
            in0 => \N__43360\,
            in1 => \N__48303\,
            in2 => \N__42264\,
            in3 => \N__50290\,
            lcout => \c0.data_out_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49827\,
            ce => \N__50548\,
            sr => \_gnd_net_\
        );

    \i51_4_lut_adj_778_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__46294\,
            in1 => \N__46403\,
            in2 => \N__42246\,
            in3 => \N__42678\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9889_3_lut_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48652\,
            in1 => \N__46750\,
            in2 => \_gnd_net_\,
            in3 => \N__47820\,
            lcout => OPEN,
            ltout => \n5_adj_2448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i53_4_lut_adj_776_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__47874\,
            in1 => \N__47821\,
            in2 => \N__42684\,
            in3 => \N__47484\,
            lcout => OPEN,
            ltout => \n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i49_4_lut_adj_777_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__43563\,
            in1 => \N__47485\,
            in2 => \N__42681\,
            in3 => \N__46293\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i146_4_lut_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__42816\,
            in1 => \N__43041\,
            in2 => \N__50722\,
            in3 => \N__42672\,
            lcout => n450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i15099_4_lut_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42642\,
            in1 => \N__43938\,
            in2 => \N__42591\,
            in3 => \N__42554\,
            lcout => OPEN,
            ltout => \c0.tx.n17673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i29_3_lut_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__44179\,
            in1 => \_gnd_net_\,
            in2 => \N__42522\,
            in3 => \N__50823\,
            lcout => \c0.tx.n12_adj_2134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47106\,
            in1 => \N__49084\,
            in2 => \N__42519\,
            in3 => \N__47313\,
            lcout => \c0.n17126\,
            ltout => \c0.n17126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15003_3_lut_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000001010"
        )
    port map (
            in0 => \N__48313\,
            in1 => \_gnd_net_\,
            in2 => \N__42477\,
            in3 => \N__46509\,
            lcout => \c0.n17651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__42735\,
            in1 => \N__42460\,
            in2 => \N__42966\,
            in3 => \N__42365\,
            lcout => byte_transmit_counter_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_2_lut_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44022\,
            in2 => \N__47825\,
            in3 => \_gnd_net_\,
            lcout => \tx_transmit_N_1947_0\,
            ltout => OPEN,
            carryin => \bfn_14_30_0_\,
            carryout => \c0.n16110\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_3_lut_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47483\,
            in2 => \_gnd_net_\,
            in3 => \N__42747\,
            lcout => \tx_transmit_N_1947_1\,
            ltout => OPEN,
            carryin => \c0.n16110\,
            carryout => \c0.n16111\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_4_lut_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46291\,
            in2 => \_gnd_net_\,
            in3 => \N__42744\,
            lcout => \tx_transmit_N_1947_2\,
            ltout => OPEN,
            carryin => \c0.n16111\,
            carryout => \c0.n16112\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_5_lut_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46401\,
            in2 => \_gnd_net_\,
            in3 => \N__42741\,
            lcout => \tx_transmit_N_1947_3\,
            ltout => OPEN,
            carryin => \c0.n16112\,
            carryout => \c0.n16113\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_6_lut_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43836\,
            in2 => \_gnd_net_\,
            in3 => \N__42738\,
            lcout => \tx_transmit_N_1947_4\,
            ltout => OPEN,
            carryin => \c0.n16113\,
            carryout => \c0.n16114\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_7_lut_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42734\,
            in2 => \_gnd_net_\,
            in3 => \N__42723\,
            lcout => \tx_transmit_N_1947_5\,
            ltout => OPEN,
            carryin => \c0.n16114\,
            carryout => \c0.n16115\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_8_lut_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42720\,
            in2 => \_gnd_net_\,
            in3 => \N__42702\,
            lcout => \tx_transmit_N_1947_6\,
            ltout => OPEN,
            carryin => \c0.n16115\,
            carryout => \c0.n16116\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2506_9_lut_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42698\,
            in2 => \_gnd_net_\,
            in3 => \N__42687\,
            lcout => \tx_transmit_N_1947_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_14_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__43043\,
            in1 => \N__43008\,
            in2 => \N__43002\,
            in3 => \N__42875\,
            lcout => OPEN,
            ltout => \c0.n68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_2168_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__48110\,
            in1 => \N__42918\,
            in2 => \N__43080\,
            in3 => \N__43077\,
            lcout => \c0.r_SM_Main_2_N_2034_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__43059\
        );

    \c0.i2_3_lut_adj_766_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__48022\,
            in1 => \N__48314\,
            in2 => \_gnd_net_\,
            in3 => \N__50276\,
            lcout => \c0.n4650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i90_4_lut_LC_14_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110010"
        )
    port map (
            in0 => \N__50275\,
            in1 => \N__43042\,
            in2 => \N__48379\,
            in3 => \N__42842\,
            lcout => \c0.n59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_768_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__42843\,
            in1 => \N__48315\,
            in2 => \_gnd_net_\,
            in3 => \N__50277\,
            lcout => \c0.n65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14627_4_lut_LC_14_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42985\,
            in1 => \N__42962\,
            in2 => \N__50720\,
            in3 => \N__42935\,
            lcout => \c0.n17404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10986_2_lut_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42905\,
            in2 => \_gnd_net_\,
            in3 => \N__42887\,
            lcout => \c0.n13662\,
            ltout => \c0.n13662_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11047_2_lut_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42855\,
            in3 => \N__42841\,
            lcout => \c0.n13726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15194_2_lut_LC_14_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__50322\,
            in1 => \N__50492\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n10815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__3__2253_LC_14_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50323\,
            in2 => \N__50546\,
            in3 => \N__42761\,
            lcout => data_out_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_790_LC_14_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__45330\,
            in1 => \N__46414\,
            in2 => \N__44223\,
            in3 => \N__46292\,
            lcout => n10_adj_2483,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__6__2226_LC_14_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__50319\,
            in1 => \N__48416\,
            in2 => \N__50547\,
            in3 => \N__43280\,
            lcout => \c0.data_out_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i25_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45030\,
            in1 => \N__44737\,
            in2 => \N__43266\,
            in3 => \N__44605\,
            lcout => \c0.FRAME_MATCHER_state_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49749\,
            ce => 'H',
            sr => \N__43242\
        );

    \c0.FRAME_MATCHER_state_i26_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__45029\,
            in1 => \N__43225\,
            in2 => \N__44604\,
            in3 => \N__44738\,
            lcout => \c0.FRAME_MATCHER_state_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49761\,
            ce => 'H',
            sr => \N__43203\
        );

    \c0.FRAME_MATCHER_state_i15_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45018\,
            in1 => \N__44702\,
            in2 => \N__43190\,
            in3 => \N__44573\,
            lcout => \c0.FRAME_MATCHER_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49774\,
            ce => 'H',
            sr => \N__43164\
        );

    \c0.FRAME_MATCHER_state_i21_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__44976\,
            in1 => \N__44678\,
            in2 => \N__43157\,
            in3 => \N__44511\,
            lcout => \c0.FRAME_MATCHER_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49786\,
            ce => 'H',
            sr => \N__43131\
        );

    \c0.FRAME_MATCHER_state_i24_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45028\,
            in1 => \N__44675\,
            in2 => \N__43114\,
            in3 => \N__44583\,
            lcout => \c0.FRAME_MATCHER_state_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49796\,
            ce => 'H',
            sr => \N__43089\
        );

    \c0.data_out_10__4__2172_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43415\,
            in1 => \N__46726\,
            in2 => \_gnd_net_\,
            in3 => \N__47265\,
            lcout => \c0.data_out_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => \N__49980\,
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_421_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43406\,
            in1 => \N__47132\,
            in2 => \N__45843\,
            in3 => \N__45420\,
            lcout => \c0.n17201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__7__2177_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43416\,
            in1 => \N__43491\,
            in2 => \N__43485\,
            in3 => \N__47277\,
            lcout => \c0.data_out_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => \N__49980\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_435_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47536\,
            in2 => \_gnd_net_\,
            in3 => \N__43470\,
            lcout => \c0.n10316\,
            ltout => \c0.n10316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__4__2180_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__43425\,
            in1 => \N__43551\,
            in2 => \N__43419\,
            in3 => \N__45743\,
            lcout => \c0.data_out_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49813\,
            ce => \N__49980\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_731_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47038\,
            in1 => \N__46825\,
            in2 => \N__47199\,
            in3 => \N__47014\,
            lcout => \c0.n17177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43399\,
            in1 => \N__45435\,
            in2 => \_gnd_net_\,
            in3 => \N__47791\,
            lcout => \c0.n8_adj_2157\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_694_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43359\,
            in1 => \N__43398\,
            in2 => \_gnd_net_\,
            in3 => \N__45614\,
            lcout => \c0.n26_adj_2165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9952_3_lut_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43549\,
            in1 => \N__43358\,
            in2 => \_gnd_net_\,
            in3 => \N__47487\,
            lcout => \c0.n12630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_471_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__43320\,
            in1 => \N__47264\,
            in2 => \_gnd_net_\,
            in3 => \N__43624\,
            lcout => \c0.n10179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__1__2255_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__50262\,
            in1 => \N__50537\,
            in2 => \_gnd_net_\,
            in3 => \N__43575\,
            lcout => data_out_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_8__5__2187_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49977\,
            in1 => \N__43743\,
            in2 => \_gnd_net_\,
            in3 => \N__45615\,
            lcout => data_out_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__5__2195_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__43625\,
            in1 => \N__43717\,
            in2 => \N__43650\,
            in3 => \N__46898\,
            lcout => \c0.data_out_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__46176\,
            in1 => \N__43601\,
            in2 => \N__44098\,
            in3 => \N__43844\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43587\,
            in1 => \N__43574\,
            in2 => \_gnd_net_\,
            in3 => \N__47803\,
            lcout => n1_adj_2449,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9953_4_lut_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__47804\,
            in1 => \N__43557\,
            in2 => \N__46832\,
            in3 => \N__47495\,
            lcout => n6_adj_2446,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_453_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43550\,
            in1 => \N__45590\,
            in2 => \N__45464\,
            in3 => \N__43529\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_454_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__49033\,
            in1 => \_gnd_net_\,
            in2 => \N__43518\,
            in3 => \N__48896\,
            lcout => \data_out_9__2__N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__43511\,
            in1 => \N__45750\,
            in2 => \N__44097\,
            in3 => \N__43843\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__47805\,
            in1 => \N__43497\,
            in2 => \N__49040\,
            in3 => \N__47496\,
            lcout => n10_adj_2422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i5_3_lut_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__46051\,
            in1 => \N__45784\,
            in2 => \_gnd_net_\,
            in3 => \N__43851\,
            lcout => OPEN,
            ltout => \c0.tx.n77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i101_4_lut_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45990\,
            in1 => \N__46021\,
            in2 => \N__43899\,
            in3 => \N__46546\,
            lcout => \c0.tx.n83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45522\,
            in2 => \_gnd_net_\,
            in3 => \N__46123\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__45945\,
            in1 => \N__43862\,
            in2 => \_gnd_net_\,
            in3 => \N__43896\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46153\,
            in1 => \N__46084\,
            in2 => \N__45543\,
            in3 => \N__45568\,
            lcout => \c0.tx.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46005\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__43840\,
            in1 => \N__43764\,
            in2 => \N__44075\,
            in3 => \N__43757\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__46124\,
            in1 => \_gnd_net_\,
            in2 => \N__46035\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_402_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43986\,
            in2 => \_gnd_net_\,
            in3 => \N__43936\,
            lcout => \c0.tx.n13702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100010000"
        )
    port map (
            in0 => \N__43937\,
            in1 => \N__45941\,
            in2 => \N__44004\,
            in3 => \N__44115\,
            lcout => \c0.tx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45552\,
            in2 => \_gnd_net_\,
            in3 => \N__46111\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46627\,
            in1 => \N__45838\,
            in2 => \_gnd_net_\,
            in3 => \N__47833\,
            lcout => OPEN,
            ltout => \c0.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_15_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__47834\,
            in1 => \N__48446\,
            in2 => \N__44109\,
            in3 => \N__47494\,
            lcout => n10_adj_2413,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_3_lut_4_lut_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__50819\,
            in1 => \N__44178\,
            in2 => \N__44003\,
            in3 => \N__45940\,
            lcout => n9257,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43985\,
            in2 => \_gnd_net_\,
            in3 => \N__50818\,
            lcout => \c0.tx.n6759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__43999\,
            in1 => \N__45926\,
            in2 => \N__44193\,
            in3 => \N__43952\,
            lcout => \c0.tx.r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_401_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44295\,
            in2 => \_gnd_net_\,
            in3 => \N__50762\,
            lcout => \c0.n65_adj_2192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_4_lut_4_lut_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__43998\,
            in1 => \N__45924\,
            in2 => \N__44191\,
            in3 => \N__43951\,
            lcout => n5142,
            ltout => \n5142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45849\,
            in2 => \N__44313\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_399_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__44310\,
            in1 => \N__44301\,
            in2 => \N__44192\,
            in3 => \N__45925\,
            lcout => \c0.tx.n10613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_2167_LC_15_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50763\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15104_2_lut_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44289\,
            lcout => OPEN,
            ltout => \c0.n17581_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15361_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__44238\,
            in1 => \N__46299\,
            in2 => \N__44226\,
            in3 => \N__47507\,
            lcout => \c0.n18088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__7__2225_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__48112\,
            in1 => \N__50317\,
            in2 => \N__50529\,
            in3 => \N__46530\,
            lcout => data_out_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__44325\,
            in1 => \N__47508\,
            in2 => \N__48687\,
            in3 => \N__47827\,
            lcout => n10_adj_2432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_15_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010001110100"
        )
    port map (
            in0 => \N__44180\,
            in1 => \N__44121\,
            in2 => \N__50781\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_15_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45323\,
            in1 => \N__50007\,
            in2 => \_gnd_net_\,
            in3 => \N__47828\,
            lcout => OPEN,
            ltout => \c0.n2_adj_2164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18088_bdd_4_lut_LC_15_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__45354\,
            in1 => \N__45339\,
            in2 => \N__45333\,
            in3 => \N__46321\,
            lcout => n18091,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__5__2227_LC_15_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__45324\,
            in1 => \N__48113\,
            in2 => \N__50333\,
            in3 => \N__50418\,
            lcout => data_out_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__6__2250_LC_15_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__48383\,
            in1 => \N__50324\,
            in2 => \N__50471\,
            in3 => \N__45308\,
            lcout => \c0.data_out_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__45293\,
            in1 => \N__45259\,
            in2 => \N__45097\,
            in3 => \N__45176\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__6__2242_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__48168\,
            in1 => \N__50291\,
            in2 => \N__50583\,
            in3 => \N__45050\,
            lcout => data_out_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i22_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__45031\,
            in1 => \N__44724\,
            in2 => \N__44371\,
            in3 => \N__44617\,
            lcout => \c0.FRAME_MATCHER_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49814\,
            ce => 'H',
            sr => \N__44349\
        );

    \c0.data_out_1__7__2241_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__50533\,
            in1 => \N__50292\,
            in2 => \_gnd_net_\,
            in3 => \N__44334\,
            lcout => data_out_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15018_2_lut_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__47839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44333\,
            lcout => \c0.n17607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48533\,
            in1 => \N__45616\,
            in2 => \_gnd_net_\,
            in3 => \N__47838\,
            lcout => \c0.n8_adj_2352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__2__2174_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45434\,
            in1 => \N__45509\,
            in2 => \N__46965\,
            in3 => \N__49168\,
            lcout => \c0.data_out_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49829\,
            ce => \N__49988\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_497_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45433\,
            in2 => \_gnd_net_\,
            in3 => \N__45656\,
            lcout => \c0.n17209\,
            ltout => \c0.n17209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__6__2170_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45441\,
            in1 => \N__45494\,
            in2 => \N__45468\,
            in3 => \N__47015\,
            lcout => \c0.data_out_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49829\,
            ce => \N__49988\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_501_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45414\,
            in2 => \_gnd_net_\,
            in3 => \N__45463\,
            lcout => \c0.n6_adj_2216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__6__2178_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__48616\,
            in1 => \N__46574\,
            in2 => \N__48948\,
            in3 => \N__48572\,
            lcout => \c0.data_out_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49829\,
            ce => \N__49988\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_425_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__48571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48615\,
            lcout => \c0.n17200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i51_4_lut_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__47832\,
            in1 => \N__45378\,
            in2 => \N__47195\,
            in3 => \N__47513\,
            lcout => n32,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9896_3_lut_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45413\,
            in1 => \N__48614\,
            in2 => \_gnd_net_\,
            in3 => \N__47831\,
            lcout => n8_adj_2445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i52_3_lut_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45372\,
            in1 => \N__45366\,
            in2 => \_gnd_net_\,
            in3 => \N__46322\,
            lcout => OPEN,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i49_4_lut_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__46323\,
            in1 => \N__45759\,
            in2 => \N__45753\,
            in3 => \N__46415\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_742_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48659\,
            in1 => \N__48926\,
            in2 => \N__48620\,
            in3 => \N__45744\,
            lcout => \c0.n10196\,
            ltout => \c0.n10196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_448_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48447\,
            in2 => \N__45681\,
            in3 => \N__45678\,
            lcout => \c0.n17243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__0__2184_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__45657\,
            in1 => \N__45621\,
            in2 => \N__46662\,
            in3 => \N__45591\,
            lcout => \c0.data_out_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49835\,
            ce => \N__49979\,
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46086\,
            in1 => \N__46085\,
            in2 => \N__45958\,
            in3 => \N__45576\,
            lcout => n10994,
            ltout => OPEN,
            carryin => \bfn_16_28_0_\,
            carryout => \c0.tx.n16117\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45786\,
            in1 => \N__45785\,
            in2 => \N__45963\,
            in3 => \N__45573\,
            lcout => n10951,
            ltout => OPEN,
            carryin => \c0.tx.n16117\,
            carryout => \c0.tx.n16118\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45570\,
            in1 => \N__45569\,
            in2 => \N__45959\,
            in3 => \N__45546\,
            lcout => n10954,
            ltout => OPEN,
            carryin => \c0.tx.n16118\,
            carryout => \c0.tx.n16119\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45542\,
            in1 => \N__45541\,
            in2 => \N__45964\,
            in3 => \N__45516\,
            lcout => n10957,
            ltout => OPEN,
            carryin => \c0.tx.n16119\,
            carryout => \c0.tx.n16120\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46155\,
            in1 => \N__46154\,
            in2 => \N__45960\,
            in3 => \N__46059\,
            lcout => n10960,
            ltout => OPEN,
            carryin => \c0.tx.n16120\,
            carryout => \c0.tx.n16121\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46055\,
            in1 => \N__46056\,
            in2 => \N__45965\,
            in3 => \N__46026\,
            lcout => n10963,
            ltout => OPEN,
            carryin => \c0.tx.n16121\,
            carryout => \c0.tx.n16122\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46023\,
            in1 => \N__46022\,
            in2 => \N__45961\,
            in3 => \N__45996\,
            lcout => n10966,
            ltout => OPEN,
            carryin => \c0.tx.n16122\,
            carryout => \c0.tx.n16123\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46551\,
            in1 => \N__46547\,
            in2 => \N__45966\,
            in3 => \N__45993\,
            lcout => n10969,
            ltout => OPEN,
            carryin => \c0.tx.n16123\,
            carryout => \c0.tx.n16124\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45985\,
            in1 => \N__45986\,
            in2 => \N__45962\,
            in3 => \N__45852\,
            lcout => n10972,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_468_LC_16_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46833\,
            in1 => \N__48971\,
            in2 => \_gnd_net_\,
            in3 => \N__47322\,
            lcout => \c0.n17197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_423_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48683\,
            in2 => \_gnd_net_\,
            in3 => \N__45839\,
            lcout => \c0.n6_adj_2169\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45792\,
            in2 => \_gnd_net_\,
            in3 => \N__46121\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_16_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46122\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45768\,
            lcout => \c0.tx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_16_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47829\,
            in1 => \N__46529\,
            in2 => \_gnd_net_\,
            in3 => \N__46517\,
            lcout => \c0.n2_adj_2156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__7__2233_LC_16_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__46518\,
            in1 => \_gnd_net_\,
            in2 => \N__50470\,
            in3 => \N__50244\,
            lcout => data_out_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15148_2_lut_LC_16_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46508\,
            in2 => \_gnd_net_\,
            in3 => \N__47830\,
            lcout => OPEN,
            ltout => \c0.n17747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_15445_LC_16_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__46449\,
            in1 => \N__46313\,
            in2 => \N__46437\,
            in3 => \N__47509\,
            lcout => OPEN,
            ltout => \c0.n18220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n18220_bdd_4_lut_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__46314\,
            in1 => \N__46434\,
            in2 => \N__46428\,
            in3 => \N__46425\,
            lcout => OPEN,
            ltout => \n18223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_16_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__46416\,
            in1 => \N__46332\,
            in2 => \N__46326\,
            in3 => \N__46315\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_16_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46164\,
            in2 => \_gnd_net_\,
            in3 => \N__46120\,
            lcout => \c0.tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_16_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46134\,
            in2 => \_gnd_net_\,
            in3 => \N__46119\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15208_4_lut_2_lut_3_lut_LC_16_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__48372\,
            in1 => \N__48111\,
            in2 => \_gnd_net_\,
            in3 => \N__50236\,
            lcout => n10596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15202_2_lut_3_lut_LC_16_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__50390\,
            in1 => \N__48382\,
            in2 => \_gnd_net_\,
            in3 => \N__50237\,
            lcout => \c0.n10595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_727_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46704\,
            in1 => \N__48534\,
            in2 => \N__46734\,
            in3 => \N__46766\,
            lcout => \c0.n17252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_479_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46824\,
            in2 => \_gnd_net_\,
            in3 => \N__47016\,
            lcout => OPEN,
            ltout => \c0.n10447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_440_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46788\,
            in1 => \N__48770\,
            in2 => \N__46773\,
            in3 => \N__49014\,
            lcout => \c0.n12_adj_2180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_490_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__46770\,
            in1 => \N__46727\,
            in2 => \_gnd_net_\,
            in3 => \N__46703\,
            lcout => \c0.n17180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_688_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47546\,
            in1 => \N__48826\,
            in2 => \N__47194\,
            in3 => \N__48728\,
            lcout => \c0.n17222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_461_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46658\,
            in1 => \N__48570\,
            in2 => \N__46646\,
            in3 => \N__46589\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_462_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__46578\,
            in1 => \N__48884\,
            in2 => \N__46554\,
            in3 => \N__47331\,
            lcout => \c0.n17261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47048\,
            in1 => \N__48473\,
            in2 => \_gnd_net_\,
            in3 => \N__47840\,
            lcout => OPEN,
            ltout => \c0.n8_adj_2198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__47841\,
            in1 => \N__47547\,
            in2 => \N__47517\,
            in3 => \N__47514\,
            lcout => n10_adj_2430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_457_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48791\,
            in1 => \N__47337\,
            in2 => \_gnd_net_\,
            in3 => \N__49865\,
            lcout => \c0.n17297\,
            ltout => \c0.n17297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_436_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48532\,
            in2 => \N__47325\,
            in3 => \N__47320\,
            lcout => \c0.n14_adj_2176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__0__2176_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47163\,
            in1 => \N__47263\,
            in2 => \N__47211\,
            in3 => \N__46943\,
            lcout => data_out_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49842\,
            ce => \N__49984\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_738_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47162\,
            in1 => \N__47131\,
            in2 => \N__49161\,
            in3 => \N__49113\,
            lcout => \c0.n17162\,
            ltout => \c0.n17162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_466_LC_17_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47058\,
            in1 => \N__47049\,
            in2 => \N__47019\,
            in3 => \N__47013\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__1__2175_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46958\,
            in2 => \N__46947\,
            in3 => \N__46944\,
            lcout => data_out_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49842\,
            ce => \N__49984\,
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_17_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48933\,
            in1 => \N__48903\,
            in2 => \N__48792\,
            in3 => \N__48885\,
            lcout => OPEN,
            ltout => \c0.n10_adj_2166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__1__2183_LC_17_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__48834\,
            in1 => \_gnd_net_\,
            in2 => \N__48795\,
            in3 => \N__48483\,
            lcout => \c0.data_out_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49847\,
            ce => \N__49989\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_455_LC_17_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__48745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48673\,
            lcout => \c0.n10170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_10__5__2171_LC_17_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48774\,
            in1 => \N__48746\,
            in2 => \_gnd_net_\,
            in3 => \N__48732\,
            lcout => \c0.data_out_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49847\,
            ce => \N__49989\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_444_LC_17_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48660\,
            in2 => \_gnd_net_\,
            in3 => \N__48621\,
            lcout => OPEN,
            ltout => \c0.n17150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__5__2179_LC_17_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48591\,
            in1 => \N__48582\,
            in2 => \N__48576\,
            in3 => \N__48566\,
            lcout => \c0.data_out_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49847\,
            ce => \N__49989\,
            sr => \_gnd_net_\
        );

    \c0.data_out_10__7__2169_LC_17_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48510\,
            in2 => \_gnd_net_\,
            in3 => \N__48482\,
            lcout => \c0.data_out_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49847\,
            ce => \N__49989\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__1__2215_LC_17_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__48412\,
            in1 => \N__48134\,
            in2 => \N__47901\,
            in3 => \N__50316\,
            lcout => data_out_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49850\,
            ce => \N__50491\,
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_403_LC_17_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50816\,
            in2 => \_gnd_net_\,
            in3 => \N__50773\,
            lcout => n444,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__5__2235_LC_17_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__50411\,
            in1 => \N__50318\,
            in2 => \_gnd_net_\,
            in3 => \N__50003\,
            lcout => data_out_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_9__2__2182_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49978\,
            in1 => \N__49151\,
            in2 => \_gnd_net_\,
            in3 => \N__49866\,
            lcout => data_out_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_443_LC_18_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49147\,
            in2 => \_gnd_net_\,
            in3 => \N__49112\,
            lcout => OPEN,
            ltout => \c0.n10204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_426_LC_18_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49041\,
            in1 => \N__49013\,
            in2 => \N__48981\,
            in3 => \N__48978\,
            lcout => \c0.n10_adj_2172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
