-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 12 2019 16:24:44

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : inout std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : inout std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : inout std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__35917\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal data_in_10_1 : std_logic;
signal data_in_11_1 : std_logic;
signal data_in_14_1 : std_logic;
signal data_in_13_1 : std_logic;
signal data_in_12_1 : std_logic;
signal data_in_7_4 : std_logic;
signal data_in_8_4 : std_logic;
signal data_in_9_4 : std_logic;
signal data_in_10_4 : std_logic;
signal data_in_11_4 : std_logic;
signal data_in_12_4 : std_logic;
signal data_in_5_1 : std_logic;
signal data_in_6_1 : std_logic;
signal data_in_7_1 : std_logic;
signal data_in_9_1 : std_logic;
signal data_in_8_1 : std_logic;
signal \c0.n4431_cascade_\ : std_logic;
signal n1902 : std_logic;
signal data_in_6_4 : std_logic;
signal \c0.n24_cascade_\ : std_logic;
signal \c0.n4_adj_1594_cascade_\ : std_logic;
signal \c0.n9674_cascade_\ : std_logic;
signal \c0.n9677_cascade_\ : std_logic;
signal \c0.n4431\ : std_logic;
signal \c0.n8849_cascade_\ : std_logic;
signal \c0.n20_adj_1622_cascade_\ : std_logic;
signal \c0.data_in_frame_19_5\ : std_logic;
signal \c0.n10_adj_1637_cascade_\ : std_logic;
signal \c0.data_in_frame_19_3\ : std_logic;
signal \c0.n9686_cascade_\ : std_logic;
signal \c0.n9689_cascade_\ : std_logic;
signal \c0.n10_adj_1646\ : std_logic;
signal \c0.n8779\ : std_logic;
signal \c0.n54_cascade_\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.n9001\ : std_logic;
signal \c0.n9001_cascade_\ : std_logic;
signal \c0.n9464_cascade_\ : std_logic;
signal \c0.n9470_cascade_\ : std_logic;
signal \c0.n9216\ : std_logic;
signal \c0.n9213_cascade_\ : std_logic;
signal \c0.n9210\ : std_logic;
signal \c0.n9458_cascade_\ : std_logic;
signal \c0.n9461_cascade_\ : std_logic;
signal \c0.n9530_cascade_\ : std_logic;
signal \c0.n9524_cascade_\ : std_logic;
signal \c0.n9183\ : std_logic;
signal \c0.n9186_cascade_\ : std_logic;
signal \c0.n9518_cascade_\ : std_logic;
signal \c0.n22_adj_1680\ : std_logic;
signal \c0.n9521_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_0\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal \c0.tx2.n8105\ : std_logic;
signal \c0.tx2.n8106\ : std_logic;
signal \c0.tx2.n8107\ : std_logic;
signal \c0.tx2.n8108\ : std_logic;
signal \c0.tx2.n8109\ : std_logic;
signal \c0.tx2.n8110\ : std_logic;
signal \c0.tx2.n8111\ : std_logic;
signal \c0.tx2.n8112\ : std_logic;
signal \bfn_1_32_0_\ : std_logic;
signal data_in_7_7 : std_logic;
signal data_in_10_7 : std_logic;
signal data_in_11_7 : std_logic;
signal data_in_12_7 : std_logic;
signal data_in_13_4 : std_logic;
signal data_in_14_4 : std_logic;
signal data_in_10_0 : std_logic;
signal data_in_11_0 : std_logic;
signal \c0.n9548_cascade_\ : std_logic;
signal \c0.n9177\ : std_logic;
signal \c0.data_in_field_10\ : std_logic;
signal \c0.n8801_cascade_\ : std_logic;
signal \c0.data_in_field_11\ : std_logic;
signal \c0.n4276\ : std_logic;
signal \c0.n4276_cascade_\ : std_logic;
signal \c0.n12_adj_1633_cascade_\ : std_logic;
signal \c0.n4327\ : std_logic;
signal \c0.n4434_cascade_\ : std_logic;
signal \c0.n8766\ : std_logic;
signal \c0.n9482_cascade_\ : std_logic;
signal \c0.n9207\ : std_logic;
signal n1894 : std_logic;
signal \c0.n9542_cascade_\ : std_logic;
signal \c0.n9180\ : std_logic;
signal \c0.n4114_cascade_\ : std_logic;
signal \c0.n17_cascade_\ : std_logic;
signal \c0.n4324_cascade_\ : std_logic;
signal \c0.n8951\ : std_logic;
signal \c0.n8951_cascade_\ : std_logic;
signal \c0.n48\ : std_logic;
signal \c0.n4406\ : std_logic;
signal \c0.n4406_cascade_\ : std_logic;
signal \c0.n43_adj_1610\ : std_logic;
signal \c0.data_in_frame_20_5\ : std_logic;
signal \c0.n4215_cascade_\ : std_logic;
signal \c0.n18_adj_1593_cascade_\ : std_logic;
signal \c0.n20_adj_1596\ : std_logic;
signal \c0.n4568_cascade_\ : std_logic;
signal \c0.n46\ : std_logic;
signal data_in_6_7 : std_logic;
signal \c0.n8816\ : std_logic;
signal \c0.n4282_cascade_\ : std_logic;
signal \c0.n4577\ : std_logic;
signal \c0.n4282\ : std_logic;
signal \c0.n4476_cascade_\ : std_logic;
signal \c0.n19_adj_1623\ : std_logic;
signal data_in_5_7 : std_logic;
signal tx2_enable : std_logic;
signal \c0.tx2.r_Clock_Count_2\ : std_logic;
signal \c0.tx2.r_Clock_Count_6\ : std_logic;
signal \c0.tx2.r_Clock_Count_1\ : std_logic;
signal \c0.tx2.r_Clock_Count_3\ : std_logic;
signal \c0.tx2.r_Clock_Count_4\ : std_logic;
signal \c0.tx2.r_Clock_Count_5\ : std_logic;
signal \c0.tx2.n5_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_7\ : std_logic;
signal \c0.tx2.n4081\ : std_logic;
signal \c0.tx2.n4081_cascade_\ : std_logic;
signal \c0.tx2.n7\ : std_logic;
signal \c0.tx2.n8196_cascade_\ : std_logic;
signal \c0.tx2.n5146\ : std_logic;
signal \n9075_cascade_\ : std_logic;
signal \c0.tx2.r_Clock_Count_8\ : std_logic;
signal \c0.tx2.n7399\ : std_logic;
signal \c0.tx2.n7236\ : std_logic;
signal \c0.tx2.n7236_cascade_\ : std_logic;
signal \n3220_cascade_\ : std_logic;
signal data_in_9_7 : std_logic;
signal data_in_8_7 : std_logic;
signal n1900 : std_logic;
signal data_in_7_3 : std_logic;
signal data_in_8_3 : std_logic;
signal data_in_9_0 : std_logic;
signal data_in_8_0 : std_logic;
signal data_in_7_0 : std_logic;
signal data_in_1_5 : std_logic;
signal data_in_12_0 : std_logic;
signal \c0.n14_adj_1670\ : std_logic;
signal \c0.n14_adj_1669\ : std_logic;
signal \c0.n26_adj_1673\ : std_logic;
signal \c0.n25_adj_1675\ : std_logic;
signal \c0.n9033_cascade_\ : std_logic;
signal \c0.n9578\ : std_logic;
signal \c0.n8794\ : std_logic;
signal data_in_3_1 : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n4381\ : std_logic;
signal \c0.n4381_cascade_\ : std_logic;
signal \c0.data_in_field_20\ : std_logic;
signal data_in_4_1 : std_logic;
signal \c0.data_in_field_35\ : std_logic;
signal \c0.n4154_cascade_\ : std_logic;
signal \c0.data_in_field_19\ : std_logic;
signal \c0.n14\ : std_logic;
signal \c0.n10_adj_1631_cascade_\ : std_logic;
signal data_in_1_1 : std_logic;
signal data_in_4_7 : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.data_in_field_4\ : std_logic;
signal data_in_0_7 : std_logic;
signal \c0.n8776\ : std_logic;
signal \c0.n4131_cascade_\ : std_logic;
signal \c0.n8927_cascade_\ : std_logic;
signal n1896 : std_logic;
signal data_in_2_7 : std_logic;
signal data_in_0_6 : std_logic;
signal \c0.n10_adj_1647_cascade_\ : std_logic;
signal \c0.data_in_frame_19_1\ : std_logic;
signal \c0.n9704_cascade_\ : std_logic;
signal \c0.data_in_frame_20_1\ : std_logic;
signal \c0.n9707_cascade_\ : std_logic;
signal \c0.n22_adj_1682\ : std_logic;
signal \c0.n9722_cascade_\ : std_logic;
signal \c0.data_in_field_7\ : std_logic;
signal \c0.data_in_field_23\ : std_logic;
signal \c0.n4514\ : std_logic;
signal \c0.n9007\ : std_logic;
signal \c0.n18_adj_1589_cascade_\ : std_logic;
signal \c0.n20_adj_1590_cascade_\ : std_logic;
signal \c0.n29\ : std_logic;
signal \c0.n4114\ : std_logic;
signal \c0.n4448\ : std_logic;
signal \c0.n4445\ : std_logic;
signal \c0.n8896\ : std_logic;
signal n6164 : std_logic;
signal data_in_field_105 : std_logic;
signal \c0.n8890_cascade_\ : std_logic;
signal \c0.n14_adj_1638\ : std_logic;
signal \c0.n4285\ : std_logic;
signal data_in_field_83 : std_logic;
signal \c0.n9126\ : std_logic;
signal \c0.n9123_cascade_\ : std_logic;
signal \c0.n9240\ : std_logic;
signal \c0.n9644_cascade_\ : std_logic;
signal \c0.n9647_cascade_\ : std_logic;
signal \c0.n9656\ : std_logic;
signal \c0.n9752_cascade_\ : std_logic;
signal \c0.data_in_field_39\ : std_logic;
signal \c0.n9120\ : std_logic;
signal \c0.tx2.r_Tx_Data_3\ : std_logic;
signal \c0.tx2.r_Tx_Data_1\ : std_logic;
signal \c0.tx2.n9692_cascade_\ : std_logic;
signal \c0.tx2.n9695_cascade_\ : std_logic;
signal \c0.tx2.o_Tx_Serial_N_1511_cascade_\ : std_logic;
signal \n2207_cascade_\ : std_logic;
signal \r_Bit_Index_2_adj_1741\ : std_logic;
signal \r_SM_Main_0_adj_1740\ : std_logic;
signal \r_SM_Main_2_N_1480_1_adj_1744\ : std_logic;
signal data_in_13_7 : std_logic;
signal data_in_16_6 : std_logic;
signal data_in_9_6 : std_logic;
signal data_in_10_6 : std_logic;
signal data_in_11_6 : std_logic;
signal data_in_13_6 : std_logic;
signal data_in_12_6 : std_logic;
signal data_in_15_6 : std_logic;
signal data_in_14_6 : std_logic;
signal data_in_20_4 : std_logic;
signal data_in_3_0 : std_logic;
signal data_in_0_5 : std_logic;
signal \c0.n28_adj_1668_cascade_\ : std_logic;
signal \c0.n30_adj_1674\ : std_logic;
signal \c0.n22_adj_1667\ : std_logic;
signal data_in_0_0 : std_logic;
signal data_in_13_0 : std_logic;
signal data_in_4_0 : std_logic;
signal \c0.n13_adj_1671\ : std_logic;
signal \c0.n13_adj_1672\ : std_logic;
signal data_in_1_2 : std_logic;
signal data_in_6_3 : std_logic;
signal data_in_1_3 : std_logic;
signal data_in_2_3 : std_logic;
signal \c0.n4495\ : std_logic;
signal \c0.data_in_field_2\ : std_logic;
signal \c0.data_in_field_33\ : std_logic;
signal \c0.n6_adj_1632_cascade_\ : std_logic;
signal \c0.n8804\ : std_logic;
signal data_in_1_6 : std_logic;
signal data_in_3_7 : std_logic;
signal \c0.n4127\ : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.data_in_field_3\ : std_logic;
signal \c0.n20_adj_1597\ : std_logic;
signal \c0.n22_adj_1595\ : std_logic;
signal data_in_2_6 : std_logic;
signal \n9069_cascade_\ : std_logic;
signal data_in_3_3 : std_logic;
signal \c0.n8849\ : std_logic;
signal \n4_adj_1750_cascade_\ : std_logic;
signal n1892 : std_logic;
signal n1891 : std_logic;
signal \c0.n8831\ : std_logic;
signal \c0.data_in_field_9\ : std_logic;
signal \c0.n8831_cascade_\ : std_logic;
signal data_in_1_0 : std_logic;
signal n1888 : std_logic;
signal data_in_5_3 : std_logic;
signal data_in_4_3 : std_logic;
signal \c0.n4131\ : std_logic;
signal \c0.n4224\ : std_logic;
signal \c0.n10_adj_1640_cascade_\ : std_logic;
signal \c0.n4434\ : std_logic;
signal \c0.n8933_cascade_\ : std_logic;
signal \c0.n8822\ : std_logic;
signal \c0.n8314_cascade_\ : std_logic;
signal data_in_field_145 : std_logic;
signal \c0.n4556\ : std_logic;
signal \c0.n8861\ : std_logic;
signal \c0.n6\ : std_logic;
signal \c0.n4452_cascade_\ : std_logic;
signal \c0.n8906\ : std_logic;
signal \c0.n4452\ : std_logic;
signal \c0.n4253_cascade_\ : std_logic;
signal data_in_field_71 : std_logic;
signal data_in_field_147 : std_logic;
signal data_in_field_127 : std_logic;
signal \c0.n9650\ : std_logic;
signal \c0.n16_adj_1598\ : std_logic;
signal \c0.n9016\ : std_logic;
signal \c0.n6_adj_1645_cascade_\ : std_logic;
signal \c0.n4154\ : std_logic;
signal \c0.n8788_cascade_\ : std_logic;
signal \c0.n14_adj_1648\ : std_logic;
signal \c0.n8936\ : std_logic;
signal \c0.n24_adj_1600_cascade_\ : std_logic;
signal \c0.n18_adj_1603\ : std_logic;
signal \c0.n4107\ : std_logic;
signal \c0.tx2_transmit_N_1334_cascade_\ : std_logic;
signal \c0.n8980\ : std_logic;
signal \c0.n22_adj_1601_cascade_\ : std_logic;
signal \c0.n26\ : std_logic;
signal \c0.n16\ : std_logic;
signal data_in_field_115 : std_logic;
signal \c0.n4574_cascade_\ : std_logic;
signal data_in_field_81 : std_logic;
signal data_in_field_47 : std_logic;
signal \c0.n4333\ : std_logic;
signal \c0.n4333_cascade_\ : std_logic;
signal n3_adj_1749 : std_logic;
signal tx2_o : std_logic;
signal \c0.n24_adj_1615\ : std_logic;
signal \c0.n34\ : std_logic;
signal \r_SM_Main_1_adj_1739\ : std_logic;
signal n8747 : std_logic;
signal \c0.tx2.r_Tx_Data_7\ : std_logic;
signal \c0.tx2.n9716_cascade_\ : std_logic;
signal \c0.tx2.n9719\ : std_logic;
signal \n4691_cascade_\ : std_logic;
signal \r_Bit_Index_0_adj_1743\ : std_logic;
signal n9075 : std_logic;
signal n5346 : std_logic;
signal \r_Bit_Index_1_adj_1742\ : std_logic;
signal data_in_15_1 : std_logic;
signal data_in_5_4 : std_logic;
signal data_in_17_1 : std_logic;
signal data_in_16_1 : std_logic;
signal data_in_14_7 : std_logic;
signal data_in_15_7 : std_logic;
signal data_in_16_7 : std_logic;
signal data_in_15_4 : std_logic;
signal data_in_17_4 : std_logic;
signal data_in_16_4 : std_logic;
signal data_in_17_7 : std_logic;
signal data_in_19_4 : std_logic;
signal data_in_18_4 : std_logic;
signal data_in_2_5 : std_logic;
signal data_in_5_6 : std_logic;
signal data_in_4_6 : std_logic;
signal data_in_6_6 : std_logic;
signal data_in_8_6 : std_logic;
signal data_in_7_6 : std_logic;
signal data_in_3_5 : std_logic;
signal data_in_3_6 : std_logic;
signal \c0.n8843_cascade_\ : std_logic;
signal \c0.data_in_field_31\ : std_logic;
signal \c0.n4151_cascade_\ : std_logic;
signal \c0.data_in_field_30\ : std_logic;
signal \c0.data_in_field_22\ : std_logic;
signal \c0.data_in_field_14\ : std_logic;
signal \c0.n9638_cascade_\ : std_logic;
signal \c0.data_in_field_6\ : std_logic;
signal data_in_2_0 : std_logic;
signal \c0.data_in_field_26\ : std_logic;
signal \c0.data_in_field_18\ : std_logic;
signal \c0.n9512\ : std_logic;
signal data_in_2_1 : std_logic;
signal \c0.n4492\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.n8902\ : std_logic;
signal \c0.n4492_cascade_\ : std_logic;
signal \c0.n8948_cascade_\ : std_logic;
signal \c0.n8858\ : std_logic;
signal \c0.n19_adj_1602\ : std_logic;
signal data_in_0_1 : std_logic;
signal \c0.data_in_field_1\ : std_logic;
signal data_in_1_7 : std_logic;
signal \c0.data_in_field_15\ : std_logic;
signal \n1895_cascade_\ : std_logic;
signal n1889 : std_logic;
signal n1897 : std_logic;
signal data_in_4_4 : std_logic;
signal \c0.n9506_cascade_\ : std_logic;
signal \c0.data_in_field_34\ : std_logic;
signal \c0.n4_adj_1592_cascade_\ : std_logic;
signal \c0.n4324\ : std_logic;
signal \c0.n21_adj_1599\ : std_logic;
signal \c0.n4200\ : std_logic;
signal \c0.n28\ : std_logic;
signal \c0.n23_adj_1608\ : std_logic;
signal \c0.n8864\ : std_logic;
signal \c0.n8843\ : std_logic;
signal \c0.n8930\ : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.n21_cascade_\ : std_logic;
signal \c0.n19\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n8421_cascade_\ : std_logic;
signal \c0.tx2_transmit_N_1334\ : std_logic;
signal \c0.n24_adj_1605\ : std_logic;
signal data_in_field_75 : std_logic;
signal data_in_field_67 : std_logic;
signal \c0.n6_adj_1654\ : std_logic;
signal \c0.n4253\ : std_logic;
signal \c0.n4151\ : std_logic;
signal \c0.data_in_field_17\ : std_logic;
signal \c0.n45\ : std_logic;
signal \c0.n4183\ : std_logic;
signal data_in_field_63 : std_logic;
signal data_in_field_59 : std_logic;
signal data_in_field_51 : std_logic;
signal \c0.n4302\ : std_logic;
signal data_in_field_79 : std_logic;
signal data_in_field_139 : std_logic;
signal \c0.n8825\ : std_logic;
signal data_in_field_111 : std_logic;
signal \c0.n4525_cascade_\ : std_logic;
signal data_in_field_107 : std_logic;
signal data_in_field_137 : std_logic;
signal \c0.n8874_cascade_\ : std_logic;
signal data_in_field_55 : std_logic;
signal \c0.n6_adj_1636\ : std_logic;
signal \c0.n8989\ : std_logic;
signal \c0.n6_adj_1604_cascade_\ : std_logic;
signal \c0.n8983\ : std_logic;
signal \c0.n8948\ : std_logic;
signal \c0.n8945\ : std_logic;
signal \c0.n8983_cascade_\ : std_logic;
signal \c0.n9004\ : std_logic;
signal data_in_field_89 : std_logic;
signal \c0.n4203\ : std_logic;
signal \c0.n8890\ : std_logic;
signal \c0.n8874\ : std_logic;
signal \c0.n24_adj_1607\ : std_logic;
signal \c0.n23\ : std_logic;
signal \c0.n25_cascade_\ : std_logic;
signal \c0.n26_adj_1606\ : std_logic;
signal \c0.data_in_frame_20_3\ : std_logic;
signal \c0.n8974\ : std_logic;
signal \c0.n22_adj_1617\ : std_logic;
signal \c0.n8933\ : std_logic;
signal \c0.data_in_frame_20_7\ : std_logic;
signal \c0.n3056_cascade_\ : std_logic;
signal \c0.n22_adj_1676\ : std_logic;
signal \c0.n38_adj_1616\ : std_logic;
signal \c0.n36\ : std_logic;
signal \c0.n37\ : std_logic;
signal \c0.data_in_frame_19_7\ : std_logic;
signal data_in_field_135 : std_logic;
signal \c0.n9662_cascade_\ : std_logic;
signal \c0.n9665\ : std_logic;
signal data_in_13_3 : std_logic;
signal data_in_14_3 : std_logic;
signal data_in_16_3 : std_logic;
signal data_in_15_3 : std_logic;
signal data_in_17_3 : std_logic;
signal data_in_18_3 : std_logic;
signal data_in_19_3 : std_logic;
signal data_in_20_3 : std_logic;
signal data_in_19_5 : std_logic;
signal data_in_17_6 : std_logic;
signal data_in_10_3 : std_logic;
signal data_in_9_3 : std_logic;
signal data_in_20_5 : std_logic;
signal data_in_5_5 : std_logic;
signal data_in_4_5 : std_logic;
signal data_in_6_5 : std_logic;
signal data_in_7_5 : std_logic;
signal data_in_8_5 : std_logic;
signal data_in_9_5 : std_logic;
signal data_in_14_0 : std_logic;
signal data_in_15_0 : std_logic;
signal data_in_2_2 : std_logic;
signal data_in_16_0 : std_logic;
signal data_in_20_0 : std_logic;
signal n1898 : std_logic;
signal \c0.n9746_cascade_\ : std_logic;
signal \c0.data_in_field_32\ : std_logic;
signal data_in_field_42 : std_logic;
signal data_in_field_40 : std_logic;
signal \c0.n4208\ : std_logic;
signal data_in_3_4 : std_logic;
signal data_in_3_2 : std_logic;
signal data_in_2_4 : std_logic;
signal data_in_17_0 : std_logic;
signal \c0.n8960\ : std_logic;
signal data_in_0_4 : std_logic;
signal n1890 : std_logic;
signal data_in_1_4 : std_logic;
signal n9069 : std_logic;
signal data_in_field_45 : std_logic;
signal \c0.n9602\ : std_logic;
signal \c0.data_in_field_12\ : std_logic;
signal \c0.n9019\ : std_logic;
signal \c0.data_in_field_28\ : std_logic;
signal n9091 : std_logic;
signal \n9092_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal n8761 : std_logic;
signal data_in_field_48 : std_logic;
signal \c0.n4897_cascade_\ : std_logic;
signal \bfn_6_27_0_\ : std_logic;
signal n8155 : std_logic;
signal n8156 : std_logic;
signal n8157 : std_logic;
signal n8158 : std_logic;
signal rand_data_5 : std_logic;
signal n8159 : std_logic;
signal n8160 : std_logic;
signal n8161 : std_logic;
signal n8162 : std_logic;
signal \bfn_6_28_0_\ : std_logic;
signal n8163 : std_logic;
signal n8164 : std_logic;
signal n8165 : std_logic;
signal n8166 : std_logic;
signal n8167 : std_logic;
signal rand_data_14 : std_logic;
signal n8168 : std_logic;
signal n8169 : std_logic;
signal n8170 : std_logic;
signal \bfn_6_29_0_\ : std_logic;
signal n8171 : std_logic;
signal n8172 : std_logic;
signal rand_data_19 : std_logic;
signal n8173 : std_logic;
signal n8174 : std_logic;
signal n8175 : std_logic;
signal n8176 : std_logic;
signal n8177 : std_logic;
signal n8178 : std_logic;
signal \bfn_6_30_0_\ : std_logic;
signal rand_data_25 : std_logic;
signal n8179 : std_logic;
signal n8180 : std_logic;
signal rand_data_27 : std_logic;
signal n8181 : std_logic;
signal n8182 : std_logic;
signal n8183 : std_logic;
signal n8184 : std_logic;
signal n8185 : std_logic;
signal rand_data_31 : std_logic;
signal data_in_field_104 : std_logic;
signal \c0.n9734_cascade_\ : std_logic;
signal data_in_field_141 : std_logic;
signal rand_data_21 : std_logic;
signal rand_data_17 : std_logic;
signal data_in_field_113 : std_logic;
signal data_in_field_149 : std_logic;
signal \c0.n1893_adj_1635\ : std_logic;
signal rand_data_23 : std_logic;
signal data_in_field_85 : std_logic;
signal \c0.n9596_cascade_\ : std_logic;
signal data_in_field_117 : std_logic;
signal \c0.n9590_cascade_\ : std_logic;
signal \c0.n9153\ : std_logic;
signal \c0.n9156_cascade_\ : std_logic;
signal \c0.n9584_cascade_\ : std_logic;
signal \c0.n9150\ : std_logic;
signal \c0.n22_adj_1678\ : std_logic;
signal \c0.n9587_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_5\ : std_logic;
signal data_in_10_5 : std_logic;
signal data_in_11_5 : std_logic;
signal data_in_13_5 : std_logic;
signal data_in_12_5 : std_logic;
signal data_in_14_5 : std_logic;
signal data_in_15_5 : std_logic;
signal data_in_16_5 : std_logic;
signal data_in_18_5 : std_logic;
signal data_in_17_5 : std_logic;
signal data_in_18_6 : std_logic;
signal data_in_18_1 : std_logic;
signal data_in_19_1 : std_logic;
signal data_in_20_1 : std_logic;
signal rx_data_2 : std_logic;
signal data_in_12_3 : std_logic;
signal data_in_11_3 : std_logic;
signal n4 : std_logic;
signal rx_data_3 : std_logic;
signal data_in_19_6 : std_logic;
signal rx_data_0 : std_logic;
signal data_in_18_7 : std_logic;
signal data_in_20_6 : std_logic;
signal n4_adj_1725 : std_logic;
signal \n4_adj_1725_cascade_\ : std_logic;
signal rx_data_1 : std_logic;
signal \n4044_cascade_\ : std_logic;
signal rx_data_6 : std_logic;
signal rx_data_4 : std_logic;
signal rx_data_7 : std_logic;
signal data_in_20_7 : std_logic;
signal data_in_19_7 : std_logic;
signal n4044 : std_logic;
signal rx_data_5 : std_logic;
signal n4049 : std_logic;
signal \c0.n9476\ : std_logic;
signal rand_data_24 : std_logic;
signal n1903 : std_logic;
signal data_in_field_129 : std_logic;
signal \c0.n8791\ : std_logic;
signal data_in_6_0 : std_logic;
signal data_in_5_0 : std_logic;
signal \c0.n19_adj_1665_cascade_\ : std_logic;
signal tx2_active : std_logic;
signal \c0.r_SM_Main_2_N_1483_0\ : std_logic;
signal \c0.n19_adj_1665\ : std_logic;
signal \c0.n7194_cascade_\ : std_logic;
signal \c0.n8449\ : std_logic;
signal n4839 : std_logic;
signal \n4839_cascade_\ : std_logic;
signal n31 : std_logic;
signal data_in_field_65 : std_logic;
signal \c0.tx2_transmit_N_1444\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \c0.n8113\ : std_logic;
signal \c0.n8114\ : std_logic;
signal \c0.n8115\ : std_logic;
signal \c0.n8116\ : std_logic;
signal \c0.byte_transmit_counter2_5\ : std_logic;
signal \c0.n8117\ : std_logic;
signal \c0.byte_transmit_counter2_6\ : std_logic;
signal \c0.n8118\ : std_logic;
signal \c0.n8119\ : std_logic;
signal \c0.byte_transmit_counter2_7\ : std_logic;
signal \c0.n4897\ : std_logic;
signal \c0.n5154\ : std_logic;
signal rand_data_8 : std_logic;
signal rand_data_22 : std_logic;
signal rand_data_3 : std_logic;
signal \c0.n8992\ : std_logic;
signal \c0.n21_adj_1624\ : std_logic;
signal rand_data_7 : std_logic;
signal rand_data_1 : std_logic;
signal rand_data_15 : std_logic;
signal data_in_field_143 : std_logic;
signal rand_data_28 : std_logic;
signal rand_data_13 : std_logic;
signal \c0.data_in_field_29\ : std_logic;
signal \c0.data_in_field_21\ : std_logic;
signal \c0.n9608_cascade_\ : std_logic;
signal \c0.data_in_field_5\ : std_logic;
signal \c0.n9147\ : std_logic;
signal rand_data_29 : std_logic;
signal data_in_field_109 : std_logic;
signal rand_data_4 : std_logic;
signal \c0.n8942\ : std_logic;
signal data_in_field_57 : std_logic;
signal data_in_field_93 : std_logic;
signal \c0.n4390\ : std_logic;
signal data_in_field_87 : std_logic;
signal data_in_field_91 : std_logic;
signal \c0.n8909\ : std_logic;
signal \c0.n4197\ : std_logic;
signal data_in_field_60 : std_logic;
signal \c0.n4197_cascade_\ : std_logic;
signal \c0.n4399\ : std_logic;
signal data_in_field_61 : std_logic;
signal \c0.n4399_cascade_\ : std_logic;
signal \c0.n4288\ : std_logic;
signal \c0.n10\ : std_logic;
signal rand_data_9 : std_logic;
signal data_in_field_121 : std_logic;
signal data_in_field_44 : std_logic;
signal \c0.n9572\ : std_logic;
signal data_in_field_77 : std_logic;
signal data_in_field_49 : std_logic;
signal \c0.n8887_cascade_\ : std_logic;
signal data_in_field_120 : std_logic;
signal rand_data_30 : std_logic;
signal \c0.n8785\ : std_logic;
signal \c0.n8887\ : std_logic;
signal \c0.n4240_cascade_\ : std_logic;
signal \c0.data_in_field_13\ : std_logic;
signal \c0.n44_adj_1609\ : std_logic;
signal \c0.n4553\ : std_logic;
signal data_in_field_53 : std_logic;
signal \c0.n8964\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \c0.n18_adj_1666\ : std_logic;
signal data_in_field_36 : std_logic;
signal \c0.n1645\ : std_logic;
signal data_in_field_62 : std_logic;
signal data_in_field_46 : std_logic;
signal \c0.n9632_cascade_\ : std_logic;
signal \c0.data_in_field_38\ : std_logic;
signal data_in_field_126 : std_logic;
signal \c0.n9620_cascade_\ : std_logic;
signal data_in_field_94 : std_logic;
signal \c0.n9626_cascade_\ : std_logic;
signal \c0.n9141\ : std_logic;
signal \c0.n9138_cascade_\ : std_logic;
signal \c0.n9132\ : std_logic;
signal \c0.n9135\ : std_logic;
signal \c0.n9614_cascade_\ : std_logic;
signal \c0.n9617_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_6\ : std_logic;
signal data_in_11_2 : std_logic;
signal data_in_12_2 : std_logic;
signal data_in_13_2 : std_logic;
signal data_in_14_2 : std_logic;
signal data_in_15_2 : std_logic;
signal data_in_16_2 : std_logic;
signal data_in_18_2 : std_logic;
signal data_in_17_2 : std_logic;
signal data_in_20_2 : std_logic;
signal data_in_19_2 : std_logic;
signal n7171 : std_logic;
signal \c0.n9668\ : std_logic;
signal \c0.n8878\ : std_logic;
signal \c0.n8813\ : std_logic;
signal data_in_field_43 : std_logic;
signal \c0.n28_adj_1619\ : std_logic;
signal \c0.n29_adj_1620_cascade_\ : std_logic;
signal \c0.data_in_frame_19_6\ : std_logic;
signal n1901 : std_logic;
signal \FRAME_MATCHER_state_2\ : std_logic;
signal \c0.n7194\ : std_logic;
signal n9262 : std_logic;
signal data_in_6_2 : std_logic;
signal \FRAME_MATCHER_state_0\ : std_logic;
signal n1893 : std_logic;
signal data_in_7_2 : std_logic;
signal data_in_8_2 : std_logic;
signal data_in_10_2 : std_logic;
signal data_in_9_2 : std_logic;
signal \c0.n8921\ : std_logic;
signal \c0.n4562_cascade_\ : std_logic;
signal \c0.n4479\ : std_logic;
signal \c0.n4235_cascade_\ : std_logic;
signal \c0.n4562\ : std_logic;
signal data_in_field_99 : std_logic;
signal data_in_field_131 : std_logic;
signal \c0.n8846\ : std_logic;
signal rand_data_2 : std_logic;
signal \c0.n30\ : std_logic;
signal rand_data_26 : std_logic;
signal data_in_field_58 : std_logic;
signal data_in_field_118 : std_logic;
signal \c0.n4534\ : std_logic;
signal \c0.n27_adj_1621\ : std_logic;
signal rand_data_10 : std_logic;
signal \c0.n4473\ : std_logic;
signal \c0.n4473_cascade_\ : std_logic;
signal \c0.n9010\ : std_logic;
signal \c0.n4244_cascade_\ : std_logic;
signal rand_data_6 : std_logic;
signal data_in_field_102 : std_logic;
signal data_in_field_125 : std_logic;
signal data_in_field_73 : std_logic;
signal \c0.n18_adj_1618\ : std_logic;
signal data_in_field_54 : std_logic;
signal data_in_field_69 : std_logic;
signal \c0.n8998\ : std_logic;
signal \c0.n16_adj_1591\ : std_logic;
signal rand_data_20 : std_logic;
signal data_in_field_124 : std_logic;
signal data_in_field_116 : std_logic;
signal data_in_field_56 : std_logic;
signal data_in_field_101 : std_logic;
signal rand_data_16 : std_logic;
signal \c0.n8788\ : std_logic;
signal \c0.n8828\ : std_logic;
signal \c0.n8855\ : std_logic;
signal \c0.n35\ : std_logic;
signal data_in_field_84 : std_logic;
signal data_in_field_92 : std_logic;
signal \c0.n9560\ : std_logic;
signal data_in_field_108 : std_logic;
signal data_in_field_100 : std_logic;
signal \c0.n8927\ : std_logic;
signal \c0.n8837\ : std_logic;
signal data_in_field_41 : std_logic;
signal \c0.n16_adj_1629\ : std_logic;
signal \c0.n8977\ : std_logic;
signal \c0.n17_adj_1630\ : std_logic;
signal \c0.data_in_frame_19_4\ : std_logic;
signal \c0.data_in_frame_20_4\ : std_logic;
signal data_in_field_68 : std_logic;
signal data_in_field_76 : std_logic;
signal \c0.n9566\ : std_logic;
signal \c0.n9171\ : std_logic;
signal \c0.n9168_cascade_\ : std_logic;
signal \c0.n9165\ : std_logic;
signal \c0.n9162\ : std_logic;
signal \c0.n9554\ : std_logic;
signal \c0.n22_adj_1679\ : std_logic;
signal \c0.n9557_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_Data_4\ : std_logic;
signal \n5185_cascade_\ : std_logic;
signal data_in_field_150 : std_logic;
signal data_in_field_52 : std_logic;
signal data_in_field_151 : std_logic;
signal data_in_field_86 : std_logic;
signal \c0.n8915\ : std_logic;
signal n9077 : std_logic;
signal n5185 : std_logic;
signal \r_Bit_Index_0_adj_1733\ : std_logic;
signal \r_Bit_Index_1_adj_1732\ : std_logic;
signal n4_adj_1724 : std_logic;
signal data_in_field_134 : std_logic;
signal data_in_field_119 : std_logic;
signal \c0.n8883\ : std_logic;
signal \c0.n8770\ : std_logic;
signal \c0.n8810\ : std_logic;
signal \c0.n8899\ : std_logic;
signal \c0.n16_adj_1657\ : std_logic;
signal \c0.n22_adj_1655_cascade_\ : std_logic;
signal data_in_field_37 : std_logic;
signal \c0.n24_adj_1658\ : std_logic;
signal \c0.n8939\ : std_logic;
signal \c0.n20_adj_1659\ : std_logic;
signal \c0.data_in_frame_19_0\ : std_logic;
signal data_in_field_136 : std_logic;
signal \c0.n9536_cascade_\ : std_logic;
signal data_in_field_128 : std_logic;
signal \c0.n9539_cascade_\ : std_logic;
signal rand_data_18 : std_logic;
signal data_in_field_114 : std_logic;
signal data_in_field_144 : std_logic;
signal \c0.n8971\ : std_logic;
signal \c0.n6_adj_1628\ : std_logic;
signal rand_data_0 : std_logic;
signal \c0.n8918\ : std_logic;
signal \c0.n8840_cascade_\ : std_logic;
signal \c0.n4511\ : std_logic;
signal \c0.n4309\ : std_logic;
signal rand_data_11 : std_logic;
signal data_in_field_123 : std_logic;
signal data_in_field_146 : std_logic;
signal data_in_field_130 : std_logic;
signal \c0.n9698_cascade_\ : std_logic;
signal data_in_field_138 : std_logic;
signal \c0.n9701_cascade_\ : std_logic;
signal data_in_field_142 : std_logic;
signal data_in_field_78 : std_logic;
signal \c0.n4215\ : std_logic;
signal \c0.n8912\ : std_logic;
signal \c0.n8954\ : std_logic;
signal \c0.n8819_cascade_\ : std_logic;
signal \c0.n4365\ : std_logic;
signal \c0.n21_adj_1644_cascade_\ : std_logic;
signal \c0.n19_adj_1643\ : std_logic;
signal \c0.data_in_frame_19_2\ : std_logic;
signal \c0.n8782\ : std_logic;
signal \c0.n8807\ : std_logic;
signal data_in_field_110 : std_logic;
signal \c0.n8819\ : std_logic;
signal \c0.n8893\ : std_logic;
signal \c0.n8427\ : std_logic;
signal \c0.n28_adj_1612\ : std_logic;
signal \c0.n26_adj_1613\ : std_logic;
signal \c0.n27_cascade_\ : std_logic;
signal \c0.n25_adj_1614\ : std_logic;
signal \c0.data_in_frame_20_0\ : std_logic;
signal \c0.n8995\ : std_logic;
signal \c0.n8834\ : std_logic;
signal \c0.n8924\ : std_logic;
signal \c0.n8852\ : std_logic;
signal \c0.n9013\ : std_logic;
signal data_in_field_70 : std_logic;
signal \c0.n12_cascade_\ : std_logic;
signal data_in_field_112 : std_logic;
signal \c0.data_in_frame_20_2\ : std_logic;
signal data_in_5_2 : std_logic;
signal data_in_4_2 : std_logic;
signal \r_SM_Main_2_adj_1738\ : std_logic;
signal \c0.tx2.n4880\ : std_logic;
signal \c0.n4525\ : std_logic;
signal \c0.n4244\ : std_logic;
signal data_in_field_50 : std_logic;
signal \c0.n20_adj_1642\ : std_logic;
signal \n12_adj_1753_cascade_\ : std_logic;
signal \r_SM_Main_2_N_1537_2_cascade_\ : std_logic;
signal \c0.rx.n4090\ : std_logic;
signal \c0.rx.n7393\ : std_logic;
signal data_in_field_122 : std_logic;
signal \c0.n4537\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_1543_0_cascade_\ : std_logic;
signal \n6_adj_1751_cascade_\ : std_logic;
signal \n30_cascade_\ : std_logic;
signal data_in_field_97 : std_logic;
signal data_in_field_95 : std_logic;
signal data_in_field_96 : std_logic;
signal \c0.n4296\ : std_logic;
signal \c0.rx.n12\ : std_logic;
signal tx_enable : std_logic;
signal n2185 : std_logic;
signal \r_Bit_Index_2_adj_1731\ : std_logic;
signal \n7415_cascade_\ : std_logic;
signal \n9301_cascade_\ : std_logic;
signal n1 : std_logic;
signal \r_Rx_Data\ : std_logic;
signal \c0.rx.r_SM_Main_2_N_1543_0\ : std_logic;
signal n9300 : std_logic;
signal \c0.data_in_field_24\ : std_logic;
signal \c0.data_in_field_16\ : std_logic;
signal \c0.data_in_field_8\ : std_logic;
signal \c0.data_in_field_0\ : std_logic;
signal \c0.n9446_cascade_\ : std_logic;
signal \c0.n9228\ : std_logic;
signal \c0.n9449_cascade_\ : std_logic;
signal data_in_field_80 : std_logic;
signal data_in_field_72 : std_logic;
signal \c0.n9740_cascade_\ : std_logic;
signal data_in_field_64 : std_logic;
signal \c0.n9234\ : std_logic;
signal \c0.n9231_cascade_\ : std_logic;
signal \c0.n9728\ : std_logic;
signal \c0.n22_adj_1661\ : std_logic;
signal \c0.n9731\ : std_logic;
signal \c0.tx2.r_Tx_Data_0\ : std_logic;
signal rx_data_ready : std_logic;
signal data_in_19_0 : std_logic;
signal data_in_18_0 : std_logic;
signal rand_data_12 : std_logic;
signal n4806 : std_logic;
signal data_in_field_88 : std_logic;
signal \c0.n4292\ : std_logic;
signal \c0.n8957\ : std_logic;
signal \c0.data_in_field_27\ : std_logic;
signal \c0.data_in_field_25\ : std_logic;
signal \c0.n8871\ : std_logic;
signal n26 : std_logic;
signal \bfn_11_27_0_\ : std_logic;
signal n25_adj_1722 : std_logic;
signal n8130 : std_logic;
signal n24 : std_logic;
signal n8131 : std_logic;
signal n23 : std_logic;
signal n8132 : std_logic;
signal n22 : std_logic;
signal n8133 : std_logic;
signal n21 : std_logic;
signal n8134 : std_logic;
signal n20 : std_logic;
signal n8135 : std_logic;
signal n19 : std_logic;
signal n8136 : std_logic;
signal n8137 : std_logic;
signal n18 : std_logic;
signal \bfn_11_28_0_\ : std_logic;
signal n17 : std_logic;
signal n8138 : std_logic;
signal n16 : std_logic;
signal n8139 : std_logic;
signal n15 : std_logic;
signal n8140 : std_logic;
signal n14 : std_logic;
signal n8141 : std_logic;
signal n13 : std_logic;
signal n8142 : std_logic;
signal n12 : std_logic;
signal n8143 : std_logic;
signal n11 : std_logic;
signal n8144 : std_logic;
signal n8145 : std_logic;
signal n10 : std_logic;
signal \bfn_11_29_0_\ : std_logic;
signal n9 : std_logic;
signal n8146 : std_logic;
signal n8 : std_logic;
signal n8147 : std_logic;
signal n7 : std_logic;
signal n8148 : std_logic;
signal n6 : std_logic;
signal n8149 : std_logic;
signal blink_counter_21 : std_logic;
signal n8150 : std_logic;
signal blink_counter_22 : std_logic;
signal n8151 : std_logic;
signal blink_counter_23 : std_logic;
signal n8152 : std_logic;
signal n8153 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_11_30_0_\ : std_logic;
signal n8154 : std_logic;
signal blink_counter_25 : std_logic;
signal \r_SM_Main_1_adj_1735\ : std_logic;
signal n9246 : std_logic;
signal \r_SM_Main_0_adj_1736\ : std_logic;
signal \n44_cascade_\ : std_logic;
signal \r_SM_Main_2_adj_1734\ : std_logic;
signal \r_SM_Main_2_N_1537_2\ : std_logic;
signal n9245 : std_logic;
signal \r_Clock_Count_0_adj_1730\ : std_logic;
signal n226 : std_logic;
signal \bfn_11_31_0_\ : std_logic;
signal \r_Clock_Count_1\ : std_logic;
signal n225 : std_logic;
signal \c0.rx.n8098\ : std_logic;
signal \r_Clock_Count_2\ : std_logic;
signal n224 : std_logic;
signal \c0.rx.n8099\ : std_logic;
signal \r_Clock_Count_3\ : std_logic;
signal n223 : std_logic;
signal \c0.rx.n8100\ : std_logic;
signal \c0.rx.n8101\ : std_logic;
signal \c0.rx.n8102\ : std_logic;
signal \r_Clock_Count_6_adj_1728\ : std_logic;
signal n220 : std_logic;
signal \c0.rx.n8103\ : std_logic;
signal \r_Clock_Count_7_adj_1727\ : std_logic;
signal \c0.rx.n8104\ : std_logic;
signal n219 : std_logic;
signal n4084 : std_logic;
signal n221 : std_logic;
signal \r_Clock_Count_5\ : std_logic;
signal n30 : std_logic;
signal n222 : std_logic;
signal n44 : std_logic;
signal \r_Clock_Count_4_adj_1729\ : std_logic;
signal \c0.n9192\ : std_logic;
signal \c0.n9195\ : std_logic;
signal \c0.n22_adj_1681\ : std_logic;
signal \c0.n9491_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2_4\ : std_logic;
signal \c0.tx2.r_Tx_Data_2\ : std_logic;
signal \c0.tx2.n3760\ : std_logic;
signal data_in_field_82 : std_logic;
signal data_in_field_90 : std_logic;
signal \c0.byte_transmit_counter2_0\ : std_logic;
signal data_in_field_66 : std_logic;
signal data_in_field_74 : std_logic;
signal \c0.n9500\ : std_logic;
signal \c0.byte_transmit_counter2_3\ : std_logic;
signal \c0.n9198_cascade_\ : std_logic;
signal \c0.n9488\ : std_logic;
signal data_in_field_98 : std_logic;
signal \c0.n9494\ : std_logic;
signal data_in_field_106 : std_logic;
signal \c0.n9201\ : std_logic;
signal \c0.n3056\ : std_logic;
signal \c0.n9671\ : std_logic;
signal \c0.data_in_frame_20_6\ : std_logic;
signal \c0.byte_transmit_counter2_2\ : std_logic;
signal \c0.n22_adj_1677\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \c0.n8083\ : std_logic;
signal \c0.n8084\ : std_logic;
signal \c0.n8085\ : std_logic;
signal \c0.n8086\ : std_logic;
signal \c0.n8087\ : std_logic;
signal \c0.n8088\ : std_logic;
signal \c0.n8089\ : std_logic;
signal \c0.n11_cascade_\ : std_logic;
signal \tx_data_3_N_keep_cascade_\ : std_logic;
signal \tx_data_0_N_keep\ : std_logic;
signal data_in_field_133 : std_logic;
signal data_in_field_103 : std_logic;
signal data_in_field_148 : std_logic;
signal \c0.n8986\ : std_logic;
signal \c0.n45_adj_1656\ : std_logic;
signal \tx_data_5_N_keep_cascade_\ : std_logic;
signal \c0.n11\ : std_logic;
signal \tx_data_2_N_keep_cascade_\ : std_logic;
signal \tx_data_6_N_keep\ : std_logic;
signal \n8705_cascade_\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal data_in_field_132 : std_logic;
signal \c0.n9680\ : std_logic;
signal data_in_field_140 : std_logic;
signal \c0.byte_transmit_counter2_1\ : std_logic;
signal \c0.n9683\ : std_logic;
signal \c0.n17_adj_1663_cascade_\ : std_logic;
signal \c0.n123_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.data_out_6_7_N_965_3\ : std_logic;
signal \c0.data_out_6_7_N_965_2\ : std_logic;
signal \c0.data_out_6_7_N_965_0\ : std_logic;
signal \c0.data_out_6_7_N_965_6\ : std_logic;
signal \c0.data_out_6_7_N_965_4\ : std_logic;
signal \c0.data_out_6_7_N_965_7\ : std_logic;
signal \c0.n7_cascade_\ : std_logic;
signal \c0.n8\ : std_logic;
signal \c0.n7814_cascade_\ : std_logic;
signal \data_out_6_7_N_965_5\ : std_logic;
signal \n7204_cascade_\ : std_logic;
signal byte_transmit_counter_5 : std_logic;
signal \c0.data_out_6_7_N_965_1\ : std_logic;
signal n7204 : std_logic;
signal \tx_data_1_N_keep_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n7779_cascade_\ : std_logic;
signal \tx_data_1_N_keep\ : std_logic;
signal \c0.data_out_6__7__N_973\ : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.byte_transmit_counter_4\ : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal \c0.byte_transmit_counter_3\ : std_logic;
signal \c0.n9291\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \tx_data_7_N_keep\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal n9710 : std_logic;
signal \n9713_cascade_\ : std_logic;
signal \n5_cascade_\ : std_logic;
signal \n3_cascade_\ : std_logic;
signal tx_o_adj_1726 : std_logic;
signal n9452 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal n9455 : std_logic;
signal \tx_data_4_N_keep\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal n9073 : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal n5062 : std_logic;
signal \n9073_cascade_\ : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal n3892 : std_logic;
signal \c0.n18_adj_1662\ : std_logic;
signal \c0.n19_adj_1664\ : std_logic;
signal \c0.n123\ : std_logic;
signal \c0.n7814\ : std_logic;
signal \c0.n117\ : std_logic;
signal n3747 : std_logic;
signal \c0.tx_active_prev\ : std_logic;
signal \n8749_cascade_\ : std_logic;
signal tx_active : std_logic;
signal \c0.tx.n8_cascade_\ : std_logic;
signal \c0.tx.n9059\ : std_logic;
signal n28 : std_logic;
signal \c0.tx_transmit\ : std_logic;
signal \n3151_cascade_\ : std_logic;
signal n11_adj_1752 : std_logic;
signal \c0.tx.n5_cascade_\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \c0.tx.n23_cascade_\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal n9259 : std_logic;
signal \c0.tx.n9027\ : std_logic;
signal \bfn_15_30_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \c0.tx.n9290\ : std_logic;
signal \c0.tx.n8090\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n9313\ : std_logic;
signal \c0.tx.n8091\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx.n9281\ : std_logic;
signal \c0.tx.n8092\ : std_logic;
signal \c0.tx.n8093\ : std_logic;
signal \c0.tx.n8094\ : std_logic;
signal \r_Clock_Count_6\ : std_logic;
signal n9304 : std_logic;
signal \c0.tx.n8095\ : std_logic;
signal \c0.tx.n8096\ : std_logic;
signal \c0.tx.n8097\ : std_logic;
signal \c0.tx.n7916\ : std_logic;
signal \bfn_15_31_0_\ : std_logic;
signal n9249 : std_logic;
signal \r_Clock_Count_0\ : std_logic;
signal n9266 : std_logic;
signal \c0.n900\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.delay_counter_0\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \c0.n21_adj_1653\ : std_logic;
signal \c0.delay_counter_1\ : std_logic;
signal \c0.n8120\ : std_logic;
signal \c0.n20_adj_1652\ : std_logic;
signal \c0.delay_counter_2\ : std_logic;
signal \c0.n8121\ : std_logic;
signal \c0.n19_adj_1651\ : std_logic;
signal \c0.delay_counter_3\ : std_logic;
signal \c0.n8122\ : std_logic;
signal \c0.n18_adj_1650\ : std_logic;
signal \c0.delay_counter_4\ : std_logic;
signal \c0.n8123\ : std_logic;
signal \c0.n17_adj_1649\ : std_logic;
signal \c0.delay_counter_5\ : std_logic;
signal \c0.n8124\ : std_logic;
signal \c0.n16_adj_1641\ : std_logic;
signal \c0.delay_counter_6\ : std_logic;
signal \c0.n8125\ : std_logic;
signal \c0.n15\ : std_logic;
signal \c0.delay_counter_7\ : std_logic;
signal \c0.n8126\ : std_logic;
signal \c0.n8127\ : std_logic;
signal \c0.n14_adj_1639\ : std_logic;
signal \c0.delay_counter_8\ : std_logic;
signal \bfn_16_26_0_\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.delay_counter_9\ : std_logic;
signal \c0.n8128\ : std_logic;
signal \c0.n12_adj_1634\ : std_logic;
signal \c0.n8129\ : std_logic;
signal \c0.delay_counter_10\ : std_logic;
signal \UART_TRANSMITTER_state_0\ : std_logic;
signal \r_SM_Main_2_N_1480_1\ : std_logic;
signal \c0.tx.n23\ : std_logic;
signal \r_Clock_Count_8\ : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \c0.tx.n9310\ : std_logic;
signal n9305 : std_logic;
signal \r_Clock_Count_4\ : std_logic;
signal \c0.tx.n9314\ : std_logic;
signal \c0.tx.r_Clock_Count_5\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal n9303 : std_logic;
signal \r_Clock_Count_7\ : std_logic;
signal \CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35917\,
            DIN => \N__35916\,
            DOUT => \N__35915\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35917\,
            PADOUT => \N__35916\,
            PADIN => \N__35915\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19242\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35908\,
            DIN => \N__35907\,
            DOUT => \N__35906\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35908\,
            PADOUT => \N__35907\,
            PADIN => \N__35906\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__35899\,
            DIN => \N__35898\,
            DOUT => \N__35897\,
            PACKAGEPIN => PIN_2
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35899\,
            PADOUT => \N__35898\,
            PADIN => \N__35897\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \c0.rx.r_Rx_Data_R\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__35382\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx2_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__35890\,
            DIN => \N__35889\,
            DOUT => \N__35888\,
            PACKAGEPIN => PIN_3
        );

    \tx2_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35890\,
            PADOUT => \N__35889\,
            PADIN => \N__35888\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15786\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__13179\
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__35881\,
            DIN => \N__35880\,
            DOUT => \N__35879\,
            PACKAGEPIN => PIN_1
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35881\,
            PADOUT => \N__35880\,
            PADIN => \N__35879\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__34119\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__27585\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35872\,
            DIN => \N__35871\,
            DOUT => \N__35870\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35872\,
            PADOUT => \N__35871\,
            PADIN => \N__35870\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__8861\ : InMux
    port map (
            O => \N__35853\,
            I => \c0.n8129\
        );

    \I__8860\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35847\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35843\
        );

    \I__8858\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35840\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__35843\,
            I => \N__35837\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__35840\,
            I => \c0.delay_counter_10\
        );

    \I__8855\ : Odrv4
    port map (
            O => \N__35837\,
            I => \c0.delay_counter_10\
        );

    \I__8854\ : CEMux
    port map (
            O => \N__35832\,
            I => \N__35828\
        );

    \I__8853\ : CEMux
    port map (
            O => \N__35831\,
            I => \N__35824\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__35828\,
            I => \N__35821\
        );

    \I__8851\ : CascadeMux
    port map (
            O => \N__35827\,
            I => \N__35818\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__35824\,
            I => \N__35809\
        );

    \I__8849\ : Span4Mux_h
    port map (
            O => \N__35821\,
            I => \N__35806\
        );

    \I__8848\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35799\
        );

    \I__8847\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35799\
        );

    \I__8846\ : InMux
    port map (
            O => \N__35816\,
            I => \N__35799\
        );

    \I__8845\ : CascadeMux
    port map (
            O => \N__35815\,
            I => \N__35796\
        );

    \I__8844\ : CascadeMux
    port map (
            O => \N__35814\,
            I => \N__35793\
        );

    \I__8843\ : CascadeMux
    port map (
            O => \N__35813\,
            I => \N__35790\
        );

    \I__8842\ : CascadeMux
    port map (
            O => \N__35812\,
            I => \N__35787\
        );

    \I__8841\ : Span4Mux_h
    port map (
            O => \N__35809\,
            I => \N__35781\
        );

    \I__8840\ : Sp12to4
    port map (
            O => \N__35806\,
            I => \N__35778\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__35799\,
            I => \N__35775\
        );

    \I__8838\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35772\
        );

    \I__8837\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35769\
        );

    \I__8836\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35758\
        );

    \I__8835\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35758\
        );

    \I__8834\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35758\
        );

    \I__8833\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35758\
        );

    \I__8832\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35758\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__35781\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__8830\ : Odrv12
    port map (
            O => \N__35778\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__8829\ : Odrv4
    port map (
            O => \N__35775\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__35772\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__35769\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__35758\,
            I => \UART_TRANSMITTER_state_0\
        );

    \I__8825\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35741\
        );

    \I__8824\ : CascadeMux
    port map (
            O => \N__35744\,
            I => \N__35738\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__35741\,
            I => \N__35732\
        );

    \I__8822\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35725\
        );

    \I__8821\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35725\
        );

    \I__8820\ : InMux
    port map (
            O => \N__35736\,
            I => \N__35725\
        );

    \I__8819\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35722\
        );

    \I__8818\ : Span4Mux_v
    port map (
            O => \N__35732\,
            I => \N__35719\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__35725\,
            I => \r_SM_Main_2_N_1480_1\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__35722\,
            I => \r_SM_Main_2_N_1480_1\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__35719\,
            I => \r_SM_Main_2_N_1480_1\
        );

    \I__8814\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35704\
        );

    \I__8813\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35704\
        );

    \I__8812\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35699\
        );

    \I__8811\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35699\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__35704\,
            I => \c0.tx.n23\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__35699\,
            I => \c0.tx.n23\
        );

    \I__8808\ : CascadeMux
    port map (
            O => \N__35694\,
            I => \N__35691\
        );

    \I__8807\ : InMux
    port map (
            O => \N__35691\,
            I => \N__35684\
        );

    \I__8806\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35684\
        );

    \I__8805\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35678\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35675\
        );

    \I__8803\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35672\
        );

    \I__8802\ : InMux
    port map (
            O => \N__35682\,
            I => \N__35669\
        );

    \I__8801\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35666\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__35678\,
            I => \N__35661\
        );

    \I__8799\ : Span4Mux_h
    port map (
            O => \N__35675\,
            I => \N__35661\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__35672\,
            I => \N__35658\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__35669\,
            I => \r_Clock_Count_8\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__35666\,
            I => \r_Clock_Count_8\
        );

    \I__8795\ : Odrv4
    port map (
            O => \N__35661\,
            I => \r_Clock_Count_8\
        );

    \I__8794\ : Odrv12
    port map (
            O => \N__35658\,
            I => \r_Clock_Count_8\
        );

    \I__8793\ : InMux
    port map (
            O => \N__35649\,
            I => \N__35646\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__35646\,
            I => \N__35642\
        );

    \I__8791\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35639\
        );

    \I__8790\ : Span4Mux_v
    port map (
            O => \N__35642\,
            I => \N__35633\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__35639\,
            I => \N__35633\
        );

    \I__8788\ : InMux
    port map (
            O => \N__35638\,
            I => \N__35627\
        );

    \I__8787\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35624\
        );

    \I__8786\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35617\
        );

    \I__8785\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35617\
        );

    \I__8784\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35617\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__35627\,
            I => \r_Bit_Index_2\
        );

    \I__8782\ : Odrv4
    port map (
            O => \N__35624\,
            I => \r_Bit_Index_2\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__35617\,
            I => \r_Bit_Index_2\
        );

    \I__8780\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35607\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__35607\,
            I => \c0.tx.n9310\
        );

    \I__8778\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35601\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__35601\,
            I => n9305
        );

    \I__8776\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35593\
        );

    \I__8775\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35590\
        );

    \I__8774\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35587\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__35593\,
            I => \r_Clock_Count_4\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__35590\,
            I => \r_Clock_Count_4\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__35587\,
            I => \r_Clock_Count_4\
        );

    \I__8770\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35577\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__35577\,
            I => \c0.tx.n9314\
        );

    \I__8768\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35569\
        );

    \I__8767\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35566\
        );

    \I__8766\ : InMux
    port map (
            O => \N__35572\,
            I => \N__35563\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__35569\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__35566\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__35563\,
            I => \c0.tx.r_Clock_Count_5\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__35556\,
            I => \N__35547\
        );

    \I__8761\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35540\
        );

    \I__8760\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35540\
        );

    \I__8759\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35531\
        );

    \I__8758\ : InMux
    port map (
            O => \N__35552\,
            I => \N__35526\
        );

    \I__8757\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35526\
        );

    \I__8756\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35517\
        );

    \I__8755\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35517\
        );

    \I__8754\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35517\
        );

    \I__8753\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35517\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__35540\,
            I => \N__35509\
        );

    \I__8751\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35506\
        );

    \I__8750\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35503\
        );

    \I__8749\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35498\
        );

    \I__8748\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35498\
        );

    \I__8747\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35493\
        );

    \I__8746\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35493\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35486\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__35526\,
            I => \N__35486\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__35517\,
            I => \N__35486\
        );

    \I__8742\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35475\
        );

    \I__8741\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35475\
        );

    \I__8740\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35475\
        );

    \I__8739\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35475\
        );

    \I__8738\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35475\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__35509\,
            I => \r_SM_Main_2\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__35506\,
            I => \r_SM_Main_2\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__35503\,
            I => \r_SM_Main_2\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__35498\,
            I => \r_SM_Main_2\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__35493\,
            I => \r_SM_Main_2\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__35486\,
            I => \r_SM_Main_2\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__35475\,
            I => \r_SM_Main_2\
        );

    \I__8730\ : InMux
    port map (
            O => \N__35460\,
            I => \N__35457\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__35457\,
            I => n9303
        );

    \I__8728\ : InMux
    port map (
            O => \N__35454\,
            I => \N__35449\
        );

    \I__8727\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35446\
        );

    \I__8726\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35443\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__35449\,
            I => \r_Clock_Count_7\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__35446\,
            I => \r_Clock_Count_7\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__35443\,
            I => \r_Clock_Count_7\
        );

    \I__8722\ : ClkMux
    port map (
            O => \N__35436\,
            I => \N__34995\
        );

    \I__8721\ : ClkMux
    port map (
            O => \N__35435\,
            I => \N__34995\
        );

    \I__8720\ : ClkMux
    port map (
            O => \N__35434\,
            I => \N__34995\
        );

    \I__8719\ : ClkMux
    port map (
            O => \N__35433\,
            I => \N__34995\
        );

    \I__8718\ : ClkMux
    port map (
            O => \N__35432\,
            I => \N__34995\
        );

    \I__8717\ : ClkMux
    port map (
            O => \N__35431\,
            I => \N__34995\
        );

    \I__8716\ : ClkMux
    port map (
            O => \N__35430\,
            I => \N__34995\
        );

    \I__8715\ : ClkMux
    port map (
            O => \N__35429\,
            I => \N__34995\
        );

    \I__8714\ : ClkMux
    port map (
            O => \N__35428\,
            I => \N__34995\
        );

    \I__8713\ : ClkMux
    port map (
            O => \N__35427\,
            I => \N__34995\
        );

    \I__8712\ : ClkMux
    port map (
            O => \N__35426\,
            I => \N__34995\
        );

    \I__8711\ : ClkMux
    port map (
            O => \N__35425\,
            I => \N__34995\
        );

    \I__8710\ : ClkMux
    port map (
            O => \N__35424\,
            I => \N__34995\
        );

    \I__8709\ : ClkMux
    port map (
            O => \N__35423\,
            I => \N__34995\
        );

    \I__8708\ : ClkMux
    port map (
            O => \N__35422\,
            I => \N__34995\
        );

    \I__8707\ : ClkMux
    port map (
            O => \N__35421\,
            I => \N__34995\
        );

    \I__8706\ : ClkMux
    port map (
            O => \N__35420\,
            I => \N__34995\
        );

    \I__8705\ : ClkMux
    port map (
            O => \N__35419\,
            I => \N__34995\
        );

    \I__8704\ : ClkMux
    port map (
            O => \N__35418\,
            I => \N__34995\
        );

    \I__8703\ : ClkMux
    port map (
            O => \N__35417\,
            I => \N__34995\
        );

    \I__8702\ : ClkMux
    port map (
            O => \N__35416\,
            I => \N__34995\
        );

    \I__8701\ : ClkMux
    port map (
            O => \N__35415\,
            I => \N__34995\
        );

    \I__8700\ : ClkMux
    port map (
            O => \N__35414\,
            I => \N__34995\
        );

    \I__8699\ : ClkMux
    port map (
            O => \N__35413\,
            I => \N__34995\
        );

    \I__8698\ : ClkMux
    port map (
            O => \N__35412\,
            I => \N__34995\
        );

    \I__8697\ : ClkMux
    port map (
            O => \N__35411\,
            I => \N__34995\
        );

    \I__8696\ : ClkMux
    port map (
            O => \N__35410\,
            I => \N__34995\
        );

    \I__8695\ : ClkMux
    port map (
            O => \N__35409\,
            I => \N__34995\
        );

    \I__8694\ : ClkMux
    port map (
            O => \N__35408\,
            I => \N__34995\
        );

    \I__8693\ : ClkMux
    port map (
            O => \N__35407\,
            I => \N__34995\
        );

    \I__8692\ : ClkMux
    port map (
            O => \N__35406\,
            I => \N__34995\
        );

    \I__8691\ : ClkMux
    port map (
            O => \N__35405\,
            I => \N__34995\
        );

    \I__8690\ : ClkMux
    port map (
            O => \N__35404\,
            I => \N__34995\
        );

    \I__8689\ : ClkMux
    port map (
            O => \N__35403\,
            I => \N__34995\
        );

    \I__8688\ : ClkMux
    port map (
            O => \N__35402\,
            I => \N__34995\
        );

    \I__8687\ : ClkMux
    port map (
            O => \N__35401\,
            I => \N__34995\
        );

    \I__8686\ : ClkMux
    port map (
            O => \N__35400\,
            I => \N__34995\
        );

    \I__8685\ : ClkMux
    port map (
            O => \N__35399\,
            I => \N__34995\
        );

    \I__8684\ : ClkMux
    port map (
            O => \N__35398\,
            I => \N__34995\
        );

    \I__8683\ : ClkMux
    port map (
            O => \N__35397\,
            I => \N__34995\
        );

    \I__8682\ : ClkMux
    port map (
            O => \N__35396\,
            I => \N__34995\
        );

    \I__8681\ : ClkMux
    port map (
            O => \N__35395\,
            I => \N__34995\
        );

    \I__8680\ : ClkMux
    port map (
            O => \N__35394\,
            I => \N__34995\
        );

    \I__8679\ : ClkMux
    port map (
            O => \N__35393\,
            I => \N__34995\
        );

    \I__8678\ : ClkMux
    port map (
            O => \N__35392\,
            I => \N__34995\
        );

    \I__8677\ : ClkMux
    port map (
            O => \N__35391\,
            I => \N__34995\
        );

    \I__8676\ : ClkMux
    port map (
            O => \N__35390\,
            I => \N__34995\
        );

    \I__8675\ : ClkMux
    port map (
            O => \N__35389\,
            I => \N__34995\
        );

    \I__8674\ : ClkMux
    port map (
            O => \N__35388\,
            I => \N__34995\
        );

    \I__8673\ : ClkMux
    port map (
            O => \N__35387\,
            I => \N__34995\
        );

    \I__8672\ : ClkMux
    port map (
            O => \N__35386\,
            I => \N__34995\
        );

    \I__8671\ : ClkMux
    port map (
            O => \N__35385\,
            I => \N__34995\
        );

    \I__8670\ : ClkMux
    port map (
            O => \N__35384\,
            I => \N__34995\
        );

    \I__8669\ : ClkMux
    port map (
            O => \N__35383\,
            I => \N__34995\
        );

    \I__8668\ : ClkMux
    port map (
            O => \N__35382\,
            I => \N__34995\
        );

    \I__8667\ : ClkMux
    port map (
            O => \N__35381\,
            I => \N__34995\
        );

    \I__8666\ : ClkMux
    port map (
            O => \N__35380\,
            I => \N__34995\
        );

    \I__8665\ : ClkMux
    port map (
            O => \N__35379\,
            I => \N__34995\
        );

    \I__8664\ : ClkMux
    port map (
            O => \N__35378\,
            I => \N__34995\
        );

    \I__8663\ : ClkMux
    port map (
            O => \N__35377\,
            I => \N__34995\
        );

    \I__8662\ : ClkMux
    port map (
            O => \N__35376\,
            I => \N__34995\
        );

    \I__8661\ : ClkMux
    port map (
            O => \N__35375\,
            I => \N__34995\
        );

    \I__8660\ : ClkMux
    port map (
            O => \N__35374\,
            I => \N__34995\
        );

    \I__8659\ : ClkMux
    port map (
            O => \N__35373\,
            I => \N__34995\
        );

    \I__8658\ : ClkMux
    port map (
            O => \N__35372\,
            I => \N__34995\
        );

    \I__8657\ : ClkMux
    port map (
            O => \N__35371\,
            I => \N__34995\
        );

    \I__8656\ : ClkMux
    port map (
            O => \N__35370\,
            I => \N__34995\
        );

    \I__8655\ : ClkMux
    port map (
            O => \N__35369\,
            I => \N__34995\
        );

    \I__8654\ : ClkMux
    port map (
            O => \N__35368\,
            I => \N__34995\
        );

    \I__8653\ : ClkMux
    port map (
            O => \N__35367\,
            I => \N__34995\
        );

    \I__8652\ : ClkMux
    port map (
            O => \N__35366\,
            I => \N__34995\
        );

    \I__8651\ : ClkMux
    port map (
            O => \N__35365\,
            I => \N__34995\
        );

    \I__8650\ : ClkMux
    port map (
            O => \N__35364\,
            I => \N__34995\
        );

    \I__8649\ : ClkMux
    port map (
            O => \N__35363\,
            I => \N__34995\
        );

    \I__8648\ : ClkMux
    port map (
            O => \N__35362\,
            I => \N__34995\
        );

    \I__8647\ : ClkMux
    port map (
            O => \N__35361\,
            I => \N__34995\
        );

    \I__8646\ : ClkMux
    port map (
            O => \N__35360\,
            I => \N__34995\
        );

    \I__8645\ : ClkMux
    port map (
            O => \N__35359\,
            I => \N__34995\
        );

    \I__8644\ : ClkMux
    port map (
            O => \N__35358\,
            I => \N__34995\
        );

    \I__8643\ : ClkMux
    port map (
            O => \N__35357\,
            I => \N__34995\
        );

    \I__8642\ : ClkMux
    port map (
            O => \N__35356\,
            I => \N__34995\
        );

    \I__8641\ : ClkMux
    port map (
            O => \N__35355\,
            I => \N__34995\
        );

    \I__8640\ : ClkMux
    port map (
            O => \N__35354\,
            I => \N__34995\
        );

    \I__8639\ : ClkMux
    port map (
            O => \N__35353\,
            I => \N__34995\
        );

    \I__8638\ : ClkMux
    port map (
            O => \N__35352\,
            I => \N__34995\
        );

    \I__8637\ : ClkMux
    port map (
            O => \N__35351\,
            I => \N__34995\
        );

    \I__8636\ : ClkMux
    port map (
            O => \N__35350\,
            I => \N__34995\
        );

    \I__8635\ : ClkMux
    port map (
            O => \N__35349\,
            I => \N__34995\
        );

    \I__8634\ : ClkMux
    port map (
            O => \N__35348\,
            I => \N__34995\
        );

    \I__8633\ : ClkMux
    port map (
            O => \N__35347\,
            I => \N__34995\
        );

    \I__8632\ : ClkMux
    port map (
            O => \N__35346\,
            I => \N__34995\
        );

    \I__8631\ : ClkMux
    port map (
            O => \N__35345\,
            I => \N__34995\
        );

    \I__8630\ : ClkMux
    port map (
            O => \N__35344\,
            I => \N__34995\
        );

    \I__8629\ : ClkMux
    port map (
            O => \N__35343\,
            I => \N__34995\
        );

    \I__8628\ : ClkMux
    port map (
            O => \N__35342\,
            I => \N__34995\
        );

    \I__8627\ : ClkMux
    port map (
            O => \N__35341\,
            I => \N__34995\
        );

    \I__8626\ : ClkMux
    port map (
            O => \N__35340\,
            I => \N__34995\
        );

    \I__8625\ : ClkMux
    port map (
            O => \N__35339\,
            I => \N__34995\
        );

    \I__8624\ : ClkMux
    port map (
            O => \N__35338\,
            I => \N__34995\
        );

    \I__8623\ : ClkMux
    port map (
            O => \N__35337\,
            I => \N__34995\
        );

    \I__8622\ : ClkMux
    port map (
            O => \N__35336\,
            I => \N__34995\
        );

    \I__8621\ : ClkMux
    port map (
            O => \N__35335\,
            I => \N__34995\
        );

    \I__8620\ : ClkMux
    port map (
            O => \N__35334\,
            I => \N__34995\
        );

    \I__8619\ : ClkMux
    port map (
            O => \N__35333\,
            I => \N__34995\
        );

    \I__8618\ : ClkMux
    port map (
            O => \N__35332\,
            I => \N__34995\
        );

    \I__8617\ : ClkMux
    port map (
            O => \N__35331\,
            I => \N__34995\
        );

    \I__8616\ : ClkMux
    port map (
            O => \N__35330\,
            I => \N__34995\
        );

    \I__8615\ : ClkMux
    port map (
            O => \N__35329\,
            I => \N__34995\
        );

    \I__8614\ : ClkMux
    port map (
            O => \N__35328\,
            I => \N__34995\
        );

    \I__8613\ : ClkMux
    port map (
            O => \N__35327\,
            I => \N__34995\
        );

    \I__8612\ : ClkMux
    port map (
            O => \N__35326\,
            I => \N__34995\
        );

    \I__8611\ : ClkMux
    port map (
            O => \N__35325\,
            I => \N__34995\
        );

    \I__8610\ : ClkMux
    port map (
            O => \N__35324\,
            I => \N__34995\
        );

    \I__8609\ : ClkMux
    port map (
            O => \N__35323\,
            I => \N__34995\
        );

    \I__8608\ : ClkMux
    port map (
            O => \N__35322\,
            I => \N__34995\
        );

    \I__8607\ : ClkMux
    port map (
            O => \N__35321\,
            I => \N__34995\
        );

    \I__8606\ : ClkMux
    port map (
            O => \N__35320\,
            I => \N__34995\
        );

    \I__8605\ : ClkMux
    port map (
            O => \N__35319\,
            I => \N__34995\
        );

    \I__8604\ : ClkMux
    port map (
            O => \N__35318\,
            I => \N__34995\
        );

    \I__8603\ : ClkMux
    port map (
            O => \N__35317\,
            I => \N__34995\
        );

    \I__8602\ : ClkMux
    port map (
            O => \N__35316\,
            I => \N__34995\
        );

    \I__8601\ : ClkMux
    port map (
            O => \N__35315\,
            I => \N__34995\
        );

    \I__8600\ : ClkMux
    port map (
            O => \N__35314\,
            I => \N__34995\
        );

    \I__8599\ : ClkMux
    port map (
            O => \N__35313\,
            I => \N__34995\
        );

    \I__8598\ : ClkMux
    port map (
            O => \N__35312\,
            I => \N__34995\
        );

    \I__8597\ : ClkMux
    port map (
            O => \N__35311\,
            I => \N__34995\
        );

    \I__8596\ : ClkMux
    port map (
            O => \N__35310\,
            I => \N__34995\
        );

    \I__8595\ : ClkMux
    port map (
            O => \N__35309\,
            I => \N__34995\
        );

    \I__8594\ : ClkMux
    port map (
            O => \N__35308\,
            I => \N__34995\
        );

    \I__8593\ : ClkMux
    port map (
            O => \N__35307\,
            I => \N__34995\
        );

    \I__8592\ : ClkMux
    port map (
            O => \N__35306\,
            I => \N__34995\
        );

    \I__8591\ : ClkMux
    port map (
            O => \N__35305\,
            I => \N__34995\
        );

    \I__8590\ : ClkMux
    port map (
            O => \N__35304\,
            I => \N__34995\
        );

    \I__8589\ : ClkMux
    port map (
            O => \N__35303\,
            I => \N__34995\
        );

    \I__8588\ : ClkMux
    port map (
            O => \N__35302\,
            I => \N__34995\
        );

    \I__8587\ : ClkMux
    port map (
            O => \N__35301\,
            I => \N__34995\
        );

    \I__8586\ : ClkMux
    port map (
            O => \N__35300\,
            I => \N__34995\
        );

    \I__8585\ : ClkMux
    port map (
            O => \N__35299\,
            I => \N__34995\
        );

    \I__8584\ : ClkMux
    port map (
            O => \N__35298\,
            I => \N__34995\
        );

    \I__8583\ : ClkMux
    port map (
            O => \N__35297\,
            I => \N__34995\
        );

    \I__8582\ : ClkMux
    port map (
            O => \N__35296\,
            I => \N__34995\
        );

    \I__8581\ : ClkMux
    port map (
            O => \N__35295\,
            I => \N__34995\
        );

    \I__8580\ : ClkMux
    port map (
            O => \N__35294\,
            I => \N__34995\
        );

    \I__8579\ : ClkMux
    port map (
            O => \N__35293\,
            I => \N__34995\
        );

    \I__8578\ : ClkMux
    port map (
            O => \N__35292\,
            I => \N__34995\
        );

    \I__8577\ : ClkMux
    port map (
            O => \N__35291\,
            I => \N__34995\
        );

    \I__8576\ : ClkMux
    port map (
            O => \N__35290\,
            I => \N__34995\
        );

    \I__8575\ : GlobalMux
    port map (
            O => \N__34995\,
            I => \N__34992\
        );

    \I__8574\ : gio2CtrlBuf
    port map (
            O => \N__34992\,
            I => \CLK_c\
        );

    \I__8573\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__34986\,
            I => \c0.n19_adj_1651\
        );

    \I__8571\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34979\
        );

    \I__8570\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34976\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__34979\,
            I => \N__34973\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__34976\,
            I => \c0.delay_counter_3\
        );

    \I__8567\ : Odrv12
    port map (
            O => \N__34973\,
            I => \c0.delay_counter_3\
        );

    \I__8566\ : InMux
    port map (
            O => \N__34968\,
            I => \c0.n8122\
        );

    \I__8565\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34962\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__34962\,
            I => \c0.n18_adj_1650\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__34959\,
            I => \N__34955\
        );

    \I__8562\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34950\
        );

    \I__8561\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34950\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__34950\,
            I => \c0.delay_counter_4\
        );

    \I__8559\ : InMux
    port map (
            O => \N__34947\,
            I => \c0.n8123\
        );

    \I__8558\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34941\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__34941\,
            I => \c0.n17_adj_1649\
        );

    \I__8556\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34934\
        );

    \I__8555\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34931\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__34934\,
            I => \c0.delay_counter_5\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__34931\,
            I => \c0.delay_counter_5\
        );

    \I__8552\ : InMux
    port map (
            O => \N__34926\,
            I => \c0.n8124\
        );

    \I__8551\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__34920\,
            I => \c0.n16_adj_1641\
        );

    \I__8549\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34913\
        );

    \I__8548\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34910\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34907\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__34910\,
            I => \c0.delay_counter_6\
        );

    \I__8545\ : Odrv12
    port map (
            O => \N__34907\,
            I => \c0.delay_counter_6\
        );

    \I__8544\ : InMux
    port map (
            O => \N__34902\,
            I => \c0.n8125\
        );

    \I__8543\ : InMux
    port map (
            O => \N__34899\,
            I => \N__34896\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__34896\,
            I => \c0.n15\
        );

    \I__8541\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34887\
        );

    \I__8540\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34887\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__34887\,
            I => \c0.delay_counter_7\
        );

    \I__8538\ : InMux
    port map (
            O => \N__34884\,
            I => \c0.n8126\
        );

    \I__8537\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__34878\,
            I => \c0.n14_adj_1639\
        );

    \I__8535\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34871\
        );

    \I__8534\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34868\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__34871\,
            I => \c0.delay_counter_8\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__34868\,
            I => \c0.delay_counter_8\
        );

    \I__8531\ : InMux
    port map (
            O => \N__34863\,
            I => \bfn_16_26_0_\
        );

    \I__8530\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__34857\,
            I => \c0.n13\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__34854\,
            I => \N__34850\
        );

    \I__8527\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34847\
        );

    \I__8526\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34844\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__34847\,
            I => \c0.delay_counter_9\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__34844\,
            I => \c0.delay_counter_9\
        );

    \I__8523\ : InMux
    port map (
            O => \N__34839\,
            I => \c0.n8128\
        );

    \I__8522\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34833\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__34833\,
            I => \c0.n12_adj_1634\
        );

    \I__8520\ : InMux
    port map (
            O => \N__34830\,
            I => \c0.tx.n8094\
        );

    \I__8519\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34822\
        );

    \I__8518\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34817\
        );

    \I__8517\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34817\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__34822\,
            I => \r_Clock_Count_6\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__34817\,
            I => \r_Clock_Count_6\
        );

    \I__8514\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34809\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__34809\,
            I => n9304
        );

    \I__8512\ : InMux
    port map (
            O => \N__34806\,
            I => \c0.tx.n8095\
        );

    \I__8511\ : InMux
    port map (
            O => \N__34803\,
            I => \c0.tx.n8096\
        );

    \I__8510\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34789\
        );

    \I__8509\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34780\
        );

    \I__8508\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34780\
        );

    \I__8507\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34780\
        );

    \I__8506\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34780\
        );

    \I__8505\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34771\
        );

    \I__8504\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34771\
        );

    \I__8503\ : InMux
    port map (
            O => \N__34793\,
            I => \N__34771\
        );

    \I__8502\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34771\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__34789\,
            I => \N__34768\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__34780\,
            I => \c0.tx.n7916\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__34771\,
            I => \c0.tx.n7916\
        );

    \I__8498\ : Odrv4
    port map (
            O => \N__34768\,
            I => \c0.tx.n7916\
        );

    \I__8497\ : InMux
    port map (
            O => \N__34761\,
            I => \bfn_15_31_0_\
        );

    \I__8496\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34755\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__34755\,
            I => n9249
        );

    \I__8494\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34748\
        );

    \I__8493\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34745\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__34748\,
            I => \r_Clock_Count_0\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__34745\,
            I => \r_Clock_Count_0\
        );

    \I__8490\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34737\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__34737\,
            I => n9266
        );

    \I__8488\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__34731\,
            I => \c0.n900\
        );

    \I__8486\ : CascadeMux
    port map (
            O => \N__34728\,
            I => \N__34725\
        );

    \I__8485\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34722\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__34722\,
            I => \c0.n22\
        );

    \I__8483\ : InMux
    port map (
            O => \N__34719\,
            I => \N__34715\
        );

    \I__8482\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34712\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__34715\,
            I => \N__34709\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__34712\,
            I => \c0.delay_counter_0\
        );

    \I__8479\ : Odrv4
    port map (
            O => \N__34709\,
            I => \c0.delay_counter_0\
        );

    \I__8478\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34701\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__34701\,
            I => \c0.n21_adj_1653\
        );

    \I__8476\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34692\
        );

    \I__8475\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34692\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__34692\,
            I => \c0.delay_counter_1\
        );

    \I__8473\ : InMux
    port map (
            O => \N__34689\,
            I => \c0.n8120\
        );

    \I__8472\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34683\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__34683\,
            I => \c0.n20_adj_1652\
        );

    \I__8470\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34674\
        );

    \I__8469\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34674\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__34674\,
            I => \c0.delay_counter_2\
        );

    \I__8467\ : InMux
    port map (
            O => \N__34671\,
            I => \c0.n8121\
        );

    \I__8466\ : InMux
    port map (
            O => \N__34668\,
            I => \N__34665\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__34665\,
            I => \c0.tx.n9027\
        );

    \I__8464\ : InMux
    port map (
            O => \N__34662\,
            I => \bfn_15_30_0_\
        );

    \I__8463\ : CascadeMux
    port map (
            O => \N__34659\,
            I => \N__34654\
        );

    \I__8462\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34651\
        );

    \I__8461\ : InMux
    port map (
            O => \N__34657\,
            I => \N__34648\
        );

    \I__8460\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34645\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__34651\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__34648\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__34645\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__8456\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34635\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__34635\,
            I => \c0.tx.n9290\
        );

    \I__8454\ : InMux
    port map (
            O => \N__34632\,
            I => \c0.tx.n8090\
        );

    \I__8453\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34624\
        );

    \I__8452\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34619\
        );

    \I__8451\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34619\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__34624\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__34619\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__8448\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34611\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__34611\,
            I => \c0.tx.n9313\
        );

    \I__8446\ : InMux
    port map (
            O => \N__34608\,
            I => \c0.tx.n8091\
        );

    \I__8445\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34600\
        );

    \I__8444\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34595\
        );

    \I__8443\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34595\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__34600\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__34595\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__8440\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34587\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__34587\,
            I => \c0.tx.n9281\
        );

    \I__8438\ : InMux
    port map (
            O => \N__34584\,
            I => \c0.tx.n8092\
        );

    \I__8437\ : InMux
    port map (
            O => \N__34581\,
            I => \c0.tx.n8093\
        );

    \I__8436\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__34575\,
            I => \c0.tx.n9059\
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__34572\,
            I => \N__34569\
        );

    \I__8433\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34565\
        );

    \I__8432\ : CascadeMux
    port map (
            O => \N__34568\,
            I => \N__34562\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34559\
        );

    \I__8430\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34556\
        );

    \I__8429\ : Span4Mux_h
    port map (
            O => \N__34559\,
            I => \N__34551\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__34556\,
            I => \N__34551\
        );

    \I__8427\ : Odrv4
    port map (
            O => \N__34551\,
            I => n28
        );

    \I__8426\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34544\
        );

    \I__8425\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34537\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34534\
        );

    \I__8423\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34531\
        );

    \I__8422\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34524\
        );

    \I__8421\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34524\
        );

    \I__8420\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34524\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__34537\,
            I => \c0.tx_transmit\
        );

    \I__8418\ : Odrv4
    port map (
            O => \N__34534\,
            I => \c0.tx_transmit\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__34531\,
            I => \c0.tx_transmit\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__34524\,
            I => \c0.tx_transmit\
        );

    \I__8415\ : CascadeMux
    port map (
            O => \N__34515\,
            I => \n3151_cascade_\
        );

    \I__8414\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34509\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__34509\,
            I => n11_adj_1752
        );

    \I__8412\ : CascadeMux
    port map (
            O => \N__34506\,
            I => \c0.tx.n5_cascade_\
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__34503\,
            I => \N__34496\
        );

    \I__8410\ : CascadeMux
    port map (
            O => \N__34502\,
            I => \N__34493\
        );

    \I__8409\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34490\
        );

    \I__8408\ : CascadeMux
    port map (
            O => \N__34500\,
            I => \N__34487\
        );

    \I__8407\ : CascadeMux
    port map (
            O => \N__34499\,
            I => \N__34480\
        );

    \I__8406\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34474\
        );

    \I__8405\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34474\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__34490\,
            I => \N__34471\
        );

    \I__8403\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34468\
        );

    \I__8402\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34463\
        );

    \I__8401\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34463\
        );

    \I__8400\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34454\
        );

    \I__8399\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34454\
        );

    \I__8398\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34454\
        );

    \I__8397\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34454\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__34474\,
            I => \r_SM_Main_0\
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__34471\,
            I => \r_SM_Main_0\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__34468\,
            I => \r_SM_Main_0\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__34463\,
            I => \r_SM_Main_0\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__34454\,
            I => \r_SM_Main_0\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__34443\,
            I => \c0.tx.n23_cascade_\
        );

    \I__8390\ : CascadeMux
    port map (
            O => \N__34440\,
            I => \N__34436\
        );

    \I__8389\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34433\
        );

    \I__8388\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34430\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34414\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__34430\,
            I => \N__34414\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__34429\,
            I => \N__34411\
        );

    \I__8384\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34407\
        );

    \I__8383\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34404\
        );

    \I__8382\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34397\
        );

    \I__8381\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34397\
        );

    \I__8380\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34397\
        );

    \I__8379\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34394\
        );

    \I__8378\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34389\
        );

    \I__8377\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34389\
        );

    \I__8376\ : InMux
    port map (
            O => \N__34420\,
            I => \N__34384\
        );

    \I__8375\ : InMux
    port map (
            O => \N__34419\,
            I => \N__34384\
        );

    \I__8374\ : Span4Mux_h
    port map (
            O => \N__34414\,
            I => \N__34381\
        );

    \I__8373\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34376\
        );

    \I__8372\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34376\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__34407\,
            I => \r_SM_Main_1\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__34404\,
            I => \r_SM_Main_1\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__34397\,
            I => \r_SM_Main_1\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__34394\,
            I => \r_SM_Main_1\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__34389\,
            I => \r_SM_Main_1\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__34384\,
            I => \r_SM_Main_1\
        );

    \I__8365\ : Odrv4
    port map (
            O => \N__34381\,
            I => \r_SM_Main_1\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__34376\,
            I => \r_SM_Main_1\
        );

    \I__8363\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34356\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__34356\,
            I => n9259
        );

    \I__8361\ : CascadeMux
    port map (
            O => \N__34353\,
            I => \N__34344\
        );

    \I__8360\ : CascadeMux
    port map (
            O => \N__34352\,
            I => \N__34341\
        );

    \I__8359\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34329\
        );

    \I__8358\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34322\
        );

    \I__8357\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34322\
        );

    \I__8356\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34322\
        );

    \I__8355\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34319\
        );

    \I__8354\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34308\
        );

    \I__8353\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34308\
        );

    \I__8352\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34308\
        );

    \I__8351\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34308\
        );

    \I__8350\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34308\
        );

    \I__8349\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34295\
        );

    \I__8348\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34295\
        );

    \I__8347\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34295\
        );

    \I__8346\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34295\
        );

    \I__8345\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34295\
        );

    \I__8344\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34295\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__34329\,
            I => \c0.n123\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__34322\,
            I => \c0.n123\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__34319\,
            I => \c0.n123\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__34308\,
            I => \c0.n123\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__34295\,
            I => \c0.n123\
        );

    \I__8338\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34268\
        );

    \I__8337\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34265\
        );

    \I__8336\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34254\
        );

    \I__8335\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34254\
        );

    \I__8334\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34254\
        );

    \I__8333\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34254\
        );

    \I__8332\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34254\
        );

    \I__8331\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34239\
        );

    \I__8330\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34239\
        );

    \I__8329\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34239\
        );

    \I__8328\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34239\
        );

    \I__8327\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34239\
        );

    \I__8326\ : InMux
    port map (
            O => \N__34272\,
            I => \N__34239\
        );

    \I__8325\ : InMux
    port map (
            O => \N__34271\,
            I => \N__34239\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__34268\,
            I => \c0.n7814\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__34265\,
            I => \c0.n7814\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__34254\,
            I => \c0.n7814\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__34239\,
            I => \c0.n7814\
        );

    \I__8320\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34227\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__34224\,
            I => \c0.n117\
        );

    \I__8317\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34213\
        );

    \I__8316\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34213\
        );

    \I__8315\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34208\
        );

    \I__8314\ : InMux
    port map (
            O => \N__34218\,
            I => \N__34208\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__34213\,
            I => \N__34204\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34201\
        );

    \I__8311\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34197\
        );

    \I__8310\ : Span4Mux_v
    port map (
            O => \N__34204\,
            I => \N__34192\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__34201\,
            I => \N__34189\
        );

    \I__8308\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34186\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__34197\,
            I => \N__34183\
        );

    \I__8306\ : InMux
    port map (
            O => \N__34196\,
            I => \N__34178\
        );

    \I__8305\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34178\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__34192\,
            I => n3747
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__34189\,
            I => n3747
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__34186\,
            I => n3747
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__34183\,
            I => n3747
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__34178\,
            I => n3747
        );

    \I__8299\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34164\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__34164\,
            I => \c0.tx_active_prev\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__34161\,
            I => \n8749_cascade_\
        );

    \I__8296\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34150\
        );

    \I__8295\ : InMux
    port map (
            O => \N__34157\,
            I => \N__34147\
        );

    \I__8294\ : InMux
    port map (
            O => \N__34156\,
            I => \N__34140\
        );

    \I__8293\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34140\
        );

    \I__8292\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34140\
        );

    \I__8291\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34137\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__34150\,
            I => tx_active
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__34147\,
            I => tx_active
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__34140\,
            I => tx_active
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__34137\,
            I => tx_active
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__34128\,
            I => \c0.tx.n8_cascade_\
        );

    \I__8285\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__34122\,
            I => \c0.n19_adj_1664\
        );

    \I__8283\ : IoInMux
    port map (
            O => \N__34119\,
            I => \N__34116\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__34116\,
            I => \N__34113\
        );

    \I__8281\ : Span4Mux_s0_v
    port map (
            O => \N__34113\,
            I => \N__34109\
        );

    \I__8280\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34106\
        );

    \I__8279\ : Span4Mux_h
    port map (
            O => \N__34109\,
            I => \N__34101\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__34106\,
            I => \N__34101\
        );

    \I__8277\ : Span4Mux_h
    port map (
            O => \N__34101\,
            I => \N__34098\
        );

    \I__8276\ : Span4Mux_v
    port map (
            O => \N__34098\,
            I => \N__34094\
        );

    \I__8275\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34091\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__34094\,
            I => tx_o_adj_1726
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__34091\,
            I => tx_o_adj_1726
        );

    \I__8272\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34083\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__34083\,
            I => n9452
        );

    \I__8270\ : CascadeMux
    port map (
            O => \N__34080\,
            I => \N__34076\
        );

    \I__8269\ : InMux
    port map (
            O => \N__34079\,
            I => \N__34073\
        );

    \I__8268\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34070\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__34073\,
            I => \r_Tx_Data_0\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__34070\,
            I => \r_Tx_Data_0\
        );

    \I__8265\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34062\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__34062\,
            I => n9455
        );

    \I__8263\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34056\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__34056\,
            I => \tx_data_4_N_keep\
        );

    \I__8261\ : InMux
    port map (
            O => \N__34053\,
            I => \N__34047\
        );

    \I__8260\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34047\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__34047\,
            I => \r_Tx_Data_4\
        );

    \I__8258\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34038\
        );

    \I__8257\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34038\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__34038\,
            I => n9073
        );

    \I__8255\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34028\
        );

    \I__8254\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34025\
        );

    \I__8253\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34022\
        );

    \I__8252\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34017\
        );

    \I__8251\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34017\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__34028\,
            I => \r_Bit_Index_0\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__34025\,
            I => \r_Bit_Index_0\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__34022\,
            I => \r_Bit_Index_0\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__34017\,
            I => \r_Bit_Index_0\
        );

    \I__8246\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__34000\
        );

    \I__8244\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33995\
        );

    \I__8243\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33995\
        );

    \I__8242\ : Odrv4
    port map (
            O => \N__34000\,
            I => n5062
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__33995\,
            I => n5062
        );

    \I__8240\ : CascadeMux
    port map (
            O => \N__33990\,
            I => \n9073_cascade_\
        );

    \I__8239\ : CascadeMux
    port map (
            O => \N__33987\,
            I => \N__33981\
        );

    \I__8238\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33977\
        );

    \I__8237\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33974\
        );

    \I__8236\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33969\
        );

    \I__8235\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33966\
        );

    \I__8234\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33963\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__33977\,
            I => \N__33958\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__33974\,
            I => \N__33958\
        );

    \I__8231\ : InMux
    port map (
            O => \N__33973\,
            I => \N__33953\
        );

    \I__8230\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33953\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__33969\,
            I => \N__33950\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__33966\,
            I => \N__33947\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__33963\,
            I => \r_Bit_Index_1\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__33958\,
            I => \r_Bit_Index_1\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__33953\,
            I => \r_Bit_Index_1\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__33950\,
            I => \r_Bit_Index_1\
        );

    \I__8223\ : Odrv4
    port map (
            O => \N__33947\,
            I => \r_Bit_Index_1\
        );

    \I__8222\ : CascadeMux
    port map (
            O => \N__33936\,
            I => \N__33933\
        );

    \I__8221\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__33930\,
            I => n3892
        );

    \I__8219\ : InMux
    port map (
            O => \N__33927\,
            I => \N__33924\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__33924\,
            I => \c0.n18_adj_1662\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__33921\,
            I => \N__33914\
        );

    \I__8216\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33907\
        );

    \I__8215\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33900\
        );

    \I__8214\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33900\
        );

    \I__8213\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33900\
        );

    \I__8212\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33897\
        );

    \I__8211\ : InMux
    port map (
            O => \N__33913\,
            I => \N__33893\
        );

    \I__8210\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33890\
        );

    \I__8209\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33885\
        );

    \I__8208\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33885\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__33907\,
            I => \N__33878\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__33900\,
            I => \N__33878\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__33897\,
            I => \N__33878\
        );

    \I__8204\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33875\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__33893\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__33890\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__33885\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__33878\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__33875\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__33864\,
            I => \c0.n7779_cascade_\
        );

    \I__8197\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33857\
        );

    \I__8196\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33854\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__33857\,
            I => \tx_data_1_N_keep\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__33854\,
            I => \tx_data_1_N_keep\
        );

    \I__8193\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__33846\,
            I => \c0.data_out_6__7__N_973\
        );

    \I__8191\ : InMux
    port map (
            O => \N__33843\,
            I => \N__33839\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__33842\,
            I => \N__33832\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__33839\,
            I => \N__33829\
        );

    \I__8188\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33824\
        );

    \I__8187\ : InMux
    port map (
            O => \N__33837\,
            I => \N__33824\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__33836\,
            I => \N__33817\
        );

    \I__8185\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33814\
        );

    \I__8184\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33811\
        );

    \I__8183\ : Span4Mux_v
    port map (
            O => \N__33829\,
            I => \N__33806\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__33824\,
            I => \N__33806\
        );

    \I__8181\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33801\
        );

    \I__8180\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33801\
        );

    \I__8179\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33796\
        );

    \I__8178\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33796\
        );

    \I__8177\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33793\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__33814\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__33811\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8174\ : Odrv4
    port map (
            O => \N__33806\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__33801\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__33796\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__33793\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__8170\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33771\
        );

    \I__8169\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33771\
        );

    \I__8168\ : InMux
    port map (
            O => \N__33778\,
            I => \N__33767\
        );

    \I__8167\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33762\
        );

    \I__8166\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33762\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__33771\,
            I => \N__33759\
        );

    \I__8164\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33755\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__33767\,
            I => \N__33750\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33750\
        );

    \I__8161\ : Span4Mux_v
    port map (
            O => \N__33759\,
            I => \N__33747\
        );

    \I__8160\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33744\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__33755\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__33750\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__33747\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__33744\,
            I => \c0.byte_transmit_counter_4\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__8154\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33728\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__33731\,
            I => \N__33720\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33716\
        );

    \I__8151\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33713\
        );

    \I__8150\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33706\
        );

    \I__8149\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33706\
        );

    \I__8148\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33706\
        );

    \I__8147\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33701\
        );

    \I__8146\ : InMux
    port map (
            O => \N__33720\,
            I => \N__33701\
        );

    \I__8145\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33697\
        );

    \I__8144\ : Span4Mux_v
    port map (
            O => \N__33716\,
            I => \N__33688\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__33713\,
            I => \N__33688\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__33706\,
            I => \N__33688\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__33701\,
            I => \N__33688\
        );

    \I__8140\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33685\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__33697\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__33688\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__33685\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__8136\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33666\
        );

    \I__8135\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33666\
        );

    \I__8134\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33666\
        );

    \I__8133\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33661\
        );

    \I__8132\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33661\
        );

    \I__8131\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33657\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33654\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33651\
        );

    \I__8128\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33648\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__33657\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8126\ : Odrv4
    port map (
            O => \N__33654\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8125\ : Odrv4
    port map (
            O => \N__33651\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__33648\,
            I => \c0.byte_transmit_counter_3\
        );

    \I__8123\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__33636\,
            I => \c0.n9291\
        );

    \I__8121\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33629\
        );

    \I__8120\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33626\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33623\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__33626\,
            I => \r_Tx_Data_3\
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__33623\,
            I => \r_Tx_Data_3\
        );

    \I__8116\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__33615\,
            I => \tx_data_7_N_keep\
        );

    \I__8114\ : CascadeMux
    port map (
            O => \N__33612\,
            I => \N__33608\
        );

    \I__8113\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33603\
        );

    \I__8112\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33603\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__33603\,
            I => \r_Tx_Data_7\
        );

    \I__8110\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33596\
        );

    \I__8109\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33593\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33590\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__33593\,
            I => \r_Tx_Data_1\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__33590\,
            I => \r_Tx_Data_1\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__33585\,
            I => \N__33581\
        );

    \I__8104\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33578\
        );

    \I__8103\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33575\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__33578\,
            I => \r_Tx_Data_5\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__33575\,
            I => \r_Tx_Data_5\
        );

    \I__8100\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__33567\,
            I => n9710
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__33564\,
            I => \n9713_cascade_\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__33561\,
            I => \n5_cascade_\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__33558\,
            I => \n3_cascade_\
        );

    \I__8095\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33551\
        );

    \I__8094\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33548\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__33551\,
            I => \c0.data_out_6_7_N_965_6\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__33548\,
            I => \c0.data_out_6_7_N_965_6\
        );

    \I__8091\ : InMux
    port map (
            O => \N__33543\,
            I => \N__33539\
        );

    \I__8090\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33536\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__33539\,
            I => \c0.data_out_6_7_N_965_4\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__33536\,
            I => \c0.data_out_6_7_N_965_4\
        );

    \I__8087\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33527\
        );

    \I__8086\ : InMux
    port map (
            O => \N__33530\,
            I => \N__33524\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__33527\,
            I => \c0.data_out_6_7_N_965_7\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__33524\,
            I => \c0.data_out_6_7_N_965_7\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__33519\,
            I => \c0.n7_cascade_\
        );

    \I__8082\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__33513\,
            I => \c0.n8\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__33510\,
            I => \c0.n7814_cascade_\
        );

    \I__8079\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33501\
        );

    \I__8078\ : InMux
    port map (
            O => \N__33506\,
            I => \N__33501\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__33501\,
            I => \data_out_6_7_N_965_5\
        );

    \I__8076\ : CascadeMux
    port map (
            O => \N__33498\,
            I => \n7204_cascade_\
        );

    \I__8075\ : InMux
    port map (
            O => \N__33495\,
            I => \N__33491\
        );

    \I__8074\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33488\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__33491\,
            I => byte_transmit_counter_5
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__33488\,
            I => byte_transmit_counter_5
        );

    \I__8071\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33477\
        );

    \I__8070\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33477\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__33477\,
            I => \c0.data_out_6_7_N_965_1\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__33474\,
            I => \N__33470\
        );

    \I__8067\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33466\
        );

    \I__8066\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33461\
        );

    \I__8065\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33461\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__33466\,
            I => n7204
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__33461\,
            I => n7204
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__33456\,
            I => \tx_data_1_N_keep_cascade_\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__33453\,
            I => \c0.n17_adj_1663_cascade_\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__33450\,
            I => \c0.n123_cascade_\
        );

    \I__8059\ : CascadeMux
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__8058\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33440\
        );

    \I__8057\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33437\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__33440\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__33437\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__8054\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33428\
        );

    \I__8053\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33425\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__33428\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__33425\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__8050\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33416\
        );

    \I__8049\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33413\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__33416\,
            I => \c0.data_out_6_7_N_965_3\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__33413\,
            I => \c0.data_out_6_7_N_965_3\
        );

    \I__8046\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33404\
        );

    \I__8045\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33401\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__33404\,
            I => \c0.data_out_6_7_N_965_2\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__33401\,
            I => \c0.data_out_6_7_N_965_2\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__33396\,
            I => \N__33392\
        );

    \I__8041\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33387\
        );

    \I__8040\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33387\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__33387\,
            I => \c0.data_out_6_7_N_965_0\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__33384\,
            I => \tx_data_5_N_keep_cascade_\
        );

    \I__8037\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33376\
        );

    \I__8036\ : CascadeMux
    port map (
            O => \N__33380\,
            I => \N__33372\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__33379\,
            I => \N__33369\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__33376\,
            I => \N__33366\
        );

    \I__8033\ : InMux
    port map (
            O => \N__33375\,
            I => \N__33363\
        );

    \I__8032\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33358\
        );

    \I__8031\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33358\
        );

    \I__8030\ : Odrv12
    port map (
            O => \N__33366\,
            I => \c0.n11\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__33363\,
            I => \c0.n11\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__33358\,
            I => \c0.n11\
        );

    \I__8027\ : CascadeMux
    port map (
            O => \N__33351\,
            I => \tx_data_2_N_keep_cascade_\
        );

    \I__8026\ : InMux
    port map (
            O => \N__33348\,
            I => \N__33345\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__33345\,
            I => \tx_data_6_N_keep\
        );

    \I__8024\ : CascadeMux
    port map (
            O => \N__33342\,
            I => \n8705_cascade_\
        );

    \I__8023\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33333\
        );

    \I__8022\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33333\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__33333\,
            I => \r_Tx_Data_6\
        );

    \I__8020\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33324\
        );

    \I__8019\ : InMux
    port map (
            O => \N__33329\,
            I => \N__33324\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__33324\,
            I => \r_Tx_Data_2\
        );

    \I__8017\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__8015\ : Span4Mux_s2_v
    port map (
            O => \N__33315\,
            I => \N__33310\
        );

    \I__8014\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33307\
        );

    \I__8013\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33304\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__33310\,
            I => \N__33297\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__33307\,
            I => \N__33297\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__33304\,
            I => \N__33294\
        );

    \I__8009\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33291\
        );

    \I__8008\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33288\
        );

    \I__8007\ : Span4Mux_v
    port map (
            O => \N__33297\,
            I => \N__33285\
        );

    \I__8006\ : Span4Mux_h
    port map (
            O => \N__33294\,
            I => \N__33280\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__33291\,
            I => \N__33280\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__33288\,
            I => data_in_field_132
        );

    \I__8003\ : Odrv4
    port map (
            O => \N__33285\,
            I => data_in_field_132
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__33280\,
            I => data_in_field_132
        );

    \I__8001\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33270\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__33270\,
            I => \N__33267\
        );

    \I__7999\ : Span4Mux_s2_v
    port map (
            O => \N__33267\,
            I => \N__33264\
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__33264\,
            I => \c0.n9680\
        );

    \I__7997\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33258\
        );

    \I__7996\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33254\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__33257\,
            I => \N__33251\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33248\
        );

    \I__7993\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33244\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__33248\,
            I => \N__33241\
        );

    \I__7991\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33238\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__33244\,
            I => \N__33235\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__33241\,
            I => \N__33228\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33228\
        );

    \I__7987\ : Span4Mux_v
    port map (
            O => \N__33235\,
            I => \N__33225\
        );

    \I__7986\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33220\
        );

    \I__7985\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33220\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__33228\,
            I => \N__33217\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__33225\,
            I => data_in_field_140
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__33220\,
            I => data_in_field_140
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__33217\,
            I => data_in_field_140
        );

    \I__7980\ : CascadeMux
    port map (
            O => \N__33210\,
            I => \N__33205\
        );

    \I__7979\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33194\
        );

    \I__7978\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33194\
        );

    \I__7977\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33186\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__33204\,
            I => \N__33183\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__33203\,
            I => \N__33178\
        );

    \I__7974\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33164\
        );

    \I__7973\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33164\
        );

    \I__7972\ : InMux
    port map (
            O => \N__33200\,
            I => \N__33164\
        );

    \I__7971\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33164\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33161\
        );

    \I__7969\ : InMux
    port map (
            O => \N__33193\,
            I => \N__33152\
        );

    \I__7968\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33152\
        );

    \I__7967\ : InMux
    port map (
            O => \N__33191\,
            I => \N__33152\
        );

    \I__7966\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33152\
        );

    \I__7965\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33145\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33142\
        );

    \I__7963\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33139\
        );

    \I__7962\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33130\
        );

    \I__7961\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33130\
        );

    \I__7960\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33125\
        );

    \I__7959\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33125\
        );

    \I__7958\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33122\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__33175\,
            I => \N__33117\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__33174\,
            I => \N__33112\
        );

    \I__7955\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33109\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__33164\,
            I => \N__33102\
        );

    \I__7953\ : Span4Mux_v
    port map (
            O => \N__33161\,
            I => \N__33102\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__33152\,
            I => \N__33102\
        );

    \I__7951\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33099\
        );

    \I__7950\ : CascadeMux
    port map (
            O => \N__33150\,
            I => \N__33092\
        );

    \I__7949\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33085\
        );

    \I__7948\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33085\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33082\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__33142\,
            I => \N__33077\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__33139\,
            I => \N__33077\
        );

    \I__7944\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33074\
        );

    \I__7943\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33071\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__33136\,
            I => \N__33068\
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \N__33065\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__33130\,
            I => \N__33057\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__33125\,
            I => \N__33057\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__33122\,
            I => \N__33057\
        );

    \I__7937\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33054\
        );

    \I__7936\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33047\
        );

    \I__7935\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33047\
        );

    \I__7934\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33047\
        );

    \I__7933\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33042\
        );

    \I__7932\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33042\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__33109\,
            I => \N__33035\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__33102\,
            I => \N__33035\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33035\
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__33098\,
            I => \N__33025\
        );

    \I__7927\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33020\
        );

    \I__7926\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33015\
        );

    \I__7925\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33009\
        );

    \I__7924\ : InMux
    port map (
            O => \N__33092\,
            I => \N__33009\
        );

    \I__7923\ : InMux
    port map (
            O => \N__33091\,
            I => \N__33006\
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__33090\,
            I => \N__33003\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__33085\,
            I => \N__33000\
        );

    \I__7920\ : Span4Mux_h
    port map (
            O => \N__33082\,
            I => \N__32995\
        );

    \I__7919\ : Span4Mux_h
    port map (
            O => \N__33077\,
            I => \N__32995\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__33074\,
            I => \N__32992\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__33071\,
            I => \N__32989\
        );

    \I__7916\ : InMux
    port map (
            O => \N__33068\,
            I => \N__32982\
        );

    \I__7915\ : InMux
    port map (
            O => \N__33065\,
            I => \N__32979\
        );

    \I__7914\ : InMux
    port map (
            O => \N__33064\,
            I => \N__32975\
        );

    \I__7913\ : Span4Mux_v
    port map (
            O => \N__33057\,
            I => \N__32966\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__32966\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__33047\,
            I => \N__32966\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__33042\,
            I => \N__32966\
        );

    \I__7909\ : Span4Mux_v
    port map (
            O => \N__33035\,
            I => \N__32963\
        );

    \I__7908\ : InMux
    port map (
            O => \N__33034\,
            I => \N__32958\
        );

    \I__7907\ : InMux
    port map (
            O => \N__33033\,
            I => \N__32958\
        );

    \I__7906\ : CascadeMux
    port map (
            O => \N__33032\,
            I => \N__32952\
        );

    \I__7905\ : CascadeMux
    port map (
            O => \N__33031\,
            I => \N__32949\
        );

    \I__7904\ : InMux
    port map (
            O => \N__33030\,
            I => \N__32936\
        );

    \I__7903\ : InMux
    port map (
            O => \N__33029\,
            I => \N__32936\
        );

    \I__7902\ : InMux
    port map (
            O => \N__33028\,
            I => \N__32936\
        );

    \I__7901\ : InMux
    port map (
            O => \N__33025\,
            I => \N__32936\
        );

    \I__7900\ : CascadeMux
    port map (
            O => \N__33024\,
            I => \N__32933\
        );

    \I__7899\ : InMux
    port map (
            O => \N__33023\,
            I => \N__32930\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__33020\,
            I => \N__32927\
        );

    \I__7897\ : InMux
    port map (
            O => \N__33019\,
            I => \N__32922\
        );

    \I__7896\ : InMux
    port map (
            O => \N__33018\,
            I => \N__32922\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__32919\
        );

    \I__7894\ : CascadeMux
    port map (
            O => \N__33014\,
            I => \N__32915\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__33009\,
            I => \N__32912\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__32909\
        );

    \I__7891\ : InMux
    port map (
            O => \N__33003\,
            I => \N__32906\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__33000\,
            I => \N__32899\
        );

    \I__7889\ : Span4Mux_v
    port map (
            O => \N__32995\,
            I => \N__32899\
        );

    \I__7888\ : Span4Mux_h
    port map (
            O => \N__32992\,
            I => \N__32899\
        );

    \I__7887\ : Span4Mux_s3_h
    port map (
            O => \N__32989\,
            I => \N__32896\
        );

    \I__7886\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32893\
        );

    \I__7885\ : CascadeMux
    port map (
            O => \N__32987\,
            I => \N__32886\
        );

    \I__7884\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32878\
        );

    \I__7883\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32878\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32873\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32873\
        );

    \I__7880\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32867\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32860\
        );

    \I__7878\ : Span4Mux_v
    port map (
            O => \N__32966\,
            I => \N__32860\
        );

    \I__7877\ : IoSpan4Mux
    port map (
            O => \N__32963\,
            I => \N__32860\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__32958\,
            I => \N__32857\
        );

    \I__7875\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32852\
        );

    \I__7874\ : InMux
    port map (
            O => \N__32956\,
            I => \N__32852\
        );

    \I__7873\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32843\
        );

    \I__7872\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32843\
        );

    \I__7871\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32840\
        );

    \I__7870\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32835\
        );

    \I__7869\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32835\
        );

    \I__7868\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32832\
        );

    \I__7867\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32829\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__32936\,
            I => \N__32826\
        );

    \I__7865\ : InMux
    port map (
            O => \N__32933\,
            I => \N__32823\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__32930\,
            I => \N__32820\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__32927\,
            I => \N__32815\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32815\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__32919\,
            I => \N__32812\
        );

    \I__7860\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32807\
        );

    \I__7859\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32807\
        );

    \I__7858\ : Span4Mux_v
    port map (
            O => \N__32912\,
            I => \N__32799\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__32909\,
            I => \N__32799\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32799\
        );

    \I__7855\ : IoSpan4Mux
    port map (
            O => \N__32899\,
            I => \N__32796\
        );

    \I__7854\ : Span4Mux_h
    port map (
            O => \N__32896\,
            I => \N__32791\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__32893\,
            I => \N__32791\
        );

    \I__7852\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32786\
        );

    \I__7851\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32783\
        );

    \I__7850\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32780\
        );

    \I__7849\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32775\
        );

    \I__7848\ : InMux
    port map (
            O => \N__32886\,
            I => \N__32775\
        );

    \I__7847\ : InMux
    port map (
            O => \N__32885\,
            I => \N__32770\
        );

    \I__7846\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32770\
        );

    \I__7845\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32767\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__32878\,
            I => \N__32764\
        );

    \I__7843\ : Span4Mux_h
    port map (
            O => \N__32873\,
            I => \N__32761\
        );

    \I__7842\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32758\
        );

    \I__7841\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32755\
        );

    \I__7840\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32752\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32749\
        );

    \I__7838\ : Span4Mux_s2_h
    port map (
            O => \N__32860\,
            I => \N__32742\
        );

    \I__7837\ : Span4Mux_s2_h
    port map (
            O => \N__32857\,
            I => \N__32742\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__32852\,
            I => \N__32742\
        );

    \I__7835\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32733\
        );

    \I__7834\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32733\
        );

    \I__7833\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32733\
        );

    \I__7832\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32733\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32728\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32728\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32709\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__32832\,
            I => \N__32709\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32709\
        );

    \I__7826\ : Span4Mux_s1_v
    port map (
            O => \N__32826\,
            I => \N__32709\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__32823\,
            I => \N__32709\
        );

    \I__7824\ : Span4Mux_h
    port map (
            O => \N__32820\,
            I => \N__32709\
        );

    \I__7823\ : Span4Mux_h
    port map (
            O => \N__32815\,
            I => \N__32709\
        );

    \I__7822\ : Span4Mux_h
    port map (
            O => \N__32812\,
            I => \N__32709\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32709\
        );

    \I__7820\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32706\
        );

    \I__7819\ : Span4Mux_h
    port map (
            O => \N__32799\,
            I => \N__32699\
        );

    \I__7818\ : Span4Mux_s2_v
    port map (
            O => \N__32796\,
            I => \N__32699\
        );

    \I__7817\ : Span4Mux_h
    port map (
            O => \N__32791\,
            I => \N__32699\
        );

    \I__7816\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32696\
        );

    \I__7815\ : InMux
    port map (
            O => \N__32789\,
            I => \N__32693\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__32786\,
            I => \N__32678\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__32783\,
            I => \N__32678\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__32780\,
            I => \N__32678\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__32775\,
            I => \N__32678\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__32770\,
            I => \N__32678\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__32767\,
            I => \N__32678\
        );

    \I__7808\ : Span12Mux_s1_h
    port map (
            O => \N__32764\,
            I => \N__32678\
        );

    \I__7807\ : Span4Mux_v
    port map (
            O => \N__32761\,
            I => \N__32675\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__32758\,
            I => \N__32668\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__32755\,
            I => \N__32668\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__32752\,
            I => \N__32668\
        );

    \I__7803\ : Span4Mux_h
    port map (
            O => \N__32749\,
            I => \N__32663\
        );

    \I__7802\ : Span4Mux_h
    port map (
            O => \N__32742\,
            I => \N__32663\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__32733\,
            I => \N__32656\
        );

    \I__7800\ : Span12Mux_s6_h
    port map (
            O => \N__32728\,
            I => \N__32656\
        );

    \I__7799\ : Sp12to4
    port map (
            O => \N__32709\,
            I => \N__32656\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__32706\,
            I => \N__32653\
        );

    \I__7797\ : Span4Mux_v
    port map (
            O => \N__32699\,
            I => \N__32650\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__32696\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__32693\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7794\ : Odrv12
    port map (
            O => \N__32678\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__32675\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7792\ : Odrv4
    port map (
            O => \N__32668\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7791\ : Odrv4
    port map (
            O => \N__32663\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7790\ : Odrv12
    port map (
            O => \N__32656\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7789\ : Odrv4
    port map (
            O => \N__32653\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7788\ : Odrv4
    port map (
            O => \N__32650\,
            I => \c0.byte_transmit_counter2_1\
        );

    \I__7787\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32628\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__32628\,
            I => \N__32625\
        );

    \I__7785\ : Span4Mux_h
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__32622\,
            I => \c0.n9683\
        );

    \I__7783\ : CascadeMux
    port map (
            O => \N__32619\,
            I => \c0.n11_cascade_\
        );

    \I__7782\ : CascadeMux
    port map (
            O => \N__32616\,
            I => \tx_data_3_N_keep_cascade_\
        );

    \I__7781\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32610\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__32610\,
            I => \tx_data_0_N_keep\
        );

    \I__7779\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32603\
        );

    \I__7778\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32600\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32595\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__32600\,
            I => \N__32592\
        );

    \I__7775\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32587\
        );

    \I__7774\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32587\
        );

    \I__7773\ : Span4Mux_h
    port map (
            O => \N__32595\,
            I => \N__32583\
        );

    \I__7772\ : Span4Mux_h
    port map (
            O => \N__32592\,
            I => \N__32580\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__32587\,
            I => \N__32577\
        );

    \I__7770\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32574\
        );

    \I__7769\ : Span4Mux_h
    port map (
            O => \N__32583\,
            I => \N__32571\
        );

    \I__7768\ : Span4Mux_v
    port map (
            O => \N__32580\,
            I => \N__32568\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__32577\,
            I => \N__32565\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__32574\,
            I => data_in_field_133
        );

    \I__7765\ : Odrv4
    port map (
            O => \N__32571\,
            I => data_in_field_133
        );

    \I__7764\ : Odrv4
    port map (
            O => \N__32568\,
            I => data_in_field_133
        );

    \I__7763\ : Odrv4
    port map (
            O => \N__32565\,
            I => data_in_field_133
        );

    \I__7762\ : InMux
    port map (
            O => \N__32556\,
            I => \N__32551\
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__32555\,
            I => \N__32548\
        );

    \I__7760\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32545\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__32551\,
            I => \N__32542\
        );

    \I__7758\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32539\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32533\
        );

    \I__7756\ : Span4Mux_h
    port map (
            O => \N__32542\,
            I => \N__32533\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32530\
        );

    \I__7754\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32527\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__32533\,
            I => \N__32524\
        );

    \I__7752\ : Span4Mux_h
    port map (
            O => \N__32530\,
            I => \N__32521\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__32527\,
            I => data_in_field_103
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__32524\,
            I => data_in_field_103
        );

    \I__7749\ : Odrv4
    port map (
            O => \N__32521\,
            I => data_in_field_103
        );

    \I__7748\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32510\
        );

    \I__7747\ : InMux
    port map (
            O => \N__32513\,
            I => \N__32504\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32501\
        );

    \I__7745\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32498\
        );

    \I__7744\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32494\
        );

    \I__7743\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32491\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32488\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__32501\,
            I => \N__32485\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__32498\,
            I => \N__32482\
        );

    \I__7739\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32479\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32474\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32474\
        );

    \I__7736\ : Span4Mux_h
    port map (
            O => \N__32488\,
            I => \N__32471\
        );

    \I__7735\ : Span4Mux_v
    port map (
            O => \N__32485\,
            I => \N__32466\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__32482\,
            I => \N__32466\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__32479\,
            I => data_in_field_148
        );

    \I__7732\ : Odrv12
    port map (
            O => \N__32474\,
            I => data_in_field_148
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__32471\,
            I => data_in_field_148
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__32466\,
            I => data_in_field_148
        );

    \I__7729\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__7727\ : Span4Mux_v
    port map (
            O => \N__32451\,
            I => \N__32448\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__32448\,
            I => \N__32444\
        );

    \I__7725\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32441\
        );

    \I__7724\ : Span4Mux_h
    port map (
            O => \N__32444\,
            I => \N__32436\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__32441\,
            I => \N__32436\
        );

    \I__7722\ : Span4Mux_v
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__7721\ : Odrv4
    port map (
            O => \N__32433\,
            I => \c0.n8986\
        );

    \I__7720\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32427\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__32427\,
            I => \c0.n45_adj_1656\
        );

    \I__7718\ : InMux
    port map (
            O => \N__32424\,
            I => \c0.n8083\
        );

    \I__7717\ : InMux
    port map (
            O => \N__32421\,
            I => \c0.n8084\
        );

    \I__7716\ : InMux
    port map (
            O => \N__32418\,
            I => \c0.n8085\
        );

    \I__7715\ : InMux
    port map (
            O => \N__32415\,
            I => \c0.n8086\
        );

    \I__7714\ : InMux
    port map (
            O => \N__32412\,
            I => \c0.n8087\
        );

    \I__7713\ : InMux
    port map (
            O => \N__32409\,
            I => \c0.n8088\
        );

    \I__7712\ : InMux
    port map (
            O => \N__32406\,
            I => \c0.n8089\
        );

    \I__7711\ : InMux
    port map (
            O => \N__32403\,
            I => \N__32400\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32397\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__32397\,
            I => \N__32394\
        );

    \I__7708\ : Odrv4
    port map (
            O => \N__32394\,
            I => \c0.n22_adj_1681\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__32391\,
            I => \c0.n9491_cascade_\
        );

    \I__7706\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32385\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32378\
        );

    \I__7704\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32374\
        );

    \I__7703\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32371\
        );

    \I__7702\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32368\
        );

    \I__7701\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32365\
        );

    \I__7700\ : Span4Mux_s3_v
    port map (
            O => \N__32378\,
            I => \N__32362\
        );

    \I__7699\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32359\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__32374\,
            I => \N__32356\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__32371\,
            I => \N__32353\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32350\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__32365\,
            I => \N__32345\
        );

    \I__7694\ : Sp12to4
    port map (
            O => \N__32362\,
            I => \N__32339\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__32359\,
            I => \N__32339\
        );

    \I__7692\ : Span4Mux_h
    port map (
            O => \N__32356\,
            I => \N__32332\
        );

    \I__7691\ : Span4Mux_s1_v
    port map (
            O => \N__32353\,
            I => \N__32332\
        );

    \I__7690\ : Span4Mux_h
    port map (
            O => \N__32350\,
            I => \N__32332\
        );

    \I__7689\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32329\
        );

    \I__7688\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32326\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__32345\,
            I => \N__32323\
        );

    \I__7686\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32320\
        );

    \I__7685\ : Span12Mux_s6_h
    port map (
            O => \N__32339\,
            I => \N__32310\
        );

    \I__7684\ : Sp12to4
    port map (
            O => \N__32332\,
            I => \N__32310\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__32329\,
            I => \N__32310\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__32326\,
            I => \N__32310\
        );

    \I__7681\ : Sp12to4
    port map (
            O => \N__32323\,
            I => \N__32305\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__32320\,
            I => \N__32305\
        );

    \I__7679\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32302\
        );

    \I__7678\ : Span12Mux_s3_v
    port map (
            O => \N__32310\,
            I => \N__32299\
        );

    \I__7677\ : Odrv12
    port map (
            O => \N__32305\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__32302\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__7675\ : Odrv12
    port map (
            O => \N__32299\,
            I => \c0.byte_transmit_counter2_4\
        );

    \I__7674\ : InMux
    port map (
            O => \N__32292\,
            I => \N__32289\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__32289\,
            I => \N__32286\
        );

    \I__7672\ : Sp12to4
    port map (
            O => \N__32286\,
            I => \N__32283\
        );

    \I__7671\ : Span12Mux_s6_v
    port map (
            O => \N__32283\,
            I => \N__32280\
        );

    \I__7670\ : Odrv12
    port map (
            O => \N__32280\,
            I => \c0.tx2.r_Tx_Data_2\
        );

    \I__7669\ : CEMux
    port map (
            O => \N__32277\,
            I => \N__32274\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__32274\,
            I => \N__32268\
        );

    \I__7667\ : CEMux
    port map (
            O => \N__32273\,
            I => \N__32265\
        );

    \I__7666\ : CEMux
    port map (
            O => \N__32272\,
            I => \N__32261\
        );

    \I__7665\ : CEMux
    port map (
            O => \N__32271\,
            I => \N__32258\
        );

    \I__7664\ : IoSpan4Mux
    port map (
            O => \N__32268\,
            I => \N__32255\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32252\
        );

    \I__7662\ : CEMux
    port map (
            O => \N__32264\,
            I => \N__32249\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__32261\,
            I => \N__32246\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__32258\,
            I => \N__32243\
        );

    \I__7659\ : Span4Mux_s0_v
    port map (
            O => \N__32255\,
            I => \N__32240\
        );

    \I__7658\ : Span4Mux_v
    port map (
            O => \N__32252\,
            I => \N__32237\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__32249\,
            I => \N__32234\
        );

    \I__7656\ : Span4Mux_v
    port map (
            O => \N__32246\,
            I => \N__32230\
        );

    \I__7655\ : Span4Mux_v
    port map (
            O => \N__32243\,
            I => \N__32225\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__32240\,
            I => \N__32218\
        );

    \I__7653\ : Span4Mux_s1_h
    port map (
            O => \N__32237\,
            I => \N__32218\
        );

    \I__7652\ : Span4Mux_v
    port map (
            O => \N__32234\,
            I => \N__32218\
        );

    \I__7651\ : CEMux
    port map (
            O => \N__32233\,
            I => \N__32215\
        );

    \I__7650\ : Span4Mux_v
    port map (
            O => \N__32230\,
            I => \N__32212\
        );

    \I__7649\ : CEMux
    port map (
            O => \N__32229\,
            I => \N__32209\
        );

    \I__7648\ : CEMux
    port map (
            O => \N__32228\,
            I => \N__32206\
        );

    \I__7647\ : Span4Mux_v
    port map (
            O => \N__32225\,
            I => \N__32203\
        );

    \I__7646\ : Span4Mux_h
    port map (
            O => \N__32218\,
            I => \N__32198\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__32215\,
            I => \N__32198\
        );

    \I__7644\ : Span4Mux_h
    port map (
            O => \N__32212\,
            I => \N__32193\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32193\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__32206\,
            I => \N__32190\
        );

    \I__7641\ : Sp12to4
    port map (
            O => \N__32203\,
            I => \N__32185\
        );

    \I__7640\ : Sp12to4
    port map (
            O => \N__32198\,
            I => \N__32185\
        );

    \I__7639\ : Span4Mux_h
    port map (
            O => \N__32193\,
            I => \N__32182\
        );

    \I__7638\ : Sp12to4
    port map (
            O => \N__32190\,
            I => \N__32179\
        );

    \I__7637\ : Odrv12
    port map (
            O => \N__32185\,
            I => \c0.tx2.n3760\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__32182\,
            I => \c0.tx2.n3760\
        );

    \I__7635\ : Odrv12
    port map (
            O => \N__32179\,
            I => \c0.tx2.n3760\
        );

    \I__7634\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32168\
        );

    \I__7633\ : InMux
    port map (
            O => \N__32171\,
            I => \N__32165\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32161\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__32165\,
            I => \N__32155\
        );

    \I__7630\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32152\
        );

    \I__7629\ : Span4Mux_v
    port map (
            O => \N__32161\,
            I => \N__32149\
        );

    \I__7628\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32146\
        );

    \I__7627\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32143\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32140\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__32155\,
            I => \N__32137\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__32152\,
            I => \N__32128\
        );

    \I__7623\ : Sp12to4
    port map (
            O => \N__32149\,
            I => \N__32128\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__32146\,
            I => \N__32128\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32128\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__32140\,
            I => data_in_field_82
        );

    \I__7619\ : Odrv4
    port map (
            O => \N__32137\,
            I => data_in_field_82
        );

    \I__7618\ : Odrv12
    port map (
            O => \N__32128\,
            I => data_in_field_82
        );

    \I__7617\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32113\
        );

    \I__7616\ : CascadeMux
    port map (
            O => \N__32120\,
            I => \N__32110\
        );

    \I__7615\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32105\
        );

    \I__7614\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32105\
        );

    \I__7613\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32101\
        );

    \I__7612\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32098\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32095\
        );

    \I__7610\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32092\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32089\
        );

    \I__7608\ : InMux
    port map (
            O => \N__32104\,
            I => \N__32086\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__32101\,
            I => \N__32081\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__32098\,
            I => \N__32081\
        );

    \I__7605\ : Span4Mux_s2_v
    port map (
            O => \N__32095\,
            I => \N__32078\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__32092\,
            I => \N__32075\
        );

    \I__7603\ : Span4Mux_h
    port map (
            O => \N__32089\,
            I => \N__32072\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32063\
        );

    \I__7601\ : Span4Mux_v
    port map (
            O => \N__32081\,
            I => \N__32063\
        );

    \I__7600\ : Span4Mux_v
    port map (
            O => \N__32078\,
            I => \N__32063\
        );

    \I__7599\ : Span4Mux_h
    port map (
            O => \N__32075\,
            I => \N__32063\
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__32072\,
            I => data_in_field_90
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__32063\,
            I => data_in_field_90
        );

    \I__7596\ : InMux
    port map (
            O => \N__32058\,
            I => \N__32047\
        );

    \I__7595\ : InMux
    port map (
            O => \N__32057\,
            I => \N__32047\
        );

    \I__7594\ : InMux
    port map (
            O => \N__32056\,
            I => \N__32027\
        );

    \I__7593\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32022\
        );

    \I__7592\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32022\
        );

    \I__7591\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32017\
        );

    \I__7590\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32017\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32008\
        );

    \I__7588\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32004\
        );

    \I__7587\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32001\
        );

    \I__7586\ : InMux
    port map (
            O => \N__32044\,
            I => \N__31997\
        );

    \I__7585\ : InMux
    port map (
            O => \N__32043\,
            I => \N__31994\
        );

    \I__7584\ : InMux
    port map (
            O => \N__32042\,
            I => \N__31987\
        );

    \I__7583\ : InMux
    port map (
            O => \N__32041\,
            I => \N__31987\
        );

    \I__7582\ : InMux
    port map (
            O => \N__32040\,
            I => \N__31984\
        );

    \I__7581\ : InMux
    port map (
            O => \N__32039\,
            I => \N__31981\
        );

    \I__7580\ : InMux
    port map (
            O => \N__32038\,
            I => \N__31978\
        );

    \I__7579\ : InMux
    port map (
            O => \N__32037\,
            I => \N__31972\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__32036\,
            I => \N__31968\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__32035\,
            I => \N__31964\
        );

    \I__7576\ : InMux
    port map (
            O => \N__32034\,
            I => \N__31961\
        );

    \I__7575\ : InMux
    port map (
            O => \N__32033\,
            I => \N__31956\
        );

    \I__7574\ : InMux
    port map (
            O => \N__32032\,
            I => \N__31956\
        );

    \I__7573\ : InMux
    port map (
            O => \N__32031\,
            I => \N__31953\
        );

    \I__7572\ : InMux
    port map (
            O => \N__32030\,
            I => \N__31949\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__31946\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__32022\,
            I => \N__31943\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__32017\,
            I => \N__31940\
        );

    \I__7568\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31937\
        );

    \I__7567\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31934\
        );

    \I__7566\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31931\
        );

    \I__7565\ : InMux
    port map (
            O => \N__32013\,
            I => \N__31928\
        );

    \I__7564\ : InMux
    port map (
            O => \N__32012\,
            I => \N__31923\
        );

    \I__7563\ : InMux
    port map (
            O => \N__32011\,
            I => \N__31923\
        );

    \I__7562\ : Span4Mux_s3_v
    port map (
            O => \N__32008\,
            I => \N__31920\
        );

    \I__7561\ : InMux
    port map (
            O => \N__32007\,
            I => \N__31917\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__31914\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31911\
        );

    \I__7558\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31907\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__31997\,
            I => \N__31904\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__31994\,
            I => \N__31901\
        );

    \I__7555\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31898\
        );

    \I__7554\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31894\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__31987\,
            I => \N__31889\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__31984\,
            I => \N__31889\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__31981\,
            I => \N__31884\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__31978\,
            I => \N__31884\
        );

    \I__7549\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31881\
        );

    \I__7548\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31878\
        );

    \I__7547\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31875\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__31972\,
            I => \N__31872\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__31971\,
            I => \N__31869\
        );

    \I__7544\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31866\
        );

    \I__7543\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31863\
        );

    \I__7542\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31860\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31853\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__31956\,
            I => \N__31853\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__31953\,
            I => \N__31853\
        );

    \I__7538\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31850\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31837\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__31946\,
            I => \N__31837\
        );

    \I__7535\ : Span4Mux_s1_v
    port map (
            O => \N__31943\,
            I => \N__31837\
        );

    \I__7534\ : Span4Mux_s1_v
    port map (
            O => \N__31940\,
            I => \N__31837\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31837\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__31934\,
            I => \N__31837\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31834\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31829\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__31923\,
            I => \N__31829\
        );

    \I__7528\ : Span4Mux_h
    port map (
            O => \N__31920\,
            I => \N__31820\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__31917\,
            I => \N__31820\
        );

    \I__7526\ : Span4Mux_s3_v
    port map (
            O => \N__31914\,
            I => \N__31820\
        );

    \I__7525\ : Span4Mux_s3_v
    port map (
            O => \N__31911\,
            I => \N__31820\
        );

    \I__7524\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31817\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__31907\,
            I => \N__31814\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__31904\,
            I => \N__31807\
        );

    \I__7521\ : Span4Mux_h
    port map (
            O => \N__31901\,
            I => \N__31807\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31807\
        );

    \I__7519\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31804\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__31894\,
            I => \N__31797\
        );

    \I__7517\ : Span4Mux_v
    port map (
            O => \N__31889\,
            I => \N__31797\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__31884\,
            I => \N__31797\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__31881\,
            I => \N__31788\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__31878\,
            I => \N__31788\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__31875\,
            I => \N__31788\
        );

    \I__7512\ : Span4Mux_s3_v
    port map (
            O => \N__31872\,
            I => \N__31788\
        );

    \I__7511\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31785\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31776\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31776\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__31860\,
            I => \N__31776\
        );

    \I__7507\ : Span12Mux_s7_v
    port map (
            O => \N__31853\,
            I => \N__31776\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__31850\,
            I => \N__31773\
        );

    \I__7505\ : Span4Mux_v
    port map (
            O => \N__31837\,
            I => \N__31770\
        );

    \I__7504\ : Span4Mux_h
    port map (
            O => \N__31834\,
            I => \N__31763\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__31829\,
            I => \N__31763\
        );

    \I__7502\ : Span4Mux_v
    port map (
            O => \N__31820\,
            I => \N__31763\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__31817\,
            I => \N__31754\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__31814\,
            I => \N__31754\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__31807\,
            I => \N__31754\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31754\
        );

    \I__7497\ : Span4Mux_h
    port map (
            O => \N__31797\,
            I => \N__31749\
        );

    \I__7496\ : Span4Mux_v
    port map (
            O => \N__31788\,
            I => \N__31749\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__31785\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7494\ : Odrv12
    port map (
            O => \N__31776\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__31773\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__31770\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__31763\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__31754\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__31749\,
            I => \c0.byte_transmit_counter2_0\
        );

    \I__7488\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31726\
        );

    \I__7487\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31726\
        );

    \I__7486\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31723\
        );

    \I__7485\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31719\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__31726\,
            I => \N__31716\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31713\
        );

    \I__7482\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31709\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__31719\,
            I => \N__31706\
        );

    \I__7480\ : Span12Mux_s3_h
    port map (
            O => \N__31716\,
            I => \N__31703\
        );

    \I__7479\ : Span4Mux_h
    port map (
            O => \N__31713\,
            I => \N__31700\
        );

    \I__7478\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31697\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__31709\,
            I => data_in_field_66
        );

    \I__7476\ : Odrv4
    port map (
            O => \N__31706\,
            I => data_in_field_66
        );

    \I__7475\ : Odrv12
    port map (
            O => \N__31703\,
            I => data_in_field_66
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__31700\,
            I => data_in_field_66
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__31697\,
            I => data_in_field_66
        );

    \I__7472\ : CascadeMux
    port map (
            O => \N__31686\,
            I => \N__31682\
        );

    \I__7471\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31679\
        );

    \I__7470\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31675\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__31679\,
            I => \N__31670\
        );

    \I__7468\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31667\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__31675\,
            I => \N__31664\
        );

    \I__7466\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31661\
        );

    \I__7465\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31658\
        );

    \I__7464\ : Span12Mux_s8_h
    port map (
            O => \N__31670\,
            I => \N__31655\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31652\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__31664\,
            I => \N__31647\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31647\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__31658\,
            I => data_in_field_74
        );

    \I__7459\ : Odrv12
    port map (
            O => \N__31655\,
            I => data_in_field_74
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__31652\,
            I => data_in_field_74
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__31647\,
            I => data_in_field_74
        );

    \I__7456\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__31635\,
            I => \c0.n9500\
        );

    \I__7454\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31620\
        );

    \I__7453\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31620\
        );

    \I__7452\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31620\
        );

    \I__7451\ : InMux
    port map (
            O => \N__31629\,
            I => \N__31607\
        );

    \I__7450\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31607\
        );

    \I__7449\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31607\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31601\
        );

    \I__7447\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31594\
        );

    \I__7446\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31594\
        );

    \I__7445\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31594\
        );

    \I__7444\ : InMux
    port map (
            O => \N__31616\,
            I => \N__31587\
        );

    \I__7443\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31587\
        );

    \I__7442\ : InMux
    port map (
            O => \N__31614\,
            I => \N__31587\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31580\
        );

    \I__7440\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31573\
        );

    \I__7439\ : InMux
    port map (
            O => \N__31605\,
            I => \N__31573\
        );

    \I__7438\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31573\
        );

    \I__7437\ : Span4Mux_s3_v
    port map (
            O => \N__31601\,
            I => \N__31564\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__31594\,
            I => \N__31564\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__31587\,
            I => \N__31561\
        );

    \I__7434\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31556\
        );

    \I__7433\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31556\
        );

    \I__7432\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31553\
        );

    \I__7431\ : InMux
    port map (
            O => \N__31583\,
            I => \N__31548\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__31580\,
            I => \N__31543\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__31573\,
            I => \N__31543\
        );

    \I__7428\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31536\
        );

    \I__7427\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31536\
        );

    \I__7426\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31536\
        );

    \I__7425\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31533\
        );

    \I__7424\ : Span4Mux_v
    port map (
            O => \N__31564\,
            I => \N__31529\
        );

    \I__7423\ : Span4Mux_s3_v
    port map (
            O => \N__31561\,
            I => \N__31526\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31521\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31521\
        );

    \I__7420\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31516\
        );

    \I__7419\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31516\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__31548\,
            I => \N__31513\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__31543\,
            I => \N__31506\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__31536\,
            I => \N__31506\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__31533\,
            I => \N__31506\
        );

    \I__7414\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31503\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__31529\,
            I => \N__31498\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__31526\,
            I => \N__31498\
        );

    \I__7411\ : Span12Mux_s7_v
    port map (
            O => \N__31521\,
            I => \N__31493\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__31516\,
            I => \N__31493\
        );

    \I__7409\ : Span4Mux_h
    port map (
            O => \N__31513\,
            I => \N__31488\
        );

    \I__7408\ : Span4Mux_v
    port map (
            O => \N__31506\,
            I => \N__31488\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__31503\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__7406\ : Odrv4
    port map (
            O => \N__31498\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__7405\ : Odrv12
    port map (
            O => \N__31493\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__31488\,
            I => \c0.byte_transmit_counter2_3\
        );

    \I__7403\ : CascadeMux
    port map (
            O => \N__31479\,
            I => \c0.n9198_cascade_\
        );

    \I__7402\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__31473\,
            I => \c0.n9488\
        );

    \I__7400\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31466\
        );

    \I__7399\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31463\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__31466\,
            I => \N__31457\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__31463\,
            I => \N__31454\
        );

    \I__7396\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31451\
        );

    \I__7395\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31446\
        );

    \I__7394\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31446\
        );

    \I__7393\ : Span12Mux_h
    port map (
            O => \N__31457\,
            I => \N__31443\
        );

    \I__7392\ : Span4Mux_h
    port map (
            O => \N__31454\,
            I => \N__31436\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__31451\,
            I => \N__31436\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__31446\,
            I => \N__31436\
        );

    \I__7389\ : Odrv12
    port map (
            O => \N__31443\,
            I => data_in_field_98
        );

    \I__7388\ : Odrv4
    port map (
            O => \N__31436\,
            I => data_in_field_98
        );

    \I__7387\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31428\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__31428\,
            I => \N__31425\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__31425\,
            I => \N__31422\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__31422\,
            I => \c0.n9494\
        );

    \I__7383\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31416\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__31416\,
            I => \N__31411\
        );

    \I__7381\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31408\
        );

    \I__7380\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31404\
        );

    \I__7379\ : Span12Mux_s4_v
    port map (
            O => \N__31411\,
            I => \N__31399\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__31408\,
            I => \N__31399\
        );

    \I__7377\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31396\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__31404\,
            I => data_in_field_106
        );

    \I__7375\ : Odrv12
    port map (
            O => \N__31399\,
            I => data_in_field_106
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__31396\,
            I => data_in_field_106
        );

    \I__7373\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__31386\,
            I => \c0.n9201\
        );

    \I__7371\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31373\
        );

    \I__7369\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31370\
        );

    \I__7368\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31367\
        );

    \I__7367\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31364\
        );

    \I__7366\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31361\
        );

    \I__7365\ : Span4Mux_v
    port map (
            O => \N__31373\,
            I => \N__31355\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31355\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__31367\,
            I => \N__31352\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31347\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__31361\,
            I => \N__31347\
        );

    \I__7360\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31344\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__31355\,
            I => \N__31340\
        );

    \I__7358\ : Span4Mux_v
    port map (
            O => \N__31352\,
            I => \N__31337\
        );

    \I__7357\ : Span4Mux_v
    port map (
            O => \N__31347\,
            I => \N__31334\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__31344\,
            I => \N__31331\
        );

    \I__7355\ : InMux
    port map (
            O => \N__31343\,
            I => \N__31328\
        );

    \I__7354\ : Span4Mux_s2_v
    port map (
            O => \N__31340\,
            I => \N__31325\
        );

    \I__7353\ : Span4Mux_v
    port map (
            O => \N__31337\,
            I => \N__31322\
        );

    \I__7352\ : Span4Mux_v
    port map (
            O => \N__31334\,
            I => \N__31319\
        );

    \I__7351\ : Span4Mux_h
    port map (
            O => \N__31331\,
            I => \N__31314\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31314\
        );

    \I__7349\ : Span4Mux_h
    port map (
            O => \N__31325\,
            I => \N__31311\
        );

    \I__7348\ : Span4Mux_s0_v
    port map (
            O => \N__31322\,
            I => \N__31308\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__31319\,
            I => \N__31303\
        );

    \I__7346\ : Span4Mux_v
    port map (
            O => \N__31314\,
            I => \N__31303\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__31311\,
            I => \c0.n3056\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__31308\,
            I => \c0.n3056\
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__31303\,
            I => \c0.n3056\
        );

    \I__7342\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31293\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__31293\,
            I => \N__31290\
        );

    \I__7340\ : Span4Mux_v
    port map (
            O => \N__31290\,
            I => \N__31287\
        );

    \I__7339\ : Span4Mux_h
    port map (
            O => \N__31287\,
            I => \N__31284\
        );

    \I__7338\ : Odrv4
    port map (
            O => \N__31284\,
            I => \c0.n9671\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__31281\,
            I => \N__31278\
        );

    \I__7336\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31275\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31272\
        );

    \I__7334\ : Span4Mux_h
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__7333\ : Span4Mux_h
    port map (
            O => \N__31269\,
            I => \N__31266\
        );

    \I__7332\ : Odrv4
    port map (
            O => \N__31266\,
            I => \c0.data_in_frame_20_6\
        );

    \I__7331\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31260\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__31260\,
            I => \N__31256\
        );

    \I__7329\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31252\
        );

    \I__7328\ : Span4Mux_s1_v
    port map (
            O => \N__31256\,
            I => \N__31249\
        );

    \I__7327\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31246\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31239\
        );

    \I__7325\ : Span4Mux_h
    port map (
            O => \N__31249\,
            I => \N__31234\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31234\
        );

    \I__7323\ : InMux
    port map (
            O => \N__31245\,
            I => \N__31226\
        );

    \I__7322\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31223\
        );

    \I__7321\ : InMux
    port map (
            O => \N__31243\,
            I => \N__31220\
        );

    \I__7320\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31217\
        );

    \I__7319\ : Span4Mux_v
    port map (
            O => \N__31239\,
            I => \N__31214\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__31234\,
            I => \N__31211\
        );

    \I__7317\ : InMux
    port map (
            O => \N__31233\,
            I => \N__31208\
        );

    \I__7316\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31205\
        );

    \I__7315\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31200\
        );

    \I__7314\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31197\
        );

    \I__7313\ : InMux
    port map (
            O => \N__31229\,
            I => \N__31194\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__31226\,
            I => \N__31189\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31186\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__31220\,
            I => \N__31183\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31180\
        );

    \I__7308\ : Sp12to4
    port map (
            O => \N__31214\,
            I => \N__31169\
        );

    \I__7307\ : Sp12to4
    port map (
            O => \N__31211\,
            I => \N__31169\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31169\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__31205\,
            I => \N__31169\
        );

    \I__7304\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31166\
        );

    \I__7303\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31163\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31156\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31156\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31156\
        );

    \I__7299\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31153\
        );

    \I__7298\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31150\
        );

    \I__7297\ : Span4Mux_h
    port map (
            O => \N__31189\,
            I => \N__31141\
        );

    \I__7296\ : Span4Mux_h
    port map (
            O => \N__31186\,
            I => \N__31141\
        );

    \I__7295\ : Span4Mux_s1_v
    port map (
            O => \N__31183\,
            I => \N__31141\
        );

    \I__7294\ : Span4Mux_h
    port map (
            O => \N__31180\,
            I => \N__31141\
        );

    \I__7293\ : InMux
    port map (
            O => \N__31179\,
            I => \N__31138\
        );

    \I__7292\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31135\
        );

    \I__7291\ : Span12Mux_h
    port map (
            O => \N__31169\,
            I => \N__31132\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__31166\,
            I => \N__31123\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31123\
        );

    \I__7288\ : Span12Mux_s7_v
    port map (
            O => \N__31156\,
            I => \N__31123\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__31153\,
            I => \N__31123\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31116\
        );

    \I__7285\ : Sp12to4
    port map (
            O => \N__31141\,
            I => \N__31116\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__31138\,
            I => \N__31116\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__31135\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7282\ : Odrv12
    port map (
            O => \N__31132\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7281\ : Odrv12
    port map (
            O => \N__31123\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7280\ : Odrv12
    port map (
            O => \N__31116\,
            I => \c0.byte_transmit_counter2_2\
        );

    \I__7279\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31104\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__31104\,
            I => \N__31101\
        );

    \I__7277\ : Span4Mux_s1_v
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__31095\,
            I => \c0.n22_adj_1677\
        );

    \I__7274\ : InMux
    port map (
            O => \N__31092\,
            I => \c0.rx.n8101\
        );

    \I__7273\ : InMux
    port map (
            O => \N__31089\,
            I => \c0.rx.n8102\
        );

    \I__7272\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31083\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__7270\ : Span4Mux_h
    port map (
            O => \N__31080\,
            I => \N__31077\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__31077\,
            I => \N__31069\
        );

    \I__7268\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31066\
        );

    \I__7267\ : InMux
    port map (
            O => \N__31075\,
            I => \N__31063\
        );

    \I__7266\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31058\
        );

    \I__7265\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31058\
        );

    \I__7264\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31055\
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__31069\,
            I => \r_Clock_Count_6_adj_1728\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__31066\,
            I => \r_Clock_Count_6_adj_1728\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__31063\,
            I => \r_Clock_Count_6_adj_1728\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__31058\,
            I => \r_Clock_Count_6_adj_1728\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__31055\,
            I => \r_Clock_Count_6_adj_1728\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__7257\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__31038\,
            I => n220
        );

    \I__7255\ : InMux
    port map (
            O => \N__31035\,
            I => \c0.rx.n8103\
        );

    \I__7254\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31029\
        );

    \I__7253\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__7251\ : Span4Mux_h
    port map (
            O => \N__31023\,
            I => \N__31017\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__31022\,
            I => \N__31013\
        );

    \I__7249\ : CascadeMux
    port map (
            O => \N__31021\,
            I => \N__31009\
        );

    \I__7248\ : InMux
    port map (
            O => \N__31020\,
            I => \N__31006\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__31017\,
            I => \N__31003\
        );

    \I__7246\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31000\
        );

    \I__7245\ : InMux
    port map (
            O => \N__31013\,
            I => \N__30997\
        );

    \I__7244\ : InMux
    port map (
            O => \N__31012\,
            I => \N__30992\
        );

    \I__7243\ : InMux
    port map (
            O => \N__31009\,
            I => \N__30992\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__31006\,
            I => \r_Clock_Count_7_adj_1727\
        );

    \I__7241\ : Odrv4
    port map (
            O => \N__31003\,
            I => \r_Clock_Count_7_adj_1727\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__31000\,
            I => \r_Clock_Count_7_adj_1727\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__30997\,
            I => \r_Clock_Count_7_adj_1727\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__30992\,
            I => \r_Clock_Count_7_adj_1727\
        );

    \I__7237\ : InMux
    port map (
            O => \N__30981\,
            I => \c0.rx.n8104\
        );

    \I__7236\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__30975\,
            I => n219
        );

    \I__7234\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__7232\ : Span4Mux_v
    port map (
            O => \N__30966\,
            I => \N__30960\
        );

    \I__7231\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30955\
        );

    \I__7230\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30955\
        );

    \I__7229\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30952\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__30960\,
            I => \N__30947\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__30955\,
            I => \N__30947\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__30952\,
            I => n4084
        );

    \I__7225\ : Odrv4
    port map (
            O => \N__30947\,
            I => n4084
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__7223\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30936\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__30933\,
            I => n221
        );

    \I__7220\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30925\
        );

    \I__7219\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30920\
        );

    \I__7218\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30920\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__30925\,
            I => \r_Clock_Count_5\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__30920\,
            I => \r_Clock_Count_5\
        );

    \I__7215\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30904\
        );

    \I__7214\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30904\
        );

    \I__7213\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30895\
        );

    \I__7212\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30895\
        );

    \I__7211\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30895\
        );

    \I__7210\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30895\
        );

    \I__7209\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30892\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__30904\,
            I => n30
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__30895\,
            I => n30
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__30892\,
            I => n30
        );

    \I__7205\ : CascadeMux
    port map (
            O => \N__30885\,
            I => \N__30882\
        );

    \I__7204\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30879\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__30879\,
            I => n222
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__30876\,
            I => \N__30870\
        );

    \I__7201\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30862\
        );

    \I__7200\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30862\
        );

    \I__7199\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30859\
        );

    \I__7198\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30856\
        );

    \I__7197\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30849\
        );

    \I__7196\ : InMux
    port map (
            O => \N__30868\,
            I => \N__30849\
        );

    \I__7195\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30849\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__30862\,
            I => \N__30846\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__30859\,
            I => n44
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__30856\,
            I => n44
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__30849\,
            I => n44
        );

    \I__7190\ : Odrv4
    port map (
            O => \N__30846\,
            I => n44
        );

    \I__7189\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30832\
        );

    \I__7188\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30827\
        );

    \I__7187\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30827\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__30832\,
            I => \r_Clock_Count_4_adj_1729\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__30827\,
            I => \r_Clock_Count_4_adj_1729\
        );

    \I__7184\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30819\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__7182\ : Span4Mux_v
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__7181\ : Sp12to4
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__7180\ : Odrv12
    port map (
            O => \N__30810\,
            I => \c0.n9192\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__7178\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__7176\ : Span12Mux_h
    port map (
            O => \N__30798\,
            I => \N__30795\
        );

    \I__7175\ : Odrv12
    port map (
            O => \N__30795\,
            I => \c0.n9195\
        );

    \I__7174\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30778\
        );

    \I__7173\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30778\
        );

    \I__7172\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30771\
        );

    \I__7171\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30771\
        );

    \I__7170\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30771\
        );

    \I__7169\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30768\
        );

    \I__7168\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30765\
        );

    \I__7167\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30760\
        );

    \I__7166\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30760\
        );

    \I__7165\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30757\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30752\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__30771\,
            I => \N__30752\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__30768\,
            I => \N__30747\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30747\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__30760\,
            I => \r_SM_Main_1_adj_1735\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30757\,
            I => \r_SM_Main_1_adj_1735\
        );

    \I__7158\ : Odrv12
    port map (
            O => \N__30752\,
            I => \r_SM_Main_1_adj_1735\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__30747\,
            I => \r_SM_Main_1_adj_1735\
        );

    \I__7156\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__30735\,
            I => n9246
        );

    \I__7154\ : CascadeMux
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__7153\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30725\
        );

    \I__7152\ : CascadeMux
    port map (
            O => \N__30728\,
            I => \N__30716\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30711\
        );

    \I__7150\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30708\
        );

    \I__7149\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30703\
        );

    \I__7148\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30703\
        );

    \I__7147\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30700\
        );

    \I__7146\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30697\
        );

    \I__7145\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30690\
        );

    \I__7144\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30690\
        );

    \I__7143\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30690\
        );

    \I__7142\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30687\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__30711\,
            I => \N__30684\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__30708\,
            I => \N__30679\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__30703\,
            I => \N__30679\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__30700\,
            I => \N__30676\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__30697\,
            I => \r_SM_Main_0_adj_1736\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__30690\,
            I => \r_SM_Main_0_adj_1736\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__30687\,
            I => \r_SM_Main_0_adj_1736\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__30684\,
            I => \r_SM_Main_0_adj_1736\
        );

    \I__7133\ : Odrv12
    port map (
            O => \N__30679\,
            I => \r_SM_Main_0_adj_1736\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__30676\,
            I => \r_SM_Main_0_adj_1736\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__30663\,
            I => \n44_cascade_\
        );

    \I__7130\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30652\
        );

    \I__7129\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30652\
        );

    \I__7128\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__30657\,
            I => \N__30643\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30636\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30636\
        );

    \I__7124\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30629\
        );

    \I__7123\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30629\
        );

    \I__7122\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30629\
        );

    \I__7121\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30626\
        );

    \I__7120\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30623\
        );

    \I__7119\ : InMux
    port map (
            O => \N__30641\,
            I => \N__30620\
        );

    \I__7118\ : Span4Mux_s2_v
    port map (
            O => \N__30636\,
            I => \N__30617\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30614\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__30626\,
            I => \N__30611\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__30623\,
            I => \N__30608\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__30620\,
            I => \N__30605\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__30617\,
            I => \N__30602\
        );

    \I__7112\ : Span4Mux_s2_v
    port map (
            O => \N__30614\,
            I => \N__30599\
        );

    \I__7111\ : Span4Mux_s2_v
    port map (
            O => \N__30611\,
            I => \N__30592\
        );

    \I__7110\ : Span4Mux_h
    port map (
            O => \N__30608\,
            I => \N__30592\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__30605\,
            I => \N__30592\
        );

    \I__7108\ : Span4Mux_h
    port map (
            O => \N__30602\,
            I => \N__30589\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__30599\,
            I => \N__30584\
        );

    \I__7106\ : Span4Mux_v
    port map (
            O => \N__30592\,
            I => \N__30584\
        );

    \I__7105\ : Odrv4
    port map (
            O => \N__30589\,
            I => \r_SM_Main_2_adj_1734\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__30584\,
            I => \r_SM_Main_2_adj_1734\
        );

    \I__7103\ : CascadeMux
    port map (
            O => \N__30579\,
            I => \N__30576\
        );

    \I__7102\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30573\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__7100\ : Span4Mux_s2_v
    port map (
            O => \N__30570\,
            I => \N__30564\
        );

    \I__7099\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30558\
        );

    \I__7098\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30558\
        );

    \I__7097\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30555\
        );

    \I__7096\ : Span4Mux_h
    port map (
            O => \N__30564\,
            I => \N__30552\
        );

    \I__7095\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30549\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__30558\,
            I => \N__30544\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__30555\,
            I => \N__30544\
        );

    \I__7092\ : Odrv4
    port map (
            O => \N__30552\,
            I => \r_SM_Main_2_N_1537_2\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__30549\,
            I => \r_SM_Main_2_N_1537_2\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__30544\,
            I => \r_SM_Main_2_N_1537_2\
        );

    \I__7089\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__30534\,
            I => n9245
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__30531\,
            I => \N__30527\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__30530\,
            I => \N__30524\
        );

    \I__7085\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30519\
        );

    \I__7084\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30516\
        );

    \I__7083\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30511\
        );

    \I__7082\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30511\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__30519\,
            I => \r_Clock_Count_0_adj_1730\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__30516\,
            I => \r_Clock_Count_0_adj_1730\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__30511\,
            I => \r_Clock_Count_0_adj_1730\
        );

    \I__7078\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30501\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__30501\,
            I => n226
        );

    \I__7076\ : InMux
    port map (
            O => \N__30498\,
            I => \bfn_11_31_0_\
        );

    \I__7075\ : CascadeMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__7074\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30485\
        );

    \I__7073\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30482\
        );

    \I__7072\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30479\
        );

    \I__7071\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30474\
        );

    \I__7070\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30474\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__30485\,
            I => \r_Clock_Count_1\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__30482\,
            I => \r_Clock_Count_1\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__30479\,
            I => \r_Clock_Count_1\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__30474\,
            I => \r_Clock_Count_1\
        );

    \I__7065\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30462\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__7063\ : Odrv4
    port map (
            O => \N__30459\,
            I => n225
        );

    \I__7062\ : InMux
    port map (
            O => \N__30456\,
            I => \c0.rx.n8098\
        );

    \I__7061\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30446\
        );

    \I__7060\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30443\
        );

    \I__7059\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30440\
        );

    \I__7058\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30435\
        );

    \I__7057\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30435\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__30446\,
            I => \r_Clock_Count_2\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__30443\,
            I => \r_Clock_Count_2\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__30440\,
            I => \r_Clock_Count_2\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__30435\,
            I => \r_Clock_Count_2\
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__7051\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30420\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__30420\,
            I => n224
        );

    \I__7049\ : InMux
    port map (
            O => \N__30417\,
            I => \c0.rx.n8099\
        );

    \I__7048\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30407\
        );

    \I__7047\ : InMux
    port map (
            O => \N__30413\,
            I => \N__30404\
        );

    \I__7046\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30401\
        );

    \I__7045\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30396\
        );

    \I__7044\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30396\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__30407\,
            I => \r_Clock_Count_3\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__30404\,
            I => \r_Clock_Count_3\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__30401\,
            I => \r_Clock_Count_3\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__30396\,
            I => \r_Clock_Count_3\
        );

    \I__7039\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30384\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__30384\,
            I => n223
        );

    \I__7037\ : InMux
    port map (
            O => \N__30381\,
            I => \c0.rx.n8100\
        );

    \I__7036\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30375\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__30375\,
            I => n7
        );

    \I__7034\ : InMux
    port map (
            O => \N__30372\,
            I => n8148
        );

    \I__7033\ : InMux
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__30366\,
            I => n6
        );

    \I__7031\ : InMux
    port map (
            O => \N__30363\,
            I => n8149
        );

    \I__7030\ : CascadeMux
    port map (
            O => \N__30360\,
            I => \N__30356\
        );

    \I__7029\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30351\
        );

    \I__7028\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30351\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__7026\ : Span4Mux_h
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__7025\ : Sp12to4
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__7024\ : Span12Mux_v
    port map (
            O => \N__30342\,
            I => \N__30338\
        );

    \I__7023\ : InMux
    port map (
            O => \N__30341\,
            I => \N__30335\
        );

    \I__7022\ : Odrv12
    port map (
            O => \N__30338\,
            I => blink_counter_21
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__30335\,
            I => blink_counter_21
        );

    \I__7020\ : InMux
    port map (
            O => \N__30330\,
            I => n8150
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__7018\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30318\
        );

    \I__7017\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30318\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__7015\ : Span4Mux_v
    port map (
            O => \N__30315\,
            I => \N__30312\
        );

    \I__7014\ : Span4Mux_h
    port map (
            O => \N__30312\,
            I => \N__30308\
        );

    \I__7013\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30305\
        );

    \I__7012\ : Odrv4
    port map (
            O => \N__30308\,
            I => blink_counter_22
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__30305\,
            I => blink_counter_22
        );

    \I__7010\ : InMux
    port map (
            O => \N__30300\,
            I => n8151
        );

    \I__7009\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30291\
        );

    \I__7008\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30291\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__30288\,
            I => \N__30285\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__30285\,
            I => \N__30281\
        );

    \I__7004\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30278\
        );

    \I__7003\ : Odrv4
    port map (
            O => \N__30281\,
            I => blink_counter_23
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__30278\,
            I => blink_counter_23
        );

    \I__7001\ : InMux
    port map (
            O => \N__30273\,
            I => n8152
        );

    \I__7000\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30264\
        );

    \I__6999\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30264\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__6997\ : Span12Mux_s10_h
    port map (
            O => \N__30261\,
            I => \N__30257\
        );

    \I__6996\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30254\
        );

    \I__6995\ : Odrv12
    port map (
            O => \N__30257\,
            I => blink_counter_24
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__30254\,
            I => blink_counter_24
        );

    \I__6993\ : InMux
    port map (
            O => \N__30249\,
            I => \bfn_11_30_0_\
        );

    \I__6992\ : InMux
    port map (
            O => \N__30246\,
            I => n8154
        );

    \I__6991\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__6989\ : Span12Mux_v
    port map (
            O => \N__30237\,
            I => \N__30233\
        );

    \I__6988\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30230\
        );

    \I__6987\ : Odrv12
    port map (
            O => \N__30233\,
            I => blink_counter_25
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__30230\,
            I => blink_counter_25
        );

    \I__6985\ : InMux
    port map (
            O => \N__30225\,
            I => \N__30222\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__30222\,
            I => n15
        );

    \I__6983\ : InMux
    port map (
            O => \N__30219\,
            I => n8140
        );

    \I__6982\ : InMux
    port map (
            O => \N__30216\,
            I => \N__30213\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__30213\,
            I => n14
        );

    \I__6980\ : InMux
    port map (
            O => \N__30210\,
            I => n8141
        );

    \I__6979\ : InMux
    port map (
            O => \N__30207\,
            I => \N__30204\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__30204\,
            I => n13
        );

    \I__6977\ : InMux
    port map (
            O => \N__30201\,
            I => n8142
        );

    \I__6976\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__30195\,
            I => n12
        );

    \I__6974\ : InMux
    port map (
            O => \N__30192\,
            I => n8143
        );

    \I__6973\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30186\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__30186\,
            I => n11
        );

    \I__6971\ : InMux
    port map (
            O => \N__30183\,
            I => n8144
        );

    \I__6970\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__30177\,
            I => n10
        );

    \I__6968\ : InMux
    port map (
            O => \N__30174\,
            I => \bfn_11_29_0_\
        );

    \I__6967\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__30168\,
            I => n9
        );

    \I__6965\ : InMux
    port map (
            O => \N__30165\,
            I => n8146
        );

    \I__6964\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30159\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__30159\,
            I => n8
        );

    \I__6962\ : InMux
    port map (
            O => \N__30156\,
            I => n8147
        );

    \I__6961\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__30150\,
            I => n24
        );

    \I__6959\ : InMux
    port map (
            O => \N__30147\,
            I => n8131
        );

    \I__6958\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__30141\,
            I => n23
        );

    \I__6956\ : InMux
    port map (
            O => \N__30138\,
            I => n8132
        );

    \I__6955\ : InMux
    port map (
            O => \N__30135\,
            I => \N__30132\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__30132\,
            I => n22
        );

    \I__6953\ : InMux
    port map (
            O => \N__30129\,
            I => n8133
        );

    \I__6952\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__30123\,
            I => n21
        );

    \I__6950\ : InMux
    port map (
            O => \N__30120\,
            I => n8134
        );

    \I__6949\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__30114\,
            I => n20
        );

    \I__6947\ : InMux
    port map (
            O => \N__30111\,
            I => n8135
        );

    \I__6946\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30105\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__30105\,
            I => n19
        );

    \I__6944\ : InMux
    port map (
            O => \N__30102\,
            I => n8136
        );

    \I__6943\ : InMux
    port map (
            O => \N__30099\,
            I => \N__30096\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__30096\,
            I => n18
        );

    \I__6941\ : InMux
    port map (
            O => \N__30093\,
            I => \bfn_11_28_0_\
        );

    \I__6940\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30087\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__30087\,
            I => n17
        );

    \I__6938\ : InMux
    port map (
            O => \N__30084\,
            I => n8138
        );

    \I__6937\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30078\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__30078\,
            I => n16
        );

    \I__6935\ : InMux
    port map (
            O => \N__30075\,
            I => n8139
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__30072\,
            I => \N__30069\
        );

    \I__6933\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30066\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30063\
        );

    \I__6931\ : Odrv4
    port map (
            O => \N__30063\,
            I => \c0.n22_adj_1661\
        );

    \I__6930\ : InMux
    port map (
            O => \N__30060\,
            I => \N__30057\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__30057\,
            I => \c0.n9731\
        );

    \I__6928\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30051\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__30051\,
            I => \N__30048\
        );

    \I__6926\ : Span4Mux_h
    port map (
            O => \N__30048\,
            I => \N__30045\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__30045\,
            I => \N__30042\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__30042\,
            I => \N__30039\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__30039\,
            I => \c0.tx2.r_Tx_Data_0\
        );

    \I__6922\ : CascadeMux
    port map (
            O => \N__30036\,
            I => \N__30025\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30015\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__30034\,
            I => \N__30012\
        );

    \I__6919\ : CascadeMux
    port map (
            O => \N__30033\,
            I => \N__30009\
        );

    \I__6918\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30002\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__30031\,
            I => \N__29999\
        );

    \I__6916\ : CascadeMux
    port map (
            O => \N__30030\,
            I => \N__29996\
        );

    \I__6915\ : CascadeMux
    port map (
            O => \N__30029\,
            I => \N__29961\
        );

    \I__6914\ : CascadeMux
    port map (
            O => \N__30028\,
            I => \N__29958\
        );

    \I__6913\ : InMux
    port map (
            O => \N__30025\,
            I => \N__29942\
        );

    \I__6912\ : InMux
    port map (
            O => \N__30024\,
            I => \N__29942\
        );

    \I__6911\ : InMux
    port map (
            O => \N__30023\,
            I => \N__29942\
        );

    \I__6910\ : InMux
    port map (
            O => \N__30022\,
            I => \N__29942\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30021\,
            I => \N__29942\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__30020\,
            I => \N__29939\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__30019\,
            I => \N__29936\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__30018\,
            I => \N__29933\
        );

    \I__6905\ : InMux
    port map (
            O => \N__30015\,
            I => \N__29908\
        );

    \I__6904\ : InMux
    port map (
            O => \N__30012\,
            I => \N__29908\
        );

    \I__6903\ : InMux
    port map (
            O => \N__30009\,
            I => \N__29908\
        );

    \I__6902\ : InMux
    port map (
            O => \N__30008\,
            I => \N__29908\
        );

    \I__6901\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29908\
        );

    \I__6900\ : InMux
    port map (
            O => \N__30006\,
            I => \N__29908\
        );

    \I__6899\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29908\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29905\
        );

    \I__6897\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29894\
        );

    \I__6896\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29894\
        );

    \I__6895\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29894\
        );

    \I__6894\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29894\
        );

    \I__6893\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29894\
        );

    \I__6892\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29887\
        );

    \I__6891\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29887\
        );

    \I__6890\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29887\
        );

    \I__6889\ : CascadeMux
    port map (
            O => \N__29989\,
            I => \N__29879\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__29988\,
            I => \N__29876\
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__29987\,
            I => \N__29867\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__29986\,
            I => \N__29863\
        );

    \I__6885\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29846\
        );

    \I__6884\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29846\
        );

    \I__6883\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29846\
        );

    \I__6882\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29846\
        );

    \I__6881\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29846\
        );

    \I__6880\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29846\
        );

    \I__6879\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29830\
        );

    \I__6878\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29830\
        );

    \I__6877\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29830\
        );

    \I__6876\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29825\
        );

    \I__6875\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29825\
        );

    \I__6874\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29816\
        );

    \I__6873\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29816\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29816\
        );

    \I__6871\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29816\
        );

    \I__6870\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29805\
        );

    \I__6869\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29805\
        );

    \I__6868\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29805\
        );

    \I__6867\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29805\
        );

    \I__6866\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29805\
        );

    \I__6865\ : CascadeMux
    port map (
            O => \N__29965\,
            I => \N__29797\
        );

    \I__6864\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29782\
        );

    \I__6863\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29782\
        );

    \I__6862\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29782\
        );

    \I__6861\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29782\
        );

    \I__6860\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29782\
        );

    \I__6859\ : CascadeMux
    port map (
            O => \N__29955\,
            I => \N__29771\
        );

    \I__6858\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29763\
        );

    \I__6857\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29760\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29756\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29743\
        );

    \I__6854\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29743\
        );

    \I__6853\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29743\
        );

    \I__6852\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29743\
        );

    \I__6851\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29743\
        );

    \I__6850\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29743\
        );

    \I__6849\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29740\
        );

    \I__6848\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29735\
        );

    \I__6847\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29735\
        );

    \I__6846\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29730\
        );

    \I__6845\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29730\
        );

    \I__6844\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29727\
        );

    \I__6843\ : InMux
    port map (
            O => \N__29923\,
            I => \N__29724\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__29908\,
            I => \N__29721\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__29905\,
            I => \N__29714\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29714\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__29887\,
            I => \N__29714\
        );

    \I__6838\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29705\
        );

    \I__6837\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29705\
        );

    \I__6836\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29705\
        );

    \I__6835\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29702\
        );

    \I__6834\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29694\
        );

    \I__6833\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29685\
        );

    \I__6832\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29685\
        );

    \I__6831\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29685\
        );

    \I__6830\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29685\
        );

    \I__6829\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29676\
        );

    \I__6828\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29676\
        );

    \I__6827\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29676\
        );

    \I__6826\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29676\
        );

    \I__6825\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29671\
        );

    \I__6824\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29671\
        );

    \I__6823\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29660\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29660\
        );

    \I__6821\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29660\
        );

    \I__6820\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29660\
        );

    \I__6819\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29660\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__29846\,
            I => \N__29657\
        );

    \I__6817\ : CascadeMux
    port map (
            O => \N__29845\,
            I => \N__29639\
        );

    \I__6816\ : CascadeMux
    port map (
            O => \N__29844\,
            I => \N__29636\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__29843\,
            I => \N__29628\
        );

    \I__6814\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29620\
        );

    \I__6813\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29617\
        );

    \I__6812\ : InMux
    port map (
            O => \N__29840\,
            I => \N__29611\
        );

    \I__6811\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29604\
        );

    \I__6810\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29604\
        );

    \I__6809\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29604\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__29830\,
            I => \N__29599\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29599\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__29816\,
            I => \N__29594\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__29805\,
            I => \N__29594\
        );

    \I__6804\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29587\
        );

    \I__6803\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29587\
        );

    \I__6802\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29587\
        );

    \I__6801\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29572\
        );

    \I__6800\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29572\
        );

    \I__6799\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29572\
        );

    \I__6798\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29572\
        );

    \I__6797\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29572\
        );

    \I__6796\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29572\
        );

    \I__6795\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29572\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__29782\,
            I => \N__29567\
        );

    \I__6793\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29560\
        );

    \I__6792\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29560\
        );

    \I__6791\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29560\
        );

    \I__6790\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29551\
        );

    \I__6789\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29551\
        );

    \I__6788\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29551\
        );

    \I__6787\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29551\
        );

    \I__6786\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29536\
        );

    \I__6785\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29536\
        );

    \I__6784\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29536\
        );

    \I__6783\ : InMux
    port map (
            O => \N__29769\,
            I => \N__29536\
        );

    \I__6782\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29536\
        );

    \I__6781\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29536\
        );

    \I__6780\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29536\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__29763\,
            I => \N__29531\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__29760\,
            I => \N__29531\
        );

    \I__6777\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29528\
        );

    \I__6776\ : Span4Mux_v
    port map (
            O => \N__29756\,
            I => \N__29521\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__29743\,
            I => \N__29521\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__29740\,
            I => \N__29521\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__29735\,
            I => \N__29508\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29508\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__29727\,
            I => \N__29508\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__29724\,
            I => \N__29508\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__29721\,
            I => \N__29508\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__29714\,
            I => \N__29508\
        );

    \I__6767\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29503\
        );

    \I__6766\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29503\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29498\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__29702\,
            I => \N__29498\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__29701\,
            I => \N__29494\
        );

    \I__6762\ : CascadeMux
    port map (
            O => \N__29700\,
            I => \N__29489\
        );

    \I__6761\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29482\
        );

    \I__6760\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29477\
        );

    \I__6759\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29477\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__29694\,
            I => \N__29472\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29472\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__29676\,
            I => \N__29467\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29467\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29464\
        );

    \I__6753\ : Span4Mux_v
    port map (
            O => \N__29657\,
            I => \N__29461\
        );

    \I__6752\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29452\
        );

    \I__6751\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29452\
        );

    \I__6750\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29452\
        );

    \I__6749\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29452\
        );

    \I__6748\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29447\
        );

    \I__6747\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29447\
        );

    \I__6746\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29444\
        );

    \I__6745\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29437\
        );

    \I__6744\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29437\
        );

    \I__6743\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29437\
        );

    \I__6742\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29428\
        );

    \I__6741\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29428\
        );

    \I__6740\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29428\
        );

    \I__6739\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29428\
        );

    \I__6738\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29425\
        );

    \I__6737\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29414\
        );

    \I__6736\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29414\
        );

    \I__6735\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29414\
        );

    \I__6734\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29414\
        );

    \I__6733\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29414\
        );

    \I__6732\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29409\
        );

    \I__6731\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29409\
        );

    \I__6730\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29400\
        );

    \I__6729\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29400\
        );

    \I__6728\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29400\
        );

    \I__6727\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29400\
        );

    \I__6726\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29397\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__29623\,
            I => \N__29390\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__29620\,
            I => \N__29384\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__29617\,
            I => \N__29381\
        );

    \I__6722\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29375\
        );

    \I__6721\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29375\
        );

    \I__6720\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29372\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29359\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__29604\,
            I => \N__29359\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__29599\,
            I => \N__29359\
        );

    \I__6716\ : Span4Mux_v
    port map (
            O => \N__29594\,
            I => \N__29359\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__29587\,
            I => \N__29359\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__29572\,
            I => \N__29359\
        );

    \I__6713\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29353\
        );

    \I__6712\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29353\
        );

    \I__6711\ : Span4Mux_v
    port map (
            O => \N__29567\,
            I => \N__29332\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__29560\,
            I => \N__29332\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__29551\,
            I => \N__29332\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__29536\,
            I => \N__29332\
        );

    \I__6707\ : Span4Mux_v
    port map (
            O => \N__29531\,
            I => \N__29332\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__29528\,
            I => \N__29332\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__29521\,
            I => \N__29332\
        );

    \I__6704\ : Span4Mux_h
    port map (
            O => \N__29508\,
            I => \N__29332\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29332\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__29498\,
            I => \N__29332\
        );

    \I__6701\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29325\
        );

    \I__6700\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29325\
        );

    \I__6699\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29325\
        );

    \I__6698\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29322\
        );

    \I__6697\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29311\
        );

    \I__6696\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29311\
        );

    \I__6695\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29311\
        );

    \I__6694\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29311\
        );

    \I__6693\ : InMux
    port map (
            O => \N__29485\,
            I => \N__29311\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__29482\,
            I => \N__29288\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__29477\,
            I => \N__29288\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__29472\,
            I => \N__29288\
        );

    \I__6689\ : Span4Mux_v
    port map (
            O => \N__29467\,
            I => \N__29288\
        );

    \I__6688\ : Span4Mux_v
    port map (
            O => \N__29464\,
            I => \N__29288\
        );

    \I__6687\ : Span4Mux_h
    port map (
            O => \N__29461\,
            I => \N__29288\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__29452\,
            I => \N__29288\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29288\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__29444\,
            I => \N__29288\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29288\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__29428\,
            I => \N__29288\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__29425\,
            I => \N__29279\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__29414\,
            I => \N__29279\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29279\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__29400\,
            I => \N__29279\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__29397\,
            I => \N__29276\
        );

    \I__6676\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29273\
        );

    \I__6675\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29270\
        );

    \I__6674\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29267\
        );

    \I__6673\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29258\
        );

    \I__6672\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29258\
        );

    \I__6671\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29258\
        );

    \I__6670\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29258\
        );

    \I__6669\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29255\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29251\
        );

    \I__6667\ : Span4Mux_v
    port map (
            O => \N__29381\,
            I => \N__29248\
        );

    \I__6666\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29245\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__29375\,
            I => \N__29238\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__29372\,
            I => \N__29238\
        );

    \I__6663\ : Span4Mux_h
    port map (
            O => \N__29359\,
            I => \N__29238\
        );

    \I__6662\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29235\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__29353\,
            I => \N__29230\
        );

    \I__6660\ : Sp12to4
    port map (
            O => \N__29332\,
            I => \N__29230\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__29325\,
            I => \N__29219\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__29322\,
            I => \N__29219\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__29311\,
            I => \N__29219\
        );

    \I__6656\ : Span4Mux_h
    port map (
            O => \N__29288\,
            I => \N__29219\
        );

    \I__6655\ : Span4Mux_s2_h
    port map (
            O => \N__29279\,
            I => \N__29219\
        );

    \I__6654\ : Span4Mux_v
    port map (
            O => \N__29276\,
            I => \N__29216\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__29273\,
            I => \N__29213\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__29270\,
            I => \N__29206\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__29267\,
            I => \N__29206\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__29258\,
            I => \N__29206\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__29255\,
            I => \N__29203\
        );

    \I__6648\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29200\
        );

    \I__6647\ : Span4Mux_s0_v
    port map (
            O => \N__29251\,
            I => \N__29195\
        );

    \I__6646\ : Span4Mux_v
    port map (
            O => \N__29248\,
            I => \N__29195\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29184\
        );

    \I__6644\ : Sp12to4
    port map (
            O => \N__29238\,
            I => \N__29184\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29184\
        );

    \I__6642\ : Span12Mux_s2_h
    port map (
            O => \N__29230\,
            I => \N__29184\
        );

    \I__6641\ : Sp12to4
    port map (
            O => \N__29219\,
            I => \N__29184\
        );

    \I__6640\ : Span4Mux_v
    port map (
            O => \N__29216\,
            I => \N__29179\
        );

    \I__6639\ : Span4Mux_s3_h
    port map (
            O => \N__29213\,
            I => \N__29179\
        );

    \I__6638\ : Span12Mux_v
    port map (
            O => \N__29206\,
            I => \N__29176\
        );

    \I__6637\ : Span12Mux_v
    port map (
            O => \N__29203\,
            I => \N__29173\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29166\
        );

    \I__6635\ : Sp12to4
    port map (
            O => \N__29195\,
            I => \N__29166\
        );

    \I__6634\ : Span12Mux_v
    port map (
            O => \N__29184\,
            I => \N__29166\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__29179\,
            I => rx_data_ready
        );

    \I__6632\ : Odrv12
    port map (
            O => \N__29176\,
            I => rx_data_ready
        );

    \I__6631\ : Odrv12
    port map (
            O => \N__29173\,
            I => rx_data_ready
        );

    \I__6630\ : Odrv12
    port map (
            O => \N__29166\,
            I => rx_data_ready
        );

    \I__6629\ : InMux
    port map (
            O => \N__29157\,
            I => \N__29154\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__6627\ : Span4Mux_h
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__6626\ : Span4Mux_v
    port map (
            O => \N__29148\,
            I => \N__29144\
        );

    \I__6625\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29141\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__29144\,
            I => data_in_19_0
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__29141\,
            I => data_in_19_0
        );

    \I__6622\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__6620\ : Span4Mux_h
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__6619\ : Span4Mux_h
    port map (
            O => \N__29127\,
            I => \N__29123\
        );

    \I__6618\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29120\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__29123\,
            I => data_in_18_0
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__29120\,
            I => data_in_18_0
        );

    \I__6615\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29112\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__29112\,
            I => \N__29109\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__29109\,
            I => \N__29104\
        );

    \I__6612\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29101\
        );

    \I__6611\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29098\
        );

    \I__6610\ : Span4Mux_h
    port map (
            O => \N__29104\,
            I => \N__29093\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__29101\,
            I => \N__29088\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29088\
        );

    \I__6607\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29085\
        );

    \I__6606\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29082\
        );

    \I__6605\ : Odrv4
    port map (
            O => \N__29093\,
            I => rand_data_12
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__29088\,
            I => rand_data_12
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__29085\,
            I => rand_data_12
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__29082\,
            I => rand_data_12
        );

    \I__6601\ : CEMux
    port map (
            O => \N__29073\,
            I => \N__29059\
        );

    \I__6600\ : CEMux
    port map (
            O => \N__29072\,
            I => \N__29049\
        );

    \I__6599\ : CascadeMux
    port map (
            O => \N__29071\,
            I => \N__29043\
        );

    \I__6598\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29039\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__29069\,
            I => \N__29036\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__29068\,
            I => \N__29033\
        );

    \I__6595\ : CEMux
    port map (
            O => \N__29067\,
            I => \N__29027\
        );

    \I__6594\ : CEMux
    port map (
            O => \N__29066\,
            I => \N__29022\
        );

    \I__6593\ : CascadeMux
    port map (
            O => \N__29065\,
            I => \N__29016\
        );

    \I__6592\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29000\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__29063\,
            I => \N__28993\
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__29062\,
            I => \N__28987\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__29059\,
            I => \N__28981\
        );

    \I__6588\ : InMux
    port map (
            O => \N__29058\,
            I => \N__28976\
        );

    \I__6587\ : InMux
    port map (
            O => \N__29057\,
            I => \N__28976\
        );

    \I__6586\ : InMux
    port map (
            O => \N__29056\,
            I => \N__28973\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__29055\,
            I => \N__28969\
        );

    \I__6584\ : CascadeMux
    port map (
            O => \N__29054\,
            I => \N__28963\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__29053\,
            I => \N__28958\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__29052\,
            I => \N__28954\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__28950\
        );

    \I__6580\ : CEMux
    port map (
            O => \N__29048\,
            I => \N__28947\
        );

    \I__6579\ : CEMux
    port map (
            O => \N__29047\,
            I => \N__28944\
        );

    \I__6578\ : InMux
    port map (
            O => \N__29046\,
            I => \N__28937\
        );

    \I__6577\ : InMux
    port map (
            O => \N__29043\,
            I => \N__28937\
        );

    \I__6576\ : InMux
    port map (
            O => \N__29042\,
            I => \N__28937\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__29039\,
            I => \N__28934\
        );

    \I__6574\ : InMux
    port map (
            O => \N__29036\,
            I => \N__28925\
        );

    \I__6573\ : InMux
    port map (
            O => \N__29033\,
            I => \N__28925\
        );

    \I__6572\ : InMux
    port map (
            O => \N__29032\,
            I => \N__28925\
        );

    \I__6571\ : InMux
    port map (
            O => \N__29031\,
            I => \N__28925\
        );

    \I__6570\ : CEMux
    port map (
            O => \N__29030\,
            I => \N__28921\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__29027\,
            I => \N__28918\
        );

    \I__6568\ : CEMux
    port map (
            O => \N__29026\,
            I => \N__28915\
        );

    \I__6567\ : CEMux
    port map (
            O => \N__29025\,
            I => \N__28912\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__28909\
        );

    \I__6565\ : CEMux
    port map (
            O => \N__29021\,
            I => \N__28906\
        );

    \I__6564\ : InMux
    port map (
            O => \N__29020\,
            I => \N__28897\
        );

    \I__6563\ : InMux
    port map (
            O => \N__29019\,
            I => \N__28897\
        );

    \I__6562\ : InMux
    port map (
            O => \N__29016\,
            I => \N__28897\
        );

    \I__6561\ : InMux
    port map (
            O => \N__29015\,
            I => \N__28897\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__29014\,
            I => \N__28893\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__29013\,
            I => \N__28889\
        );

    \I__6558\ : InMux
    port map (
            O => \N__29012\,
            I => \N__28886\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__29011\,
            I => \N__28882\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__29010\,
            I => \N__28878\
        );

    \I__6555\ : CEMux
    port map (
            O => \N__29009\,
            I => \N__28874\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__29008\,
            I => \N__28870\
        );

    \I__6553\ : CascadeMux
    port map (
            O => \N__29007\,
            I => \N__28864\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__29006\,
            I => \N__28860\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__29005\,
            I => \N__28857\
        );

    \I__6550\ : CEMux
    port map (
            O => \N__29004\,
            I => \N__28845\
        );

    \I__6549\ : CEMux
    port map (
            O => \N__29003\,
            I => \N__28842\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__29000\,
            I => \N__28839\
        );

    \I__6547\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28834\
        );

    \I__6546\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28834\
        );

    \I__6545\ : CEMux
    port map (
            O => \N__28997\,
            I => \N__28831\
        );

    \I__6544\ : CEMux
    port map (
            O => \N__28996\,
            I => \N__28828\
        );

    \I__6543\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28823\
        );

    \I__6542\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28823\
        );

    \I__6541\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28814\
        );

    \I__6540\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28814\
        );

    \I__6539\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28814\
        );

    \I__6538\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28814\
        );

    \I__6537\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28809\
        );

    \I__6536\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28809\
        );

    \I__6535\ : Span4Mux_h
    port map (
            O => \N__28981\,
            I => \N__28802\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__28976\,
            I => \N__28802\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__28973\,
            I => \N__28802\
        );

    \I__6532\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28799\
        );

    \I__6531\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28794\
        );

    \I__6530\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28794\
        );

    \I__6529\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28791\
        );

    \I__6528\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28784\
        );

    \I__6527\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28784\
        );

    \I__6526\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28784\
        );

    \I__6525\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28773\
        );

    \I__6524\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28773\
        );

    \I__6523\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28773\
        );

    \I__6522\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28773\
        );

    \I__6521\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28773\
        );

    \I__6520\ : Span4Mux_s1_v
    port map (
            O => \N__28950\,
            I => \N__28769\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__28947\,
            I => \N__28764\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28764\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__28937\,
            I => \N__28761\
        );

    \I__6516\ : Span4Mux_v
    port map (
            O => \N__28934\,
            I => \N__28756\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__28925\,
            I => \N__28756\
        );

    \I__6514\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28753\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__28921\,
            I => \N__28739\
        );

    \I__6512\ : Span4Mux_s1_h
    port map (
            O => \N__28918\,
            I => \N__28734\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__28915\,
            I => \N__28734\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__28912\,
            I => \N__28731\
        );

    \I__6509\ : Span4Mux_s1_h
    port map (
            O => \N__28909\,
            I => \N__28728\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__28906\,
            I => \N__28723\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__28897\,
            I => \N__28723\
        );

    \I__6506\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28714\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28714\
        );

    \I__6504\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28714\
        );

    \I__6503\ : InMux
    port map (
            O => \N__28889\,
            I => \N__28714\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28711\
        );

    \I__6501\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28700\
        );

    \I__6500\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28700\
        );

    \I__6499\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28700\
        );

    \I__6498\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28700\
        );

    \I__6497\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28700\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28697\
        );

    \I__6495\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28690\
        );

    \I__6494\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28690\
        );

    \I__6493\ : InMux
    port map (
            O => \N__28869\,
            I => \N__28690\
        );

    \I__6492\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28685\
        );

    \I__6491\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28685\
        );

    \I__6490\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28674\
        );

    \I__6489\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28674\
        );

    \I__6488\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28674\
        );

    \I__6487\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28674\
        );

    \I__6486\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28674\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__28855\,
            I => \N__28669\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__28854\,
            I => \N__28666\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__28853\,
            I => \N__28662\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__28852\,
            I => \N__28659\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__28851\,
            I => \N__28655\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__28850\,
            I => \N__28651\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__28849\,
            I => \N__28648\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__28848\,
            I => \N__28644\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__28845\,
            I => \N__28639\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__28842\,
            I => \N__28636\
        );

    \I__6475\ : Span4Mux_s3_h
    port map (
            O => \N__28839\,
            I => \N__28633\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28630\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__28831\,
            I => \N__28613\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28613\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28613\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28613\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28613\
        );

    \I__6468\ : Span4Mux_h
    port map (
            O => \N__28802\,
            I => \N__28613\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__28799\,
            I => \N__28613\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__28794\,
            I => \N__28613\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__28791\,
            I => \N__28606\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28606\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__28773\,
            I => \N__28606\
        );

    \I__6462\ : InMux
    port map (
            O => \N__28772\,
            I => \N__28603\
        );

    \I__6461\ : Span4Mux_v
    port map (
            O => \N__28769\,
            I => \N__28592\
        );

    \I__6460\ : Span4Mux_v
    port map (
            O => \N__28764\,
            I => \N__28592\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__28761\,
            I => \N__28592\
        );

    \I__6458\ : Span4Mux_h
    port map (
            O => \N__28756\,
            I => \N__28592\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__28753\,
            I => \N__28592\
        );

    \I__6456\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28589\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__28751\,
            I => \N__28586\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__28750\,
            I => \N__28582\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__28749\,
            I => \N__28579\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__28748\,
            I => \N__28574\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__28747\,
            I => \N__28571\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__28746\,
            I => \N__28568\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__28745\,
            I => \N__28564\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__28744\,
            I => \N__28560\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__28743\,
            I => \N__28554\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__28742\,
            I => \N__28551\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__28739\,
            I => \N__28547\
        );

    \I__6444\ : Span4Mux_h
    port map (
            O => \N__28734\,
            I => \N__28542\
        );

    \I__6443\ : Span4Mux_h
    port map (
            O => \N__28731\,
            I => \N__28542\
        );

    \I__6442\ : Span4Mux_h
    port map (
            O => \N__28728\,
            I => \N__28531\
        );

    \I__6441\ : Span4Mux_s3_v
    port map (
            O => \N__28723\,
            I => \N__28531\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__28714\,
            I => \N__28531\
        );

    \I__6439\ : Span4Mux_v
    port map (
            O => \N__28711\,
            I => \N__28531\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28531\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__28697\,
            I => \N__28526\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__28690\,
            I => \N__28526\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__28685\,
            I => \N__28521\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__28674\,
            I => \N__28521\
        );

    \I__6433\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28518\
        );

    \I__6432\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28503\
        );

    \I__6431\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28503\
        );

    \I__6430\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28503\
        );

    \I__6429\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28503\
        );

    \I__6428\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28503\
        );

    \I__6427\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28503\
        );

    \I__6426\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28503\
        );

    \I__6425\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28486\
        );

    \I__6424\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28486\
        );

    \I__6423\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28486\
        );

    \I__6422\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28486\
        );

    \I__6421\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28486\
        );

    \I__6420\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28486\
        );

    \I__6419\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28486\
        );

    \I__6418\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28486\
        );

    \I__6417\ : Span4Mux_s3_h
    port map (
            O => \N__28639\,
            I => \N__28471\
        );

    \I__6416\ : Span4Mux_s3_h
    port map (
            O => \N__28636\,
            I => \N__28471\
        );

    \I__6415\ : Span4Mux_v
    port map (
            O => \N__28633\,
            I => \N__28471\
        );

    \I__6414\ : Span4Mux_v
    port map (
            O => \N__28630\,
            I => \N__28471\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__28613\,
            I => \N__28471\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__28606\,
            I => \N__28471\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28471\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__28592\,
            I => \N__28466\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__28589\,
            I => \N__28466\
        );

    \I__6408\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28455\
        );

    \I__6407\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28455\
        );

    \I__6406\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28455\
        );

    \I__6405\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28455\
        );

    \I__6404\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28455\
        );

    \I__6403\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28440\
        );

    \I__6402\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28440\
        );

    \I__6401\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28440\
        );

    \I__6400\ : InMux
    port map (
            O => \N__28568\,
            I => \N__28440\
        );

    \I__6399\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28440\
        );

    \I__6398\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28440\
        );

    \I__6397\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28440\
        );

    \I__6396\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28425\
        );

    \I__6395\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28425\
        );

    \I__6394\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28425\
        );

    \I__6393\ : InMux
    port map (
            O => \N__28557\,
            I => \N__28425\
        );

    \I__6392\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28425\
        );

    \I__6391\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28425\
        );

    \I__6390\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28425\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__28547\,
            I => n4806
        );

    \I__6388\ : Odrv4
    port map (
            O => \N__28542\,
            I => n4806
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__28531\,
            I => n4806
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__28526\,
            I => n4806
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__28521\,
            I => n4806
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__28518\,
            I => n4806
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__28503\,
            I => n4806
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__28486\,
            I => n4806
        );

    \I__6381\ : Odrv4
    port map (
            O => \N__28471\,
            I => n4806
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__28466\,
            I => n4806
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__28455\,
            I => n4806
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__28440\,
            I => n4806
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__28425\,
            I => n4806
        );

    \I__6376\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28392\
        );

    \I__6375\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28389\
        );

    \I__6374\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28385\
        );

    \I__6373\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28382\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__28392\,
            I => \N__28378\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28375\
        );

    \I__6370\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28372\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28367\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__28382\,
            I => \N__28367\
        );

    \I__6367\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28364\
        );

    \I__6366\ : Span4Mux_h
    port map (
            O => \N__28378\,
            I => \N__28361\
        );

    \I__6365\ : Span12Mux_s6_v
    port map (
            O => \N__28375\,
            I => \N__28358\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__28372\,
            I => \N__28353\
        );

    \I__6363\ : Span4Mux_v
    port map (
            O => \N__28367\,
            I => \N__28353\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__28364\,
            I => data_in_field_88
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__28361\,
            I => data_in_field_88
        );

    \I__6360\ : Odrv12
    port map (
            O => \N__28358\,
            I => data_in_field_88
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__28353\,
            I => data_in_field_88
        );

    \I__6358\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28340\
        );

    \I__6357\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28337\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28331\
        );

    \I__6354\ : Span12Mux_s10_h
    port map (
            O => \N__28334\,
            I => \N__28328\
        );

    \I__6353\ : Span4Mux_h
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__6352\ : Odrv12
    port map (
            O => \N__28328\,
            I => \c0.n4292\
        );

    \I__6351\ : Odrv4
    port map (
            O => \N__28325\,
            I => \c0.n4292\
        );

    \I__6350\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28316\
        );

    \I__6349\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28313\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__28316\,
            I => \N__28310\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__28313\,
            I => \c0.n8957\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__28310\,
            I => \c0.n8957\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__28305\,
            I => \N__28302\
        );

    \I__6344\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28296\
        );

    \I__6343\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28293\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__28300\,
            I => \N__28289\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__28299\,
            I => \N__28286\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28283\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28280\
        );

    \I__6338\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28277\
        );

    \I__6337\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28274\
        );

    \I__6336\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28271\
        );

    \I__6335\ : Span4Mux_s3_h
    port map (
            O => \N__28283\,
            I => \N__28268\
        );

    \I__6334\ : Span12Mux_h
    port map (
            O => \N__28280\,
            I => \N__28265\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__28277\,
            I => \N__28262\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28259\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__28271\,
            I => \c0.data_in_field_27\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__28268\,
            I => \c0.data_in_field_27\
        );

    \I__6329\ : Odrv12
    port map (
            O => \N__28265\,
            I => \c0.data_in_field_27\
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__28262\,
            I => \c0.data_in_field_27\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__28259\,
            I => \c0.data_in_field_27\
        );

    \I__6326\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28241\
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__28244\,
            I => \N__28237\
        );

    \I__6323\ : Span4Mux_v
    port map (
            O => \N__28241\,
            I => \N__28234\
        );

    \I__6322\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28231\
        );

    \I__6321\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28226\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__28234\,
            I => \N__28223\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28220\
        );

    \I__6318\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28215\
        );

    \I__6317\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28215\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__28226\,
            I => \c0.data_in_field_25\
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__28223\,
            I => \c0.data_in_field_25\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__28220\,
            I => \c0.data_in_field_25\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__28215\,
            I => \c0.data_in_field_25\
        );

    \I__6312\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28203\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__28203\,
            I => \N__28200\
        );

    \I__6310\ : Sp12to4
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__6309\ : Span12Mux_s8_h
    port map (
            O => \N__28197\,
            I => \N__28194\
        );

    \I__6308\ : Odrv12
    port map (
            O => \N__28194\,
            I => \c0.n8871\
        );

    \I__6307\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28188\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__28188\,
            I => n26
        );

    \I__6305\ : InMux
    port map (
            O => \N__28185\,
            I => \bfn_11_27_0_\
        );

    \I__6304\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28179\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__28179\,
            I => n25_adj_1722
        );

    \I__6302\ : InMux
    port map (
            O => \N__28176\,
            I => n8130
        );

    \I__6301\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__28170\,
            I => n1
        );

    \I__6299\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28160\
        );

    \I__6298\ : CascadeMux
    port map (
            O => \N__28166\,
            I => \N__28153\
        );

    \I__6297\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28146\
        );

    \I__6296\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28146\
        );

    \I__6295\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28143\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__28160\,
            I => \N__28140\
        );

    \I__6293\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28133\
        );

    \I__6292\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28133\
        );

    \I__6291\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28133\
        );

    \I__6290\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28124\
        );

    \I__6289\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28124\
        );

    \I__6288\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28124\
        );

    \I__6287\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28124\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__28146\,
            I => \N__28121\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__28143\,
            I => \N__28118\
        );

    \I__6284\ : Sp12to4
    port map (
            O => \N__28140\,
            I => \N__28111\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28111\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__28124\,
            I => \N__28111\
        );

    \I__6281\ : Span4Mux_h
    port map (
            O => \N__28121\,
            I => \N__28108\
        );

    \I__6280\ : Span4Mux_h
    port map (
            O => \N__28118\,
            I => \N__28105\
        );

    \I__6279\ : Odrv12
    port map (
            O => \N__28111\,
            I => \r_Rx_Data\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__28108\,
            I => \r_Rx_Data\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__28105\,
            I => \r_Rx_Data\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28092\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28092\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__28092\,
            I => \c0.rx.r_SM_Main_2_N_1543_0\
        );

    \I__6273\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__28086\,
            I => n9300
        );

    \I__6271\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28080\,
            I => \N__28076\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__28079\,
            I => \N__28073\
        );

    \I__6268\ : Span4Mux_h
    port map (
            O => \N__28076\,
            I => \N__28070\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28066\
        );

    \I__6266\ : Span4Mux_h
    port map (
            O => \N__28070\,
            I => \N__28063\
        );

    \I__6265\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28060\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__28066\,
            I => \c0.data_in_field_24\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__28063\,
            I => \c0.data_in_field_24\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__28060\,
            I => \c0.data_in_field_24\
        );

    \I__6261\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__6259\ : Span4Mux_h
    port map (
            O => \N__28047\,
            I => \N__28044\
        );

    \I__6258\ : Span4Mux_h
    port map (
            O => \N__28044\,
            I => \N__28038\
        );

    \I__6257\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28033\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28033\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28030\
        );

    \I__6254\ : Odrv4
    port map (
            O => \N__28038\,
            I => \c0.data_in_field_16\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__28033\,
            I => \c0.data_in_field_16\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__28030\,
            I => \c0.data_in_field_16\
        );

    \I__6251\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__28020\,
            I => \N__28016\
        );

    \I__6249\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \N__28013\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__28016\,
            I => \N__28010\
        );

    \I__6247\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28006\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__28003\
        );

    \I__6245\ : InMux
    port map (
            O => \N__28009\,
            I => \N__28000\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__28006\,
            I => \c0.data_in_field_8\
        );

    \I__6243\ : Odrv4
    port map (
            O => \N__28003\,
            I => \c0.data_in_field_8\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__28000\,
            I => \c0.data_in_field_8\
        );

    \I__6241\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27990\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27986\
        );

    \I__6239\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27983\
        );

    \I__6238\ : Span4Mux_h
    port map (
            O => \N__27986\,
            I => \N__27979\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__27983\,
            I => \N__27976\
        );

    \I__6236\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27972\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__27979\,
            I => \N__27967\
        );

    \I__6234\ : Span4Mux_v
    port map (
            O => \N__27976\,
            I => \N__27967\
        );

    \I__6233\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27964\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__27972\,
            I => \c0.data_in_field_0\
        );

    \I__6231\ : Odrv4
    port map (
            O => \N__27967\,
            I => \c0.data_in_field_0\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__27964\,
            I => \c0.data_in_field_0\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__27957\,
            I => \c0.n9446_cascade_\
        );

    \I__6228\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27951\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__27951\,
            I => \N__27948\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__27948\,
            I => \N__27945\
        );

    \I__6225\ : Span4Mux_h
    port map (
            O => \N__27945\,
            I => \N__27942\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__27942\,
            I => \c0.n9228\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__27939\,
            I => \c0.n9449_cascade_\
        );

    \I__6222\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27933\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__27933\,
            I => \N__27927\
        );

    \I__6220\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27923\
        );

    \I__6219\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27920\
        );

    \I__6218\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27917\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__27927\,
            I => \N__27914\
        );

    \I__6216\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27911\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27906\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__27920\,
            I => \N__27906\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__27917\,
            I => data_in_field_80
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__27914\,
            I => data_in_field_80
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__27911\,
            I => data_in_field_80
        );

    \I__6210\ : Odrv12
    port map (
            O => \N__27906\,
            I => data_in_field_80
        );

    \I__6209\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27893\
        );

    \I__6208\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27890\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__27893\,
            I => \N__27887\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__27890\,
            I => \N__27883\
        );

    \I__6205\ : Span4Mux_h
    port map (
            O => \N__27887\,
            I => \N__27880\
        );

    \I__6204\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27876\
        );

    \I__6203\ : Span4Mux_h
    port map (
            O => \N__27883\,
            I => \N__27873\
        );

    \I__6202\ : Span4Mux_h
    port map (
            O => \N__27880\,
            I => \N__27870\
        );

    \I__6201\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27867\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__27876\,
            I => data_in_field_72
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__27873\,
            I => data_in_field_72
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__27870\,
            I => data_in_field_72
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__27867\,
            I => data_in_field_72
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__27858\,
            I => \c0.n9740_cascade_\
        );

    \I__6195\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27850\
        );

    \I__6194\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27847\
        );

    \I__6193\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27844\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__27850\,
            I => \N__27840\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__27847\,
            I => \N__27835\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__27844\,
            I => \N__27835\
        );

    \I__6189\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27832\
        );

    \I__6188\ : Span4Mux_h
    port map (
            O => \N__27840\,
            I => \N__27827\
        );

    \I__6187\ : Span4Mux_v
    port map (
            O => \N__27835\,
            I => \N__27827\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__27832\,
            I => data_in_field_64
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__27827\,
            I => data_in_field_64
        );

    \I__6184\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__6182\ : Span4Mux_v
    port map (
            O => \N__27816\,
            I => \N__27813\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__27810\,
            I => \c0.n9234\
        );

    \I__6179\ : CascadeMux
    port map (
            O => \N__27807\,
            I => \c0.n9231_cascade_\
        );

    \I__6178\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27801\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__27801\,
            I => \c0.n9728\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__27798\,
            I => \n6_adj_1751_cascade_\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__27795\,
            I => \n30_cascade_\
        );

    \I__6174\ : InMux
    port map (
            O => \N__27792\,
            I => \N__27788\
        );

    \I__6173\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27781\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__27788\,
            I => \N__27778\
        );

    \I__6171\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27775\
        );

    \I__6170\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27772\
        );

    \I__6169\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27767\
        );

    \I__6168\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27767\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27764\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__27778\,
            I => \N__27760\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__27775\,
            I => \N__27757\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__27772\,
            I => \N__27754\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27749\
        );

    \I__6162\ : Span4Mux_s2_h
    port map (
            O => \N__27764\,
            I => \N__27749\
        );

    \I__6161\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27746\
        );

    \I__6160\ : Span4Mux_h
    port map (
            O => \N__27760\,
            I => \N__27739\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__27757\,
            I => \N__27739\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__27754\,
            I => \N__27739\
        );

    \I__6157\ : Span4Mux_h
    port map (
            O => \N__27749\,
            I => \N__27736\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__27746\,
            I => data_in_field_97
        );

    \I__6155\ : Odrv4
    port map (
            O => \N__27739\,
            I => data_in_field_97
        );

    \I__6154\ : Odrv4
    port map (
            O => \N__27736\,
            I => data_in_field_97
        );

    \I__6153\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27724\
        );

    \I__6152\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27721\
        );

    \I__6151\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27717\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27714\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__27721\,
            I => \N__27711\
        );

    \I__6148\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27708\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__27717\,
            I => \N__27705\
        );

    \I__6146\ : Span4Mux_s3_h
    port map (
            O => \N__27714\,
            I => \N__27698\
        );

    \I__6145\ : Span4Mux_s2_v
    port map (
            O => \N__27711\,
            I => \N__27698\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__27708\,
            I => \N__27693\
        );

    \I__6143\ : Span4Mux_s2_v
    port map (
            O => \N__27705\,
            I => \N__27693\
        );

    \I__6142\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27690\
        );

    \I__6141\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27687\
        );

    \I__6140\ : Span4Mux_v
    port map (
            O => \N__27698\,
            I => \N__27684\
        );

    \I__6139\ : Span4Mux_v
    port map (
            O => \N__27693\,
            I => \N__27679\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__27690\,
            I => \N__27679\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__27687\,
            I => data_in_field_95
        );

    \I__6136\ : Odrv4
    port map (
            O => \N__27684\,
            I => data_in_field_95
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__27679\,
            I => data_in_field_95
        );

    \I__6134\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27668\
        );

    \I__6133\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27663\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__27668\,
            I => \N__27660\
        );

    \I__6131\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27654\
        );

    \I__6130\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27654\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27651\
        );

    \I__6128\ : Span4Mux_s3_v
    port map (
            O => \N__27660\,
            I => \N__27648\
        );

    \I__6127\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27643\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__27654\,
            I => \N__27640\
        );

    \I__6125\ : Span4Mux_s3_v
    port map (
            O => \N__27651\,
            I => \N__27635\
        );

    \I__6124\ : Span4Mux_h
    port map (
            O => \N__27648\,
            I => \N__27635\
        );

    \I__6123\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27630\
        );

    \I__6122\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27630\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__27643\,
            I => data_in_field_96
        );

    \I__6120\ : Odrv12
    port map (
            O => \N__27640\,
            I => data_in_field_96
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__27635\,
            I => data_in_field_96
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__27630\,
            I => data_in_field_96
        );

    \I__6117\ : CascadeMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__6116\ : InMux
    port map (
            O => \N__27618\,
            I => \N__27615\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__27615\,
            I => \N__27611\
        );

    \I__6114\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27608\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__27611\,
            I => \N__27605\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27602\
        );

    \I__6111\ : Span4Mux_v
    port map (
            O => \N__27605\,
            I => \N__27599\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__27602\,
            I => \c0.n4296\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__27599\,
            I => \c0.n4296\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__6107\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27588\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__27588\,
            I => \c0.rx.n12\
        );

    \I__6105\ : IoInMux
    port map (
            O => \N__27585\,
            I => \N__27582\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__27582\,
            I => \N__27579\
        );

    \I__6103\ : Span4Mux_s0_v
    port map (
            O => \N__27579\,
            I => \N__27576\
        );

    \I__6102\ : Span4Mux_h
    port map (
            O => \N__27576\,
            I => \N__27573\
        );

    \I__6101\ : Odrv4
    port map (
            O => \N__27573\,
            I => tx_enable
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__27570\,
            I => \N__27565\
        );

    \I__6099\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27562\
        );

    \I__6098\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27557\
        );

    \I__6097\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27557\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__27562\,
            I => n2185
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__27557\,
            I => n2185
        );

    \I__6094\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27548\
        );

    \I__6093\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27545\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__27548\,
            I => \N__27539\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27539\
        );

    \I__6090\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27536\
        );

    \I__6089\ : Span4Mux_h
    port map (
            O => \N__27539\,
            I => \N__27530\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__27536\,
            I => \N__27530\
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__27535\,
            I => \N__27526\
        );

    \I__6086\ : Span4Mux_v
    port map (
            O => \N__27530\,
            I => \N__27523\
        );

    \I__6085\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27520\
        );

    \I__6084\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27515\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__27523\,
            I => \N__27512\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27509\
        );

    \I__6081\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27504\
        );

    \I__6080\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27504\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__27515\,
            I => \r_Bit_Index_2_adj_1731\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__27512\,
            I => \r_Bit_Index_2_adj_1731\
        );

    \I__6077\ : Odrv12
    port map (
            O => \N__27509\,
            I => \r_Bit_Index_2_adj_1731\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__27504\,
            I => \r_Bit_Index_2_adj_1731\
        );

    \I__6075\ : CascadeMux
    port map (
            O => \N__27495\,
            I => \n7415_cascade_\
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__27492\,
            I => \n9301_cascade_\
        );

    \I__6073\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__6071\ : Odrv12
    port map (
            O => \N__27483\,
            I => \c0.n20_adj_1642\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__27480\,
            I => \n12_adj_1753_cascade_\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__27477\,
            I => \r_SM_Main_2_N_1537_2_cascade_\
        );

    \I__6068\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27470\
        );

    \I__6067\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27467\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__27470\,
            I => \N__27464\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__27467\,
            I => \N__27461\
        );

    \I__6064\ : Span4Mux_h
    port map (
            O => \N__27464\,
            I => \N__27458\
        );

    \I__6063\ : Span12Mux_s9_h
    port map (
            O => \N__27461\,
            I => \N__27455\
        );

    \I__6062\ : Span4Mux_v
    port map (
            O => \N__27458\,
            I => \N__27452\
        );

    \I__6061\ : Odrv12
    port map (
            O => \N__27455\,
            I => \c0.rx.n4090\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__27452\,
            I => \c0.rx.n4090\
        );

    \I__6059\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27444\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__6057\ : Span4Mux_h
    port map (
            O => \N__27441\,
            I => \N__27437\
        );

    \I__6056\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27434\
        );

    \I__6055\ : Odrv4
    port map (
            O => \N__27437\,
            I => \c0.rx.n7393\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__27434\,
            I => \c0.rx.n7393\
        );

    \I__6053\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27426\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__27426\,
            I => \N__27422\
        );

    \I__6051\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27419\
        );

    \I__6050\ : Span4Mux_s3_v
    port map (
            O => \N__27422\,
            I => \N__27416\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27413\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__27416\,
            I => \N__27405\
        );

    \I__6047\ : Span4Mux_s3_v
    port map (
            O => \N__27413\,
            I => \N__27405\
        );

    \I__6046\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27400\
        );

    \I__6045\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27400\
        );

    \I__6044\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27397\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__27405\,
            I => data_in_field_122
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__27400\,
            I => data_in_field_122
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__27397\,
            I => data_in_field_122
        );

    \I__6040\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27387\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27384\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__6037\ : Span4Mux_v
    port map (
            O => \N__27381\,
            I => \N__27378\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__27378\,
            I => \c0.n4537\
        );

    \I__6035\ : CascadeMux
    port map (
            O => \N__27375\,
            I => \c0.rx.r_SM_Main_2_N_1543_0_cascade_\
        );

    \I__6034\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27368\
        );

    \I__6033\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27365\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__27368\,
            I => \N__27362\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__27365\,
            I => \N__27359\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__27362\,
            I => \N__27356\
        );

    \I__6029\ : Span4Mux_h
    port map (
            O => \N__27359\,
            I => \N__27353\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__27356\,
            I => \N__27350\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__27353\,
            I => \c0.n8782\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__27350\,
            I => \c0.n8782\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__6024\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27339\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__27339\,
            I => \N__27336\
        );

    \I__6022\ : Span12Mux_v
    port map (
            O => \N__27336\,
            I => \N__27333\
        );

    \I__6021\ : Odrv12
    port map (
            O => \N__27333\,
            I => \c0.n8807\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__27330\,
            I => \N__27324\
        );

    \I__6019\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27321\
        );

    \I__6018\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27318\
        );

    \I__6017\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27315\
        );

    \I__6016\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27312\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__27321\,
            I => \N__27309\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__27318\,
            I => \N__27304\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__27315\,
            I => \N__27301\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__27312\,
            I => \N__27298\
        );

    \I__6011\ : Span4Mux_v
    port map (
            O => \N__27309\,
            I => \N__27295\
        );

    \I__6010\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27290\
        );

    \I__6009\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27290\
        );

    \I__6008\ : Span4Mux_s2_v
    port map (
            O => \N__27304\,
            I => \N__27285\
        );

    \I__6007\ : Span4Mux_s2_v
    port map (
            O => \N__27301\,
            I => \N__27285\
        );

    \I__6006\ : Odrv12
    port map (
            O => \N__27298\,
            I => data_in_field_110
        );

    \I__6005\ : Odrv4
    port map (
            O => \N__27295\,
            I => data_in_field_110
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__27290\,
            I => data_in_field_110
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__27285\,
            I => data_in_field_110
        );

    \I__6002\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27273\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__27273\,
            I => \c0.n8819\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__27270\,
            I => \N__27266\
        );

    \I__5999\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27263\
        );

    \I__5998\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27260\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27257\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27254\
        );

    \I__5995\ : Span4Mux_v
    port map (
            O => \N__27257\,
            I => \N__27251\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__27254\,
            I => \N__27248\
        );

    \I__5993\ : Span4Mux_s3_h
    port map (
            O => \N__27251\,
            I => \N__27245\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__27248\,
            I => \c0.n8893\
        );

    \I__5991\ : Odrv4
    port map (
            O => \N__27245\,
            I => \c0.n8893\
        );

    \I__5990\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27237\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__5988\ : Span12Mux_s7_v
    port map (
            O => \N__27234\,
            I => \N__27230\
        );

    \I__5987\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27227\
        );

    \I__5986\ : Odrv12
    port map (
            O => \N__27230\,
            I => \c0.n8427\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__27227\,
            I => \c0.n8427\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27219\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__5982\ : Odrv12
    port map (
            O => \N__27216\,
            I => \c0.n28_adj_1612\
        );

    \I__5981\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__27210\,
            I => \c0.n26_adj_1613\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__27207\,
            I => \c0.n27_cascade_\
        );

    \I__5978\ : InMux
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27198\
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__27198\,
            I => \c0.n25_adj_1614\
        );

    \I__5975\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__5973\ : Odrv12
    port map (
            O => \N__27189\,
            I => \c0.data_in_frame_20_0\
        );

    \I__5972\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__27183\,
            I => \N__27180\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__5969\ : Span4Mux_h
    port map (
            O => \N__27177\,
            I => \N__27173\
        );

    \I__5968\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27170\
        );

    \I__5967\ : Span4Mux_h
    port map (
            O => \N__27173\,
            I => \N__27167\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__27170\,
            I => \c0.n8995\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__27167\,
            I => \c0.n8995\
        );

    \I__5964\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27156\
        );

    \I__5963\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27156\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__27156\,
            I => \N__27153\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__27150\,
            I => \c0.n8834\
        );

    \I__5959\ : CascadeMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__5958\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__5956\ : Span4Mux_h
    port map (
            O => \N__27138\,
            I => \N__27134\
        );

    \I__5955\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27131\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__27134\,
            I => \N__27128\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__27131\,
            I => \c0.n8924\
        );

    \I__5952\ : Odrv4
    port map (
            O => \N__27128\,
            I => \c0.n8924\
        );

    \I__5951\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27116\
        );

    \I__5949\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27113\
        );

    \I__5948\ : Span12Mux_s10_v
    port map (
            O => \N__27116\,
            I => \N__27110\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__27113\,
            I => \N__27107\
        );

    \I__5946\ : Odrv12
    port map (
            O => \N__27110\,
            I => \c0.n8852\
        );

    \I__5945\ : Odrv4
    port map (
            O => \N__27107\,
            I => \c0.n8852\
        );

    \I__5944\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27099\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__27099\,
            I => \N__27095\
        );

    \I__5942\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27092\
        );

    \I__5941\ : Span4Mux_h
    port map (
            O => \N__27095\,
            I => \N__27089\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__27092\,
            I => \N__27086\
        );

    \I__5939\ : Odrv4
    port map (
            O => \N__27089\,
            I => \c0.n9013\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__27086\,
            I => \c0.n9013\
        );

    \I__5937\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27078\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__27078\,
            I => \N__27074\
        );

    \I__5935\ : InMux
    port map (
            O => \N__27077\,
            I => \N__27071\
        );

    \I__5934\ : Span4Mux_s2_v
    port map (
            O => \N__27074\,
            I => \N__27068\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__27071\,
            I => \N__27063\
        );

    \I__5932\ : Span4Mux_v
    port map (
            O => \N__27068\,
            I => \N__27060\
        );

    \I__5931\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27055\
        );

    \I__5930\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27055\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__27063\,
            I => data_in_field_70
        );

    \I__5928\ : Odrv4
    port map (
            O => \N__27060\,
            I => data_in_field_70
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__27055\,
            I => data_in_field_70
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__27048\,
            I => \c0.n12_cascade_\
        );

    \I__5925\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27042\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__27042\,
            I => \N__27038\
        );

    \I__5923\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27035\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__27038\,
            I => \N__27030\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__27035\,
            I => \N__27027\
        );

    \I__5920\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27024\
        );

    \I__5919\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27021\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__27030\,
            I => \N__27016\
        );

    \I__5917\ : Span4Mux_h
    port map (
            O => \N__27027\,
            I => \N__27016\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__27024\,
            I => data_in_field_112
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__27021\,
            I => data_in_field_112
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__27016\,
            I => data_in_field_112
        );

    \I__5913\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27006\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__27006\,
            I => \c0.data_in_frame_20_2\
        );

    \I__5911\ : InMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__5909\ : Span4Mux_v
    port map (
            O => \N__26997\,
            I => \N__26992\
        );

    \I__5908\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26987\
        );

    \I__5907\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26987\
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__26992\,
            I => data_in_5_2
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__26987\,
            I => data_in_5_2
        );

    \I__5904\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__26979\,
            I => \N__26975\
        );

    \I__5902\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26972\
        );

    \I__5901\ : Span4Mux_s3_h
    port map (
            O => \N__26975\,
            I => \N__26969\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__26972\,
            I => \N__26966\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__26969\,
            I => \N__26963\
        );

    \I__5898\ : Span4Mux_h
    port map (
            O => \N__26966\,
            I => \N__26960\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__26963\,
            I => \N__26956\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__26960\,
            I => \N__26953\
        );

    \I__5895\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26950\
        );

    \I__5894\ : Odrv4
    port map (
            O => \N__26956\,
            I => data_in_4_2
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__26953\,
            I => data_in_4_2
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__26950\,
            I => data_in_4_2
        );

    \I__5891\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26939\
        );

    \I__5890\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26935\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__26939\,
            I => \N__26931\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26928\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__26935\,
            I => \N__26925\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__26934\,
            I => \N__26922\
        );

    \I__5885\ : Span4Mux_h
    port map (
            O => \N__26931\,
            I => \N__26914\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26911\
        );

    \I__5883\ : Span12Mux_h
    port map (
            O => \N__26925\,
            I => \N__26908\
        );

    \I__5882\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26905\
        );

    \I__5881\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26898\
        );

    \I__5880\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26898\
        );

    \I__5879\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26898\
        );

    \I__5878\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26893\
        );

    \I__5877\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26893\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__26914\,
            I => \r_SM_Main_2_adj_1738\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__26911\,
            I => \r_SM_Main_2_adj_1738\
        );

    \I__5874\ : Odrv12
    port map (
            O => \N__26908\,
            I => \r_SM_Main_2_adj_1738\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__26905\,
            I => \r_SM_Main_2_adj_1738\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__26898\,
            I => \r_SM_Main_2_adj_1738\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__26893\,
            I => \r_SM_Main_2_adj_1738\
        );

    \I__5870\ : CEMux
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26873\
        );

    \I__5868\ : CEMux
    port map (
            O => \N__26876\,
            I => \N__26870\
        );

    \I__5867\ : Span4Mux_s1_v
    port map (
            O => \N__26873\,
            I => \N__26865\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__26870\,
            I => \N__26865\
        );

    \I__5865\ : Span4Mux_s1_h
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__5864\ : Span4Mux_h
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__5863\ : Span4Mux_h
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__26856\,
            I => \c0.tx2.n4880\
        );

    \I__5861\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26850\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__5859\ : Span4Mux_v
    port map (
            O => \N__26847\,
            I => \N__26844\
        );

    \I__5858\ : Span4Mux_h
    port map (
            O => \N__26844\,
            I => \N__26841\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__26841\,
            I => \c0.n4525\
        );

    \I__5856\ : CascadeMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__5855\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26832\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__26826\,
            I => \c0.n4244\
        );

    \I__5851\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26817\
        );

    \I__5849\ : Span4Mux_v
    port map (
            O => \N__26817\,
            I => \N__26810\
        );

    \I__5848\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26805\
        );

    \I__5847\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26805\
        );

    \I__5846\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26802\
        );

    \I__5845\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26799\
        );

    \I__5844\ : Span4Mux_h
    port map (
            O => \N__26810\,
            I => \N__26794\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26794\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__26802\,
            I => data_in_field_50
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__26799\,
            I => data_in_field_50
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__26794\,
            I => data_in_field_50
        );

    \I__5839\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26784\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__26784\,
            I => \N__26780\
        );

    \I__5837\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26777\
        );

    \I__5836\ : Odrv12
    port map (
            O => \N__26780\,
            I => \c0.n8918\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__26777\,
            I => \c0.n8918\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__26772\,
            I => \c0.n8840_cascade_\
        );

    \I__5833\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26765\
        );

    \I__5832\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26762\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__26765\,
            I => \c0.n4511\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__26762\,
            I => \c0.n4511\
        );

    \I__5829\ : InMux
    port map (
            O => \N__26757\,
            I => \N__26754\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__5827\ : Span12Mux_s7_h
    port map (
            O => \N__26751\,
            I => \N__26747\
        );

    \I__5826\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26744\
        );

    \I__5825\ : Odrv12
    port map (
            O => \N__26747\,
            I => \c0.n4309\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__26744\,
            I => \c0.n4309\
        );

    \I__5823\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26735\
        );

    \I__5822\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26732\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26729\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26725\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__26729\,
            I => \N__26722\
        );

    \I__5818\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26718\
        );

    \I__5817\ : Span4Mux_v
    port map (
            O => \N__26725\,
            I => \N__26714\
        );

    \I__5816\ : Sp12to4
    port map (
            O => \N__26722\,
            I => \N__26711\
        );

    \I__5815\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26708\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26705\
        );

    \I__5813\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26702\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__26714\,
            I => rand_data_11
        );

    \I__5811\ : Odrv12
    port map (
            O => \N__26711\,
            I => rand_data_11
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__26708\,
            I => rand_data_11
        );

    \I__5809\ : Odrv12
    port map (
            O => \N__26705\,
            I => rand_data_11
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__26702\,
            I => rand_data_11
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__26691\,
            I => \N__26686\
        );

    \I__5806\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26680\
        );

    \I__5805\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26680\
        );

    \I__5804\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26677\
        );

    \I__5803\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26674\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__26680\,
            I => \N__26671\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26668\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__26674\,
            I => \N__26665\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__26671\,
            I => \N__26660\
        );

    \I__5798\ : Span4Mux_s3_h
    port map (
            O => \N__26668\,
            I => \N__26660\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__26665\,
            I => \N__26656\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__26660\,
            I => \N__26651\
        );

    \I__5795\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26648\
        );

    \I__5794\ : Sp12to4
    port map (
            O => \N__26656\,
            I => \N__26645\
        );

    \I__5793\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26640\
        );

    \I__5792\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26640\
        );

    \I__5791\ : Span4Mux_v
    port map (
            O => \N__26651\,
            I => \N__26637\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__26648\,
            I => data_in_field_123
        );

    \I__5789\ : Odrv12
    port map (
            O => \N__26645\,
            I => data_in_field_123
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__26640\,
            I => data_in_field_123
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__26637\,
            I => data_in_field_123
        );

    \I__5786\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26624\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__26627\,
            I => \N__26620\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26616\
        );

    \I__5783\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26613\
        );

    \I__5782\ : InMux
    port map (
            O => \N__26620\,
            I => \N__26607\
        );

    \I__5781\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26607\
        );

    \I__5780\ : Span4Mux_h
    port map (
            O => \N__26616\,
            I => \N__26602\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__26613\,
            I => \N__26599\
        );

    \I__5778\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26596\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__26607\,
            I => \N__26593\
        );

    \I__5776\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26588\
        );

    \I__5775\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26585\
        );

    \I__5774\ : Span4Mux_v
    port map (
            O => \N__26602\,
            I => \N__26578\
        );

    \I__5773\ : Span4Mux_h
    port map (
            O => \N__26599\,
            I => \N__26578\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26578\
        );

    \I__5771\ : Span12Mux_s8_h
    port map (
            O => \N__26593\,
            I => \N__26575\
        );

    \I__5770\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26572\
        );

    \I__5769\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26569\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__26588\,
            I => data_in_field_146
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__26585\,
            I => data_in_field_146
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__26578\,
            I => data_in_field_146
        );

    \I__5765\ : Odrv12
    port map (
            O => \N__26575\,
            I => data_in_field_146
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__26572\,
            I => data_in_field_146
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__26569\,
            I => data_in_field_146
        );

    \I__5762\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26551\
        );

    \I__5761\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26548\
        );

    \I__5760\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26545\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__26551\,
            I => \N__26542\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__26548\,
            I => \N__26536\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__26545\,
            I => \N__26536\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__26542\,
            I => \N__26533\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__26541\,
            I => \N__26529\
        );

    \I__5754\ : Span4Mux_v
    port map (
            O => \N__26536\,
            I => \N__26526\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__26533\,
            I => \N__26523\
        );

    \I__5752\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26518\
        );

    \I__5751\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26518\
        );

    \I__5750\ : Span4Mux_h
    port map (
            O => \N__26526\,
            I => \N__26515\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__26523\,
            I => data_in_field_130
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__26518\,
            I => data_in_field_130
        );

    \I__5747\ : Odrv4
    port map (
            O => \N__26515\,
            I => data_in_field_130
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__26508\,
            I => \c0.n9698_cascade_\
        );

    \I__5745\ : InMux
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26497\
        );

    \I__5743\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26494\
        );

    \I__5742\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26491\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__26497\,
            I => \N__26486\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26486\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__26491\,
            I => \N__26481\
        );

    \I__5738\ : Span4Mux_h
    port map (
            O => \N__26486\,
            I => \N__26478\
        );

    \I__5737\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26473\
        );

    \I__5736\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26473\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__26481\,
            I => data_in_field_138
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__26478\,
            I => data_in_field_138
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__26473\,
            I => data_in_field_138
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__26466\,
            I => \c0.n9701_cascade_\
        );

    \I__5731\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26458\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__26462\,
            I => \N__26454\
        );

    \I__5729\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26451\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__26458\,
            I => \N__26448\
        );

    \I__5727\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26445\
        );

    \I__5726\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26442\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__26451\,
            I => \N__26438\
        );

    \I__5724\ : Span4Mux_v
    port map (
            O => \N__26448\,
            I => \N__26433\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26433\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__26442\,
            I => \N__26430\
        );

    \I__5721\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26427\
        );

    \I__5720\ : Span4Mux_h
    port map (
            O => \N__26438\,
            I => \N__26424\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__26433\,
            I => \N__26421\
        );

    \I__5718\ : Span4Mux_v
    port map (
            O => \N__26430\,
            I => \N__26418\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__26427\,
            I => data_in_field_142
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__26424\,
            I => data_in_field_142
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__26421\,
            I => data_in_field_142
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__26418\,
            I => data_in_field_142
        );

    \I__5713\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26405\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__26408\,
            I => \N__26401\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__26405\,
            I => \N__26398\
        );

    \I__5710\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26394\
        );

    \I__5709\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26391\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__26398\,
            I => \N__26388\
        );

    \I__5707\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26385\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__26394\,
            I => \N__26382\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__26391\,
            I => \N__26377\
        );

    \I__5704\ : IoSpan4Mux
    port map (
            O => \N__26388\,
            I => \N__26374\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__26385\,
            I => \N__26371\
        );

    \I__5702\ : Span4Mux_s1_v
    port map (
            O => \N__26382\,
            I => \N__26368\
        );

    \I__5701\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26365\
        );

    \I__5700\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26362\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__26377\,
            I => \N__26353\
        );

    \I__5698\ : Span4Mux_s3_h
    port map (
            O => \N__26374\,
            I => \N__26353\
        );

    \I__5697\ : Span4Mux_v
    port map (
            O => \N__26371\,
            I => \N__26353\
        );

    \I__5696\ : Span4Mux_v
    port map (
            O => \N__26368\,
            I => \N__26353\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__26365\,
            I => data_in_field_78
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__26362\,
            I => data_in_field_78
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__26353\,
            I => data_in_field_78
        );

    \I__5692\ : InMux
    port map (
            O => \N__26346\,
            I => \N__26342\
        );

    \I__5691\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26339\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__26342\,
            I => \N__26336\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26333\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__26336\,
            I => \N__26330\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__26333\,
            I => \N__26326\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__26330\,
            I => \N__26323\
        );

    \I__5685\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26320\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__26326\,
            I => \c0.n4215\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__26323\,
            I => \c0.n4215\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__26320\,
            I => \c0.n4215\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__5680\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26307\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26304\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__26304\,
            I => \N__26300\
        );

    \I__5677\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26297\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__26300\,
            I => \c0.n8912\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__26297\,
            I => \c0.n8912\
        );

    \I__5674\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26288\
        );

    \I__5673\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26285\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26282\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26279\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__26282\,
            I => \c0.n8954\
        );

    \I__5669\ : Odrv12
    port map (
            O => \N__26279\,
            I => \c0.n8954\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__26274\,
            I => \c0.n8819_cascade_\
        );

    \I__5667\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26268\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__26268\,
            I => \N__26264\
        );

    \I__5665\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26261\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__26264\,
            I => \c0.n4365\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26261\,
            I => \c0.n4365\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__26256\,
            I => \c0.n21_adj_1644_cascade_\
        );

    \I__5661\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__26241\,
            I => \c0.n19_adj_1643\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \N__26235\
        );

    \I__5655\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__26232\,
            I => \c0.data_in_frame_19_2\
        );

    \I__5653\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__26226\,
            I => \c0.data_in_frame_19_0\
        );

    \I__5651\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26220\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__26220\,
            I => \N__26216\
        );

    \I__5649\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26213\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__26216\,
            I => \N__26207\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26207\
        );

    \I__5646\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26203\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__26207\,
            I => \N__26200\
        );

    \I__5644\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26197\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__26203\,
            I => data_in_field_136
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__26200\,
            I => data_in_field_136
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__26197\,
            I => data_in_field_136
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__26190\,
            I => \c0.n9536_cascade_\
        );

    \I__5639\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26183\
        );

    \I__5638\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26180\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26176\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26173\
        );

    \I__5635\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26169\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__26176\,
            I => \N__26164\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__26173\,
            I => \N__26164\
        );

    \I__5632\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26161\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__26169\,
            I => data_in_field_128
        );

    \I__5630\ : Odrv4
    port map (
            O => \N__26164\,
            I => data_in_field_128
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__26161\,
            I => data_in_field_128
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__26154\,
            I => \c0.n9539_cascade_\
        );

    \I__5627\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26148\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__26148\,
            I => \N__26143\
        );

    \I__5625\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26140\
        );

    \I__5624\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26137\
        );

    \I__5623\ : Span4Mux_v
    port map (
            O => \N__26143\,
            I => \N__26132\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__26140\,
            I => \N__26132\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__26137\,
            I => \N__26127\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__26132\,
            I => \N__26127\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__26127\,
            I => \N__26123\
        );

    \I__5618\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26120\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__26123\,
            I => rand_data_18
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__26120\,
            I => rand_data_18
        );

    \I__5615\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26112\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__26109\
        );

    \I__5613\ : Span4Mux_s2_v
    port map (
            O => \N__26109\,
            I => \N__26105\
        );

    \I__5612\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26102\
        );

    \I__5611\ : Span4Mux_h
    port map (
            O => \N__26105\,
            I => \N__26097\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26097\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__26097\,
            I => \N__26092\
        );

    \I__5608\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26087\
        );

    \I__5607\ : InMux
    port map (
            O => \N__26095\,
            I => \N__26087\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__26092\,
            I => data_in_field_114
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__26087\,
            I => data_in_field_114
        );

    \I__5604\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26076\
        );

    \I__5603\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26073\
        );

    \I__5602\ : InMux
    port map (
            O => \N__26080\,
            I => \N__26070\
        );

    \I__5601\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26067\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26062\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__26073\,
            I => \N__26062\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26057\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__26067\,
            I => \N__26054\
        );

    \I__5596\ : Span4Mux_v
    port map (
            O => \N__26062\,
            I => \N__26051\
        );

    \I__5595\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26046\
        );

    \I__5594\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26046\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__26057\,
            I => \N__26043\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__26054\,
            I => \N__26038\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__26051\,
            I => \N__26038\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__26046\,
            I => data_in_field_144
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__26043\,
            I => data_in_field_144
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__26038\,
            I => data_in_field_144
        );

    \I__5587\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26027\
        );

    \I__5586\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26024\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__26027\,
            I => \N__26021\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__26021\,
            I => \N__26015\
        );

    \I__5582\ : Span4Mux_v
    port map (
            O => \N__26018\,
            I => \N__26012\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__26015\,
            I => \N__26009\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__26012\,
            I => \c0.n8971\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__26009\,
            I => \c0.n8971\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26004\,
            I => \N__26001\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__26001\,
            I => \c0.n6_adj_1628\
        );

    \I__5576\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25994\
        );

    \I__5575\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25991\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__25994\,
            I => \N__25988\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25984\
        );

    \I__5572\ : Span4Mux_h
    port map (
            O => \N__25988\,
            I => \N__25981\
        );

    \I__5571\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25978\
        );

    \I__5570\ : Span4Mux_v
    port map (
            O => \N__25984\,
            I => \N__25973\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__25981\,
            I => \N__25970\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__25978\,
            I => \N__25967\
        );

    \I__5567\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25964\
        );

    \I__5566\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25961\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__25973\,
            I => rand_data_0
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__25970\,
            I => rand_data_0
        );

    \I__5563\ : Odrv4
    port map (
            O => \N__25967\,
            I => rand_data_0
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__25964\,
            I => rand_data_0
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__25961\,
            I => rand_data_0
        );

    \I__5560\ : InMux
    port map (
            O => \N__25950\,
            I => \N__25938\
        );

    \I__5559\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25938\
        );

    \I__5558\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25938\
        );

    \I__5557\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25938\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__25938\,
            I => n9077
        );

    \I__5555\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25929\
        );

    \I__5554\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25929\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__25929\,
            I => n5185
        );

    \I__5552\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25922\
        );

    \I__5551\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25919\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__25922\,
            I => \N__25916\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25913\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__25916\,
            I => \N__25910\
        );

    \I__5547\ : Span4Mux_h
    port map (
            O => \N__25913\,
            I => \N__25907\
        );

    \I__5546\ : Span4Mux_v
    port map (
            O => \N__25910\,
            I => \N__25903\
        );

    \I__5545\ : Span4Mux_v
    port map (
            O => \N__25907\,
            I => \N__25900\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \N__25897\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__25903\,
            I => \N__25892\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__25900\,
            I => \N__25889\
        );

    \I__5541\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25882\
        );

    \I__5540\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25882\
        );

    \I__5539\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25882\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__25892\,
            I => \r_Bit_Index_0_adj_1733\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__25889\,
            I => \r_Bit_Index_0_adj_1733\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__25882\,
            I => \r_Bit_Index_0_adj_1733\
        );

    \I__5535\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25870\
        );

    \I__5534\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25867\
        );

    \I__5533\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25864\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__25870\,
            I => \N__25860\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__25867\,
            I => \N__25855\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__25864\,
            I => \N__25855\
        );

    \I__5529\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25852\
        );

    \I__5528\ : Span4Mux_v
    port map (
            O => \N__25860\,
            I => \N__25849\
        );

    \I__5527\ : Span12Mux_s8_h
    port map (
            O => \N__25855\,
            I => \N__25844\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__25852\,
            I => \N__25844\
        );

    \I__5525\ : Span4Mux_v
    port map (
            O => \N__25849\,
            I => \N__25839\
        );

    \I__5524\ : Span12Mux_v
    port map (
            O => \N__25844\,
            I => \N__25836\
        );

    \I__5523\ : InMux
    port map (
            O => \N__25843\,
            I => \N__25831\
        );

    \I__5522\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25831\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__25839\,
            I => \r_Bit_Index_1_adj_1732\
        );

    \I__5520\ : Odrv12
    port map (
            O => \N__25836\,
            I => \r_Bit_Index_1_adj_1732\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__25831\,
            I => \r_Bit_Index_1_adj_1732\
        );

    \I__5518\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25818\
        );

    \I__5517\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25818\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__25815\,
            I => \N__25812\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__25812\,
            I => n4_adj_1724
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__25809\,
            I => \N__25805\
        );

    \I__5512\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25801\
        );

    \I__5511\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25798\
        );

    \I__5510\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25795\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__25801\,
            I => \N__25792\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__25798\,
            I => \N__25788\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__25795\,
            I => \N__25785\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__25792\,
            I => \N__25781\
        );

    \I__5505\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25778\
        );

    \I__5504\ : Span4Mux_v
    port map (
            O => \N__25788\,
            I => \N__25773\
        );

    \I__5503\ : Span4Mux_v
    port map (
            O => \N__25785\,
            I => \N__25773\
        );

    \I__5502\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25770\
        );

    \I__5501\ : Span4Mux_v
    port map (
            O => \N__25781\,
            I => \N__25767\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25764\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__25773\,
            I => \N__25761\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__25770\,
            I => data_in_field_134
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__25767\,
            I => data_in_field_134
        );

    \I__5496\ : Odrv12
    port map (
            O => \N__25764\,
            I => data_in_field_134
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__25761\,
            I => data_in_field_134
        );

    \I__5494\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__25746\,
            I => \N__25742\
        );

    \I__5491\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25737\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__25742\,
            I => \N__25734\
        );

    \I__5489\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25729\
        );

    \I__5488\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25729\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__25737\,
            I => data_in_field_119
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__25734\,
            I => data_in_field_119
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__25729\,
            I => data_in_field_119
        );

    \I__5484\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25719\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__25719\,
            I => \N__25715\
        );

    \I__5482\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25712\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__25715\,
            I => \N__25706\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__25712\,
            I => \N__25706\
        );

    \I__5479\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25703\
        );

    \I__5478\ : Span4Mux_v
    port map (
            O => \N__25706\,
            I => \N__25700\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__25703\,
            I => \N__25697\
        );

    \I__5476\ : Span4Mux_s3_h
    port map (
            O => \N__25700\,
            I => \N__25694\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__25697\,
            I => \N__25691\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__25694\,
            I => \c0.n8883\
        );

    \I__5473\ : Odrv4
    port map (
            O => \N__25691\,
            I => \c0.n8883\
        );

    \I__5472\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__25683\,
            I => \N__25680\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__25680\,
            I => \c0.n8770\
        );

    \I__5469\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25674\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__25674\,
            I => \N__25670\
        );

    \I__5467\ : CascadeMux
    port map (
            O => \N__25673\,
            I => \N__25667\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__25670\,
            I => \N__25664\
        );

    \I__5465\ : InMux
    port map (
            O => \N__25667\,
            I => \N__25661\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__25664\,
            I => \N__25656\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__25661\,
            I => \N__25656\
        );

    \I__5462\ : Span4Mux_h
    port map (
            O => \N__25656\,
            I => \N__25653\
        );

    \I__5461\ : Span4Mux_v
    port map (
            O => \N__25653\,
            I => \N__25650\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__25650\,
            I => \c0.n8810\
        );

    \I__5459\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__25644\,
            I => \N__25641\
        );

    \I__5457\ : Span4Mux_v
    port map (
            O => \N__25641\,
            I => \N__25637\
        );

    \I__5456\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25634\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__25637\,
            I => \N__25629\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__25634\,
            I => \N__25629\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__25629\,
            I => \N__25626\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__25626\,
            I => \c0.n8899\
        );

    \I__5451\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__25620\,
            I => \c0.n16_adj_1657\
        );

    \I__5449\ : CascadeMux
    port map (
            O => \N__25617\,
            I => \c0.n22_adj_1655_cascade_\
        );

    \I__5448\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25608\
        );

    \I__5447\ : InMux
    port map (
            O => \N__25613\,
            I => \N__25605\
        );

    \I__5446\ : CascadeMux
    port map (
            O => \N__25612\,
            I => \N__25600\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__25611\,
            I => \N__25597\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25594\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__25605\,
            I => \N__25591\
        );

    \I__5442\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25586\
        );

    \I__5441\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25586\
        );

    \I__5440\ : InMux
    port map (
            O => \N__25600\,
            I => \N__25581\
        );

    \I__5439\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25581\
        );

    \I__5438\ : Odrv12
    port map (
            O => \N__25594\,
            I => data_in_field_37
        );

    \I__5437\ : Odrv4
    port map (
            O => \N__25591\,
            I => data_in_field_37
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__25586\,
            I => data_in_field_37
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__25581\,
            I => data_in_field_37
        );

    \I__5434\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__25569\,
            I => \c0.n24_adj_1658\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__25566\,
            I => \N__25563\
        );

    \I__5431\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__25557\,
            I => \N__25554\
        );

    \I__5428\ : Span4Mux_h
    port map (
            O => \N__25554\,
            I => \N__25550\
        );

    \I__5427\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25547\
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__25550\,
            I => \c0.n8939\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__25547\,
            I => \c0.n8939\
        );

    \I__5424\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__25539\,
            I => \N__25536\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__25530\,
            I => \c0.n20_adj_1659\
        );

    \I__5419\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25524\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__25524\,
            I => \N__25520\
        );

    \I__5417\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25517\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__25520\,
            I => \N__25514\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25508\
        );

    \I__5414\ : IoSpan4Mux
    port map (
            O => \N__25514\,
            I => \N__25505\
        );

    \I__5413\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25500\
        );

    \I__5412\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25500\
        );

    \I__5411\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25497\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__25508\,
            I => \N__25494\
        );

    \I__5409\ : Sp12to4
    port map (
            O => \N__25505\,
            I => \N__25489\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__25500\,
            I => \N__25489\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__25497\,
            I => data_in_field_68
        );

    \I__5406\ : Odrv4
    port map (
            O => \N__25494\,
            I => data_in_field_68
        );

    \I__5405\ : Odrv12
    port map (
            O => \N__25489\,
            I => data_in_field_68
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__25482\,
            I => \N__25477\
        );

    \I__5403\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25473\
        );

    \I__5402\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25470\
        );

    \I__5401\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25467\
        );

    \I__5400\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25464\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__25473\,
            I => \N__25461\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__25470\,
            I => \N__25458\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__25467\,
            I => \N__25455\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__25464\,
            I => \N__25445\
        );

    \I__5395\ : Span4Mux_h
    port map (
            O => \N__25461\,
            I => \N__25445\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__25458\,
            I => \N__25445\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__25455\,
            I => \N__25445\
        );

    \I__5392\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25442\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__25445\,
            I => data_in_field_76
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__25442\,
            I => data_in_field_76
        );

    \I__5389\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25434\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__25431\,
            I => \c0.n9566\
        );

    \I__5386\ : InMux
    port map (
            O => \N__25428\,
            I => \N__25425\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__25422\,
            I => \c0.n9171\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__25419\,
            I => \c0.n9168_cascade_\
        );

    \I__5382\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__5380\ : Span4Mux_s2_v
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__5379\ : Odrv4
    port map (
            O => \N__25407\,
            I => \c0.n9165\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__5377\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__5373\ : Sp12to4
    port map (
            O => \N__25389\,
            I => \N__25386\
        );

    \I__5372\ : Odrv12
    port map (
            O => \N__25386\,
            I => \c0.n9162\
        );

    \I__5371\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__25380\,
            I => \c0.n9554\
        );

    \I__5369\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__25371\,
            I => \c0.n22_adj_1679\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__25368\,
            I => \c0.n9557_cascade_\
        );

    \I__5365\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__5363\ : Span4Mux_s1_v
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__25353\,
            I => \c0.tx2.r_Tx_Data_4\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__25350\,
            I => \n5185_cascade_\
        );

    \I__5359\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25343\
        );

    \I__5358\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25340\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__25343\,
            I => \N__25335\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__25340\,
            I => \N__25331\
        );

    \I__5355\ : InMux
    port map (
            O => \N__25339\,
            I => \N__25328\
        );

    \I__5354\ : InMux
    port map (
            O => \N__25338\,
            I => \N__25325\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__25335\,
            I => \N__25322\
        );

    \I__5352\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25319\
        );

    \I__5351\ : Span4Mux_h
    port map (
            O => \N__25331\,
            I => \N__25315\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__25328\,
            I => \N__25310\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__25325\,
            I => \N__25310\
        );

    \I__5348\ : Span4Mux_v
    port map (
            O => \N__25322\,
            I => \N__25307\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__25319\,
            I => \N__25304\
        );

    \I__5346\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25300\
        );

    \I__5345\ : Span4Mux_h
    port map (
            O => \N__25315\,
            I => \N__25295\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__25310\,
            I => \N__25295\
        );

    \I__5343\ : Sp12to4
    port map (
            O => \N__25307\,
            I => \N__25290\
        );

    \I__5342\ : Span12Mux_s8_v
    port map (
            O => \N__25304\,
            I => \N__25290\
        );

    \I__5341\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25287\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__25300\,
            I => data_in_field_150
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__25295\,
            I => data_in_field_150
        );

    \I__5338\ : Odrv12
    port map (
            O => \N__25290\,
            I => data_in_field_150
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__25287\,
            I => data_in_field_150
        );

    \I__5336\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25272\
        );

    \I__5335\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25269\
        );

    \I__5334\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25266\
        );

    \I__5333\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25263\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__25272\,
            I => \N__25259\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25256\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__25266\,
            I => \N__25251\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__25263\,
            I => \N__25251\
        );

    \I__5328\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25247\
        );

    \I__5327\ : Span12Mux_s7_v
    port map (
            O => \N__25259\,
            I => \N__25244\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__25256\,
            I => \N__25241\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__25251\,
            I => \N__25238\
        );

    \I__5324\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25235\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__25247\,
            I => data_in_field_52
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__25244\,
            I => data_in_field_52
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__25241\,
            I => data_in_field_52
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__25238\,
            I => data_in_field_52
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__25235\,
            I => data_in_field_52
        );

    \I__5318\ : CascadeMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__5317\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25215\
        );

    \I__5316\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25210\
        );

    \I__5315\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25207\
        );

    \I__5314\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25204\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__25215\,
            I => \N__25201\
        );

    \I__5312\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25198\
        );

    \I__5311\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25195\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__25210\,
            I => \N__25190\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25190\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__25204\,
            I => \N__25183\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__25201\,
            I => \N__25183\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__25198\,
            I => \N__25183\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__25195\,
            I => \N__25180\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__25190\,
            I => \N__25177\
        );

    \I__5303\ : Span4Mux_v
    port map (
            O => \N__25183\,
            I => \N__25174\
        );

    \I__5302\ : Span4Mux_h
    port map (
            O => \N__25180\,
            I => \N__25171\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__25177\,
            I => \N__25167\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__25174\,
            I => \N__25161\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__25171\,
            I => \N__25161\
        );

    \I__5298\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25158\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__25167\,
            I => \N__25155\
        );

    \I__5296\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25152\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__25161\,
            I => \N__25149\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__25158\,
            I => data_in_field_151
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__25155\,
            I => data_in_field_151
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__25152\,
            I => data_in_field_151
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__25149\,
            I => data_in_field_151
        );

    \I__5290\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25135\
        );

    \I__5289\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25132\
        );

    \I__5288\ : CascadeMux
    port map (
            O => \N__25138\,
            I => \N__25129\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25125\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25122\
        );

    \I__5285\ : InMux
    port map (
            O => \N__25129\,
            I => \N__25119\
        );

    \I__5284\ : InMux
    port map (
            O => \N__25128\,
            I => \N__25115\
        );

    \I__5283\ : Span4Mux_s2_v
    port map (
            O => \N__25125\,
            I => \N__25112\
        );

    \I__5282\ : Span4Mux_s2_v
    port map (
            O => \N__25122\,
            I => \N__25109\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__25119\,
            I => \N__25106\
        );

    \I__5280\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25103\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25100\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__25112\,
            I => \N__25095\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__25109\,
            I => \N__25095\
        );

    \I__5276\ : Span4Mux_s3_v
    port map (
            O => \N__25106\,
            I => \N__25092\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__25103\,
            I => data_in_field_86
        );

    \I__5274\ : Odrv12
    port map (
            O => \N__25100\,
            I => data_in_field_86
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__25095\,
            I => data_in_field_86
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__25092\,
            I => data_in_field_86
        );

    \I__5271\ : InMux
    port map (
            O => \N__25083\,
            I => \N__25080\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__25080\,
            I => \N__25076\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__25079\,
            I => \N__25073\
        );

    \I__5268\ : Span4Mux_h
    port map (
            O => \N__25076\,
            I => \N__25070\
        );

    \I__5267\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25067\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__25070\,
            I => \N__25062\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25062\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__25062\,
            I => \c0.n8915\
        );

    \I__5263\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25053\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__25053\,
            I => \N__25050\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__25050\,
            I => \N__25047\
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__25047\,
            I => \c0.n8788\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__5257\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__25035\,
            I => \N__25031\
        );

    \I__5254\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25028\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__25031\,
            I => \c0.n8828\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__25028\,
            I => \c0.n8828\
        );

    \I__5251\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__25020\,
            I => \N__25016\
        );

    \I__5249\ : InMux
    port map (
            O => \N__25019\,
            I => \N__25013\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__25016\,
            I => \N__25010\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__25013\,
            I => \N__25007\
        );

    \I__5246\ : Span4Mux_h
    port map (
            O => \N__25010\,
            I => \N__25002\
        );

    \I__5245\ : Span4Mux_v
    port map (
            O => \N__25007\,
            I => \N__25002\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__25002\,
            I => \c0.n8855\
        );

    \I__5243\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24996\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__5241\ : Span12Mux_s3_v
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__5240\ : Odrv12
    port map (
            O => \N__24990\,
            I => \c0.n35\
        );

    \I__5239\ : CascadeMux
    port map (
            O => \N__24987\,
            I => \N__24981\
        );

    \I__5238\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24975\
        );

    \I__5237\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24975\
        );

    \I__5236\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24970\
        );

    \I__5235\ : InMux
    port map (
            O => \N__24981\,
            I => \N__24970\
        );

    \I__5234\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24967\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__24975\,
            I => data_in_field_84
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__24970\,
            I => data_in_field_84
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__24967\,
            I => data_in_field_84
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__24960\,
            I => \N__24955\
        );

    \I__5229\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24952\
        );

    \I__5228\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24949\
        );

    \I__5227\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24945\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__24952\,
            I => \N__24938\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__24949\,
            I => \N__24938\
        );

    \I__5224\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24935\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__24945\,
            I => \N__24932\
        );

    \I__5222\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24929\
        );

    \I__5221\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24926\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__24938\,
            I => \N__24923\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__24935\,
            I => \N__24918\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__24932\,
            I => \N__24918\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__24929\,
            I => data_in_field_92
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__24926\,
            I => data_in_field_92
        );

    \I__5215\ : Odrv4
    port map (
            O => \N__24923\,
            I => data_in_field_92
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__24918\,
            I => data_in_field_92
        );

    \I__5213\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__24906\,
            I => \c0.n9560\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24899\
        );

    \I__5210\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24896\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__24899\,
            I => \N__24893\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__24896\,
            I => \N__24890\
        );

    \I__5207\ : Span4Mux_h
    port map (
            O => \N__24893\,
            I => \N__24882\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__24890\,
            I => \N__24882\
        );

    \I__5205\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24877\
        );

    \I__5204\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24877\
        );

    \I__5203\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24874\
        );

    \I__5202\ : Span4Mux_v
    port map (
            O => \N__24882\,
            I => \N__24871\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24868\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__24874\,
            I => data_in_field_108
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__24871\,
            I => data_in_field_108
        );

    \I__5198\ : Odrv12
    port map (
            O => \N__24868\,
            I => data_in_field_108
        );

    \I__5197\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24857\
        );

    \I__5196\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24853\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__24857\,
            I => \N__24850\
        );

    \I__5194\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24847\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__24853\,
            I => \N__24842\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__24850\,
            I => \N__24839\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24836\
        );

    \I__5190\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24833\
        );

    \I__5189\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24830\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__24842\,
            I => \N__24827\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__24839\,
            I => \N__24820\
        );

    \I__5186\ : Span4Mux_v
    port map (
            O => \N__24836\,
            I => \N__24820\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24820\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__24830\,
            I => data_in_field_100
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__24827\,
            I => data_in_field_100
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__24820\,
            I => data_in_field_100
        );

    \I__5181\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24810\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__5179\ : Span12Mux_h
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__5178\ : Odrv12
    port map (
            O => \N__24804\,
            I => \c0.n8927\
        );

    \I__5177\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24795\
        );

    \I__5176\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24795\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__5174\ : Odrv12
    port map (
            O => \N__24792\,
            I => \c0.n8837\
        );

    \I__5173\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24782\
        );

    \I__5171\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24777\
        );

    \I__5170\ : Span4Mux_v
    port map (
            O => \N__24782\,
            I => \N__24773\
        );

    \I__5169\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24770\
        );

    \I__5168\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24767\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__24777\,
            I => \N__24764\
        );

    \I__5166\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24761\
        );

    \I__5165\ : Span4Mux_h
    port map (
            O => \N__24773\,
            I => \N__24756\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24756\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24751\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__24764\,
            I => \N__24748\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24743\
        );

    \I__5160\ : Span4Mux_v
    port map (
            O => \N__24756\,
            I => \N__24743\
        );

    \I__5159\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24738\
        );

    \I__5158\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24738\
        );

    \I__5157\ : Odrv12
    port map (
            O => \N__24751\,
            I => data_in_field_41
        );

    \I__5156\ : Odrv4
    port map (
            O => \N__24748\,
            I => data_in_field_41
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__24743\,
            I => data_in_field_41
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__24738\,
            I => data_in_field_41
        );

    \I__5153\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24726\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__24723\,
            I => \c0.n16_adj_1629\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__24720\,
            I => \N__24717\
        );

    \I__5149\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24710\
        );

    \I__5147\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24707\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__24710\,
            I => \N__24704\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24701\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__24704\,
            I => \N__24698\
        );

    \I__5143\ : Span4Mux_s3_v
    port map (
            O => \N__24701\,
            I => \N__24695\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__24698\,
            I => \c0.n8977\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__24695\,
            I => \c0.n8977\
        );

    \I__5140\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__24687\,
            I => \c0.n17_adj_1630\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__5137\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24678\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__24678\,
            I => \c0.data_in_frame_19_4\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__24675\,
            I => \N__24672\
        );

    \I__5134\ : InMux
    port map (
            O => \N__24672\,
            I => \N__24669\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__5132\ : Span4Mux_s3_v
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__24663\,
            I => \N__24660\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__24660\,
            I => \c0.data_in_frame_20_4\
        );

    \I__5129\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24651\
        );

    \I__5128\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24648\
        );

    \I__5127\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24645\
        );

    \I__5126\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24642\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24639\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24636\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__24645\,
            I => \N__24633\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__24642\,
            I => \N__24630\
        );

    \I__5121\ : Span4Mux_v
    port map (
            O => \N__24639\,
            I => \N__24626\
        );

    \I__5120\ : Span4Mux_h
    port map (
            O => \N__24636\,
            I => \N__24623\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__24633\,
            I => \N__24618\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__24630\,
            I => \N__24618\
        );

    \I__5117\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24615\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__24626\,
            I => rand_data_6
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__24623\,
            I => rand_data_6
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__24618\,
            I => rand_data_6
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__24615\,
            I => rand_data_6
        );

    \I__5112\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24601\
        );

    \I__5111\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24598\
        );

    \I__5110\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24595\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__24601\,
            I => \N__24590\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__24598\,
            I => \N__24590\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__24595\,
            I => \N__24587\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__24590\,
            I => \N__24584\
        );

    \I__5105\ : Span4Mux_s1_v
    port map (
            O => \N__24587\,
            I => \N__24581\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__24584\,
            I => \N__24576\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__24581\,
            I => \N__24573\
        );

    \I__5102\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24568\
        );

    \I__5101\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24568\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__24576\,
            I => data_in_field_102
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__24573\,
            I => data_in_field_102
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__24568\,
            I => data_in_field_102
        );

    \I__5097\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24556\
        );

    \I__5096\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24553\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__24559\,
            I => \N__24550\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__24556\,
            I => \N__24546\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__24553\,
            I => \N__24543\
        );

    \I__5092\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24540\
        );

    \I__5091\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24536\
        );

    \I__5090\ : Span4Mux_v
    port map (
            O => \N__24546\,
            I => \N__24533\
        );

    \I__5089\ : Span4Mux_s2_h
    port map (
            O => \N__24543\,
            I => \N__24530\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__24540\,
            I => \N__24527\
        );

    \I__5087\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24524\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24521\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__24533\,
            I => \N__24518\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__24530\,
            I => \N__24513\
        );

    \I__5083\ : Span4Mux_s2_v
    port map (
            O => \N__24527\,
            I => \N__24513\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__24524\,
            I => data_in_field_125
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__24521\,
            I => data_in_field_125
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__24518\,
            I => data_in_field_125
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__24513\,
            I => data_in_field_125
        );

    \I__5078\ : InMux
    port map (
            O => \N__24504\,
            I => \N__24500\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__24503\,
            I => \N__24497\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__24500\,
            I => \N__24494\
        );

    \I__5075\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24491\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__24494\,
            I => \N__24485\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24482\
        );

    \I__5072\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24479\
        );

    \I__5071\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24476\
        );

    \I__5070\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24473\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__24485\,
            I => \N__24466\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__24482\,
            I => \N__24466\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24466\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__24476\,
            I => data_in_field_73
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__24473\,
            I => data_in_field_73
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__24466\,
            I => data_in_field_73
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__5062\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24453\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__24453\,
            I => \c0.n18_adj_1618\
        );

    \I__5060\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24446\
        );

    \I__5059\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24443\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__24446\,
            I => \N__24438\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24434\
        );

    \I__5056\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24429\
        );

    \I__5055\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24429\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__24438\,
            I => \N__24426\
        );

    \I__5053\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24423\
        );

    \I__5052\ : Span4Mux_h
    port map (
            O => \N__24434\,
            I => \N__24420\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__24429\,
            I => \N__24417\
        );

    \I__5050\ : Span4Mux_v
    port map (
            O => \N__24426\,
            I => \N__24414\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__24423\,
            I => \N__24407\
        );

    \I__5048\ : Span4Mux_v
    port map (
            O => \N__24420\,
            I => \N__24407\
        );

    \I__5047\ : Span4Mux_v
    port map (
            O => \N__24417\,
            I => \N__24407\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__24414\,
            I => data_in_field_54
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__24407\,
            I => data_in_field_54
        );

    \I__5044\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24399\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__24399\,
            I => \N__24395\
        );

    \I__5042\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24392\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__24395\,
            I => \N__24387\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__24392\,
            I => \N__24384\
        );

    \I__5039\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24379\
        );

    \I__5038\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24379\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__24387\,
            I => data_in_field_69
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__24384\,
            I => data_in_field_69
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__24379\,
            I => data_in_field_69
        );

    \I__5034\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24369\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24366\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__24366\,
            I => \N__24362\
        );

    \I__5031\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24359\
        );

    \I__5030\ : Span4Mux_h
    port map (
            O => \N__24362\,
            I => \N__24354\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24354\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__24354\,
            I => \c0.n8998\
        );

    \I__5027\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24348\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__5025\ : Span4Mux_s3_h
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__5024\ : Span4Mux_h
    port map (
            O => \N__24342\,
            I => \N__24339\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__24339\,
            I => \c0.n16_adj_1591\
        );

    \I__5022\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24328\
        );

    \I__5020\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24323\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24323\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__24328\,
            I => \N__24320\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24317\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__24320\,
            I => \N__24314\
        );

    \I__5015\ : Span4Mux_v
    port map (
            O => \N__24317\,
            I => \N__24308\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__24314\,
            I => \N__24308\
        );

    \I__5013\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24305\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__24308\,
            I => rand_data_20
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__24305\,
            I => rand_data_20
        );

    \I__5010\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24293\
        );

    \I__5009\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24293\
        );

    \I__5008\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24288\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__24293\,
            I => \N__24285\
        );

    \I__5006\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24282\
        );

    \I__5005\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24278\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__24288\,
            I => \N__24273\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__24285\,
            I => \N__24273\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24270\
        );

    \I__5001\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24267\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__24278\,
            I => \N__24264\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__24273\,
            I => \N__24261\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__24270\,
            I => \N__24258\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__24267\,
            I => data_in_field_124
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__24264\,
            I => data_in_field_124
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__24261\,
            I => data_in_field_124
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__24258\,
            I => data_in_field_124
        );

    \I__4993\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__24243\,
            I => \N__24237\
        );

    \I__4990\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24230\
        );

    \I__4989\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24230\
        );

    \I__4988\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24230\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__24237\,
            I => data_in_field_116
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__24230\,
            I => data_in_field_116
        );

    \I__4985\ : InMux
    port map (
            O => \N__24225\,
            I => \N__24220\
        );

    \I__4984\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24217\
        );

    \I__4983\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24214\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__24220\,
            I => \N__24208\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__24217\,
            I => \N__24208\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24205\
        );

    \I__4979\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24202\
        );

    \I__4978\ : Span4Mux_v
    port map (
            O => \N__24208\,
            I => \N__24199\
        );

    \I__4977\ : Span4Mux_v
    port map (
            O => \N__24205\,
            I => \N__24196\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__24202\,
            I => data_in_field_56
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__24199\,
            I => data_in_field_56
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__24196\,
            I => data_in_field_56
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__24189\,
            I => \N__24185\
        );

    \I__4972\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24180\
        );

    \I__4971\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24177\
        );

    \I__4970\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24174\
        );

    \I__4969\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24171\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__24180\,
            I => \N__24168\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__24177\,
            I => \N__24165\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24162\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__24171\,
            I => \N__24159\
        );

    \I__4964\ : Span4Mux_s2_v
    port map (
            O => \N__24168\,
            I => \N__24155\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__24165\,
            I => \N__24150\
        );

    \I__4962\ : Span4Mux_v
    port map (
            O => \N__24162\,
            I => \N__24150\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__24159\,
            I => \N__24147\
        );

    \I__4960\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24144\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__24155\,
            I => \N__24141\
        );

    \I__4958\ : Span4Mux_h
    port map (
            O => \N__24150\,
            I => \N__24136\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__24147\,
            I => \N__24136\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__24144\,
            I => data_in_field_101
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__24141\,
            I => data_in_field_101
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__24136\,
            I => data_in_field_101
        );

    \I__4953\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24124\
        );

    \I__4952\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24121\
        );

    \I__4951\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24118\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__24124\,
            I => \N__24113\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24113\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__24118\,
            I => \N__24110\
        );

    \I__4947\ : Span4Mux_v
    port map (
            O => \N__24113\,
            I => \N__24107\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__24110\,
            I => \N__24103\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__24107\,
            I => \N__24100\
        );

    \I__4944\ : InMux
    port map (
            O => \N__24106\,
            I => \N__24097\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__24103\,
            I => rand_data_16
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__24100\,
            I => rand_data_16
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__24097\,
            I => rand_data_16
        );

    \I__4940\ : InMux
    port map (
            O => \N__24090\,
            I => \N__24086\
        );

    \I__4939\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24083\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__24086\,
            I => \N__24077\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__24083\,
            I => \N__24077\
        );

    \I__4936\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24074\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__24077\,
            I => \N__24071\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24067\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__24071\,
            I => \N__24064\
        );

    \I__4932\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24061\
        );

    \I__4931\ : Span12Mux_h
    port map (
            O => \N__24067\,
            I => \N__24058\
        );

    \I__4930\ : Span4Mux_s2_v
    port map (
            O => \N__24064\,
            I => \N__24055\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__24061\,
            I => rand_data_26
        );

    \I__4928\ : Odrv12
    port map (
            O => \N__24058\,
            I => rand_data_26
        );

    \I__4927\ : Odrv4
    port map (
            O => \N__24055\,
            I => rand_data_26
        );

    \I__4926\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24044\
        );

    \I__4925\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24041\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__24037\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24034\
        );

    \I__4922\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24030\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__24037\,
            I => \N__24027\
        );

    \I__4920\ : Sp12to4
    port map (
            O => \N__24034\,
            I => \N__24024\
        );

    \I__4919\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24021\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__24030\,
            I => data_in_field_58
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__24027\,
            I => data_in_field_58
        );

    \I__4916\ : Odrv12
    port map (
            O => \N__24024\,
            I => data_in_field_58
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__24021\,
            I => data_in_field_58
        );

    \I__4914\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24007\
        );

    \I__4913\ : InMux
    port map (
            O => \N__24011\,
            I => \N__24004\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__24010\,
            I => \N__24000\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__24007\,
            I => \N__23997\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__24004\,
            I => \N__23994\
        );

    \I__4909\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23991\
        );

    \I__4908\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23988\
        );

    \I__4907\ : Span4Mux_h
    port map (
            O => \N__23997\,
            I => \N__23985\
        );

    \I__4906\ : Span12Mux_s1_v
    port map (
            O => \N__23994\,
            I => \N__23980\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23980\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__23988\,
            I => data_in_field_118
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__23985\,
            I => data_in_field_118
        );

    \I__4902\ : Odrv12
    port map (
            O => \N__23980\,
            I => data_in_field_118
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__23973\,
            I => \N__23970\
        );

    \I__4900\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23967\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__23967\,
            I => \c0.n4534\
        );

    \I__4898\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__23961\,
            I => \N__23958\
        );

    \I__4896\ : Span4Mux_h
    port map (
            O => \N__23958\,
            I => \N__23955\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__23955\,
            I => \c0.n27_adj_1621\
        );

    \I__4894\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23948\
        );

    \I__4893\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23945\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23938\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23938\
        );

    \I__4890\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23933\
        );

    \I__4889\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23933\
        );

    \I__4888\ : Span12Mux_h
    port map (
            O => \N__23938\,
            I => \N__23929\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__23933\,
            I => \N__23926\
        );

    \I__4886\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23923\
        );

    \I__4885\ : Odrv12
    port map (
            O => \N__23929\,
            I => rand_data_10
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__23926\,
            I => rand_data_10
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__23923\,
            I => rand_data_10
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__23916\,
            I => \N__23913\
        );

    \I__4881\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23910\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23907\
        );

    \I__4879\ : Span12Mux_s5_v
    port map (
            O => \N__23907\,
            I => \N__23904\
        );

    \I__4878\ : Odrv12
    port map (
            O => \N__23904\,
            I => \c0.n4473\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__23901\,
            I => \c0.n4473_cascade_\
        );

    \I__4876\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23895\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__23895\,
            I => \N__23891\
        );

    \I__4874\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23888\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__23891\,
            I => \N__23885\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__23888\,
            I => \c0.n9010\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__23885\,
            I => \c0.n9010\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__23880\,
            I => \c0.n4244_cascade_\
        );

    \I__4869\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23874\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23871\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__4866\ : Span4Mux_h
    port map (
            O => \N__23868\,
            I => \N__23865\
        );

    \I__4865\ : Odrv4
    port map (
            O => \N__23865\,
            I => \c0.n4479\
        );

    \I__4864\ : CascadeMux
    port map (
            O => \N__23862\,
            I => \c0.n4235_cascade_\
        );

    \I__4863\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__23856\,
            I => \c0.n4562\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__23853\,
            I => \N__23846\
        );

    \I__4860\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23842\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23839\
        );

    \I__4858\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23834\
        );

    \I__4857\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23834\
        );

    \I__4856\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23831\
        );

    \I__4855\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23828\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__23842\,
            I => \N__23825\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23821\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23818\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__23831\,
            I => \N__23815\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__23828\,
            I => \N__23810\
        );

    \I__4849\ : Span4Mux_s3_h
    port map (
            O => \N__23825\,
            I => \N__23810\
        );

    \I__4848\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23807\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__23821\,
            I => \N__23804\
        );

    \I__4846\ : Span4Mux_h
    port map (
            O => \N__23818\,
            I => \N__23799\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__23815\,
            I => \N__23799\
        );

    \I__4844\ : Span4Mux_v
    port map (
            O => \N__23810\,
            I => \N__23796\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__23807\,
            I => data_in_field_99
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__23804\,
            I => data_in_field_99
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__23799\,
            I => data_in_field_99
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__23796\,
            I => data_in_field_99
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__23787\,
            I => \N__23783\
        );

    \I__4838\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23776\
        );

    \I__4837\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23776\
        );

    \I__4836\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23772\
        );

    \I__4835\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23769\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__23776\,
            I => \N__23766\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__23775\,
            I => \N__23763\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23759\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23756\
        );

    \I__4830\ : Span4Mux_v
    port map (
            O => \N__23766\,
            I => \N__23753\
        );

    \I__4829\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23748\
        );

    \I__4828\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23748\
        );

    \I__4827\ : Span4Mux_s3_h
    port map (
            O => \N__23759\,
            I => \N__23745\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__23756\,
            I => \N__23740\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__23753\,
            I => \N__23740\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__23748\,
            I => data_in_field_131
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__23745\,
            I => data_in_field_131
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__23740\,
            I => data_in_field_131
        );

    \I__4821\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__4819\ : Span4Mux_h
    port map (
            O => \N__23727\,
            I => \N__23724\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__23724\,
            I => \c0.n8846\
        );

    \I__4817\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23715\
        );

    \I__4816\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23715\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23711\
        );

    \I__4814\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23708\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__23711\,
            I => \N__23703\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23700\
        );

    \I__4811\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23697\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23694\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__23703\,
            I => rand_data_2
        );

    \I__4808\ : Odrv12
    port map (
            O => \N__23700\,
            I => rand_data_2
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__23697\,
            I => rand_data_2
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__23694\,
            I => rand_data_2
        );

    \I__4805\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__4803\ : Odrv12
    port map (
            O => \N__23679\,
            I => \c0.n30\
        );

    \I__4802\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__4800\ : Span4Mux_v
    port map (
            O => \N__23670\,
            I => \N__23664\
        );

    \I__4799\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23656\
        );

    \I__4798\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23653\
        );

    \I__4797\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23650\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__23664\,
            I => \N__23647\
        );

    \I__4795\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23640\
        );

    \I__4794\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23640\
        );

    \I__4793\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23640\
        );

    \I__4792\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23635\
        );

    \I__4791\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23635\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__23656\,
            I => \N__23630\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__23653\,
            I => \N__23630\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23623\
        );

    \I__4787\ : Span4Mux_h
    port map (
            O => \N__23647\,
            I => \N__23623\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23623\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__23635\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__4784\ : Odrv12
    port map (
            O => \N__23630\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__23623\,
            I => \FRAME_MATCHER_state_2\
        );

    \I__4782\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__4780\ : Span4Mux_s2_h
    port map (
            O => \N__23610\,
            I => \N__23606\
        );

    \I__4779\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23603\
        );

    \I__4778\ : Span4Mux_h
    port map (
            O => \N__23606\,
            I => \N__23600\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23597\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__23600\,
            I => \N__23594\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__23597\,
            I => \c0.n7194\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__23594\,
            I => \c0.n7194\
        );

    \I__4773\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23586\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__23583\,
            I => \N__23580\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__23580\,
            I => n9262
        );

    \I__4769\ : InMux
    port map (
            O => \N__23577\,
            I => \N__23568\
        );

    \I__4768\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23568\
        );

    \I__4767\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23568\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__23568\,
            I => data_in_6_2
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__23565\,
            I => \N__23555\
        );

    \I__4764\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23537\
        );

    \I__4763\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23528\
        );

    \I__4762\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23528\
        );

    \I__4761\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23528\
        );

    \I__4760\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23528\
        );

    \I__4759\ : CascadeMux
    port map (
            O => \N__23559\,
            I => \N__23521\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__23558\,
            I => \N__23517\
        );

    \I__4757\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23509\
        );

    \I__4756\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23509\
        );

    \I__4755\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23509\
        );

    \I__4754\ : CascadeMux
    port map (
            O => \N__23552\,
            I => \N__23503\
        );

    \I__4753\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23494\
        );

    \I__4752\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23494\
        );

    \I__4751\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23494\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__23548\,
            I => \N__23490\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__23547\,
            I => \N__23487\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__23546\,
            I => \N__23474\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23465\
        );

    \I__4746\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23460\
        );

    \I__4745\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23460\
        );

    \I__4744\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23457\
        );

    \I__4743\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23452\
        );

    \I__4742\ : InMux
    port map (
            O => \N__23540\,
            I => \N__23452\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__23537\,
            I => \N__23448\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__23528\,
            I => \N__23445\
        );

    \I__4739\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23438\
        );

    \I__4738\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23438\
        );

    \I__4737\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23438\
        );

    \I__4736\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23433\
        );

    \I__4735\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23433\
        );

    \I__4734\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23430\
        );

    \I__4733\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23424\
        );

    \I__4732\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23424\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__23509\,
            I => \N__23421\
        );

    \I__4730\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23415\
        );

    \I__4729\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23410\
        );

    \I__4728\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23410\
        );

    \I__4727\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23403\
        );

    \I__4726\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23403\
        );

    \I__4725\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23403\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__23494\,
            I => \N__23397\
        );

    \I__4723\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23386\
        );

    \I__4722\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23386\
        );

    \I__4721\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23386\
        );

    \I__4720\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23386\
        );

    \I__4719\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23386\
        );

    \I__4718\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23383\
        );

    \I__4717\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23372\
        );

    \I__4716\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23372\
        );

    \I__4715\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23372\
        );

    \I__4714\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23372\
        );

    \I__4713\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23372\
        );

    \I__4712\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23361\
        );

    \I__4711\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23361\
        );

    \I__4710\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23361\
        );

    \I__4709\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23361\
        );

    \I__4708\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23361\
        );

    \I__4707\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23350\
        );

    \I__4706\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23350\
        );

    \I__4705\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23350\
        );

    \I__4704\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23350\
        );

    \I__4703\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23350\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23345\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23345\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23342\
        );

    \I__4699\ : InMux
    port map (
            O => \N__23451\,
            I => \N__23339\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__23448\,
            I => \N__23332\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__23445\,
            I => \N__23332\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23332\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__23433\,
            I => \N__23327\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__23430\,
            I => \N__23327\
        );

    \I__4693\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23322\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__23424\,
            I => \N__23319\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__23421\,
            I => \N__23316\
        );

    \I__4690\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23313\
        );

    \I__4689\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23308\
        );

    \I__4688\ : InMux
    port map (
            O => \N__23418\,
            I => \N__23308\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__23415\,
            I => \N__23301\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__23410\,
            I => \N__23301\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23301\
        );

    \I__4684\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23294\
        );

    \I__4683\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23294\
        );

    \I__4682\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23294\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__23397\,
            I => \N__23291\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__23386\,
            I => \N__23286\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23286\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23275\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__23361\,
            I => \N__23275\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__23350\,
            I => \N__23275\
        );

    \I__4675\ : Span4Mux_h
    port map (
            O => \N__23345\,
            I => \N__23275\
        );

    \I__4674\ : Span4Mux_v
    port map (
            O => \N__23342\,
            I => \N__23275\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23268\
        );

    \I__4672\ : Span4Mux_v
    port map (
            O => \N__23332\,
            I => \N__23268\
        );

    \I__4671\ : Span4Mux_v
    port map (
            O => \N__23327\,
            I => \N__23268\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__23326\,
            I => \N__23263\
        );

    \I__4669\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23259\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23248\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__23319\,
            I => \N__23248\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__23316\,
            I => \N__23248\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23248\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__23308\,
            I => \N__23248\
        );

    \I__4663\ : Span4Mux_v
    port map (
            O => \N__23301\,
            I => \N__23241\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__23294\,
            I => \N__23241\
        );

    \I__4661\ : Span4Mux_h
    port map (
            O => \N__23291\,
            I => \N__23241\
        );

    \I__4660\ : Span4Mux_s3_h
    port map (
            O => \N__23286\,
            I => \N__23234\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__23275\,
            I => \N__23234\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__23268\,
            I => \N__23234\
        );

    \I__4657\ : InMux
    port map (
            O => \N__23267\,
            I => \N__23229\
        );

    \I__4656\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23229\
        );

    \I__4655\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23224\
        );

    \I__4654\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23224\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__23259\,
            I => \N__23219\
        );

    \I__4652\ : Sp12to4
    port map (
            O => \N__23248\,
            I => \N__23219\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__23241\,
            I => \N__23216\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__23234\,
            I => \N__23213\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__23229\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__23224\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__4647\ : Odrv12
    port map (
            O => \N__23219\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__4646\ : Odrv4
    port map (
            O => \N__23216\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__23213\,
            I => \FRAME_MATCHER_state_0\
        );

    \I__4644\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23196\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__23196\,
            I => \N__23193\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__23193\,
            I => n1893
        );

    \I__4640\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23184\
        );

    \I__4639\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23184\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__23184\,
            I => data_in_7_2
        );

    \I__4637\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23175\
        );

    \I__4636\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23175\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__23175\,
            I => data_in_8_2
        );

    \I__4634\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23169\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__23169\,
            I => \N__23166\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__23166\,
            I => \N__23162\
        );

    \I__4631\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23159\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__23162\,
            I => data_in_10_2
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__23159\,
            I => data_in_10_2
        );

    \I__4628\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23148\
        );

    \I__4627\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23148\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__23148\,
            I => data_in_9_2
        );

    \I__4625\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23141\
        );

    \I__4624\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23138\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23135\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__23138\,
            I => \N__23132\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__23135\,
            I => \N__23129\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__23132\,
            I => \N__23126\
        );

    \I__4619\ : Sp12to4
    port map (
            O => \N__23129\,
            I => \N__23121\
        );

    \I__4618\ : Sp12to4
    port map (
            O => \N__23126\,
            I => \N__23121\
        );

    \I__4617\ : Odrv12
    port map (
            O => \N__23121\,
            I => \c0.n8921\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__23118\,
            I => \c0.n4562_cascade_\
        );

    \I__4615\ : InMux
    port map (
            O => \N__23115\,
            I => \N__23109\
        );

    \I__4614\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23109\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__23109\,
            I => data_in_16_2
        );

    \I__4612\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23100\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23100\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__23100\,
            I => data_in_18_2
        );

    \I__4609\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23093\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23090\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__23093\,
            I => data_in_17_2
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__23090\,
            I => data_in_17_2
        );

    \I__4605\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23082\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__23082\,
            I => \N__23079\
        );

    \I__4603\ : Span4Mux_h
    port map (
            O => \N__23079\,
            I => \N__23075\
        );

    \I__4602\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23072\
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__23075\,
            I => data_in_20_2
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__23072\,
            I => data_in_20_2
        );

    \I__4599\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23061\
        );

    \I__4598\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23061\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__23061\,
            I => data_in_19_2
        );

    \I__4596\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23052\
        );

    \I__4595\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23052\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23049\
        );

    \I__4593\ : Span4Mux_h
    port map (
            O => \N__23049\,
            I => \N__23046\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__23046\,
            I => n7171
        );

    \I__4591\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23040\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__23037\,
            I => \c0.n9668\
        );

    \I__4588\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__4586\ : Span12Mux_h
    port map (
            O => \N__23028\,
            I => \N__23024\
        );

    \I__4585\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23021\
        );

    \I__4584\ : Odrv12
    port map (
            O => \N__23024\,
            I => \c0.n8878\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__23021\,
            I => \c0.n8878\
        );

    \I__4582\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23013\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__23013\,
            I => \N__23009\
        );

    \I__4580\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23006\
        );

    \I__4579\ : Span4Mux_h
    port map (
            O => \N__23009\,
            I => \N__23003\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__23000\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__23003\,
            I => \c0.n8813\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__23000\,
            I => \c0.n8813\
        );

    \I__4575\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22992\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__22992\,
            I => \N__22988\
        );

    \I__4573\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22985\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__22988\,
            I => \N__22978\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22978\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__22984\,
            I => \N__22973\
        );

    \I__4569\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22969\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__22978\,
            I => \N__22966\
        );

    \I__4567\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22957\
        );

    \I__4566\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22957\
        );

    \I__4565\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22957\
        );

    \I__4564\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22957\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__22969\,
            I => data_in_field_43
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__22966\,
            I => data_in_field_43
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__22957\,
            I => data_in_field_43
        );

    \I__4560\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22944\
        );

    \I__4558\ : Span4Mux_v
    port map (
            O => \N__22944\,
            I => \N__22941\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__22941\,
            I => \c0.n28_adj_1619\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__22938\,
            I => \c0.n29_adj_1620_cascade_\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__22935\,
            I => \N__22932\
        );

    \I__4554\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22929\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__4552\ : Odrv12
    port map (
            O => \N__22926\,
            I => \c0.data_in_frame_19_6\
        );

    \I__4551\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22920\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__22920\,
            I => \N__22917\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__22917\,
            I => \N__22914\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__22914\,
            I => n1901
        );

    \I__4547\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__22908\,
            I => \c0.n9141\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__22905\,
            I => \c0.n9138_cascade_\
        );

    \I__4544\ : InMux
    port map (
            O => \N__22902\,
            I => \N__22899\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__22896\,
            I => \N__22893\
        );

    \I__4541\ : Span4Mux_v
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__4540\ : Span4Mux_v
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__4539\ : Odrv4
    port map (
            O => \N__22887\,
            I => \c0.n9132\
        );

    \I__4538\ : InMux
    port map (
            O => \N__22884\,
            I => \N__22881\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__22881\,
            I => \c0.n9135\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__22878\,
            I => \c0.n9614_cascade_\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \c0.n9617_cascade_\
        );

    \I__4534\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__22866\,
            I => \c0.tx2.r_Tx_Data_6\
        );

    \I__4531\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22857\
        );

    \I__4530\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22857\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__22857\,
            I => data_in_11_2
        );

    \I__4528\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22848\
        );

    \I__4527\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22848\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__22848\,
            I => data_in_12_2
        );

    \I__4525\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22839\
        );

    \I__4524\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22839\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__22839\,
            I => data_in_13_2
        );

    \I__4522\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22830\
        );

    \I__4521\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22830\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__22830\,
            I => data_in_14_2
        );

    \I__4519\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22821\
        );

    \I__4518\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22821\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__22821\,
            I => data_in_15_2
        );

    \I__4516\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__4514\ : Odrv12
    port map (
            O => \N__22812\,
            I => \c0.n18_adj_1666\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__22809\,
            I => \N__22806\
        );

    \I__4512\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22801\
        );

    \I__4511\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22798\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__22804\,
            I => \N__22795\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__22801\,
            I => \N__22792\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__22798\,
            I => \N__22789\
        );

    \I__4507\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22786\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__22792\,
            I => \N__22783\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__22789\,
            I => \N__22780\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__22786\,
            I => \N__22774\
        );

    \I__4503\ : Span4Mux_v
    port map (
            O => \N__22783\,
            I => \N__22771\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__22780\,
            I => \N__22768\
        );

    \I__4501\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22765\
        );

    \I__4500\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22760\
        );

    \I__4499\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22760\
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__22774\,
            I => data_in_field_36
        );

    \I__4497\ : Odrv4
    port map (
            O => \N__22771\,
            I => data_in_field_36
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__22768\,
            I => data_in_field_36
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__22765\,
            I => data_in_field_36
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__22760\,
            I => data_in_field_36
        );

    \I__4493\ : InMux
    port map (
            O => \N__22749\,
            I => \N__22746\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__22740\,
            I => \c0.n1645\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__22737\,
            I => \N__22733\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__22736\,
            I => \N__22730\
        );

    \I__4487\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22725\
        );

    \I__4486\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22722\
        );

    \I__4485\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22719\
        );

    \I__4484\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22716\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__22725\,
            I => \N__22710\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__22722\,
            I => \N__22710\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__22719\,
            I => \N__22707\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22704\
        );

    \I__4479\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22701\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__22710\,
            I => \N__22698\
        );

    \I__4477\ : Span4Mux_s2_v
    port map (
            O => \N__22707\,
            I => \N__22693\
        );

    \I__4476\ : Span4Mux_h
    port map (
            O => \N__22704\,
            I => \N__22693\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__22701\,
            I => data_in_field_62
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__22698\,
            I => data_in_field_62
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__22693\,
            I => data_in_field_62
        );

    \I__4472\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22682\
        );

    \I__4471\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22679\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__22682\,
            I => \N__22676\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22668\
        );

    \I__4468\ : Span4Mux_h
    port map (
            O => \N__22676\,
            I => \N__22665\
        );

    \I__4467\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22662\
        );

    \I__4466\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22657\
        );

    \I__4465\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22657\
        );

    \I__4464\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22654\
        );

    \I__4463\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22651\
        );

    \I__4462\ : Span4Mux_v
    port map (
            O => \N__22668\,
            I => \N__22648\
        );

    \I__4461\ : Span4Mux_v
    port map (
            O => \N__22665\,
            I => \N__22643\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__22662\,
            I => \N__22643\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__22657\,
            I => \N__22640\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22637\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__22651\,
            I => data_in_field_46
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__22648\,
            I => data_in_field_46
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__22643\,
            I => data_in_field_46
        );

    \I__4454\ : Odrv12
    port map (
            O => \N__22640\,
            I => data_in_field_46
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__22637\,
            I => data_in_field_46
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__22626\,
            I => \c0.n9632_cascade_\
        );

    \I__4451\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22620\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__22620\,
            I => \N__22616\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \N__22611\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__22616\,
            I => \N__22608\
        );

    \I__4447\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22605\
        );

    \I__4446\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22601\
        );

    \I__4445\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22598\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__22608\,
            I => \N__22595\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__22605\,
            I => \N__22592\
        );

    \I__4442\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22589\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22586\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__22598\,
            I => \c0.data_in_field_38\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__22595\,
            I => \c0.data_in_field_38\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__22592\,
            I => \c0.data_in_field_38\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__22589\,
            I => \c0.data_in_field_38\
        );

    \I__4436\ : Odrv12
    port map (
            O => \N__22586\,
            I => \c0.data_in_field_38\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__22575\,
            I => \N__22571\
        );

    \I__4434\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22567\
        );

    \I__4433\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22564\
        );

    \I__4432\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22559\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__22567\,
            I => \N__22554\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__22564\,
            I => \N__22554\
        );

    \I__4429\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22549\
        );

    \I__4428\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22549\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22546\
        );

    \I__4426\ : Span12Mux_s4_v
    port map (
            O => \N__22554\,
            I => \N__22543\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__22549\,
            I => data_in_field_126
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__22546\,
            I => data_in_field_126
        );

    \I__4423\ : Odrv12
    port map (
            O => \N__22543\,
            I => data_in_field_126
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__22536\,
            I => \c0.n9620_cascade_\
        );

    \I__4421\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22528\
        );

    \I__4420\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22525\
        );

    \I__4419\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22520\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22517\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__22525\,
            I => \N__22513\
        );

    \I__4416\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22510\
        );

    \I__4415\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22507\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22502\
        );

    \I__4413\ : Span4Mux_s2_v
    port map (
            O => \N__22517\,
            I => \N__22502\
        );

    \I__4412\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22499\
        );

    \I__4411\ : Span4Mux_v
    port map (
            O => \N__22513\,
            I => \N__22494\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__22510\,
            I => \N__22494\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__22507\,
            I => \N__22489\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__22502\,
            I => \N__22489\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22484\
        );

    \I__4406\ : Span4Mux_h
    port map (
            O => \N__22494\,
            I => \N__22484\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__22489\,
            I => data_in_field_94
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__22484\,
            I => data_in_field_94
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__22479\,
            I => \c0.n9626_cascade_\
        );

    \I__4402\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22472\
        );

    \I__4401\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22469\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22464\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__22469\,
            I => \N__22460\
        );

    \I__4398\ : InMux
    port map (
            O => \N__22468\,
            I => \N__22457\
        );

    \I__4397\ : InMux
    port map (
            O => \N__22467\,
            I => \N__22454\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__22464\,
            I => \N__22451\
        );

    \I__4395\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22448\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__22460\,
            I => \N__22443\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__22457\,
            I => \N__22443\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22438\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__22451\,
            I => \N__22438\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__22448\,
            I => data_in_field_44
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__22443\,
            I => data_in_field_44
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__22438\,
            I => data_in_field_44
        );

    \I__4387\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__4385\ : Odrv12
    port map (
            O => \N__22425\,
            I => \c0.n9572\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__4383\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22415\
        );

    \I__4382\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22412\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22408\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__22412\,
            I => \N__22404\
        );

    \I__4379\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22401\
        );

    \I__4378\ : Span12Mux_s6_v
    port map (
            O => \N__22408\,
            I => \N__22398\
        );

    \I__4377\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22395\
        );

    \I__4376\ : Span4Mux_s3_v
    port map (
            O => \N__22404\,
            I => \N__22392\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__22401\,
            I => data_in_field_77
        );

    \I__4374\ : Odrv12
    port map (
            O => \N__22398\,
            I => data_in_field_77
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__22395\,
            I => data_in_field_77
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__22392\,
            I => data_in_field_77
        );

    \I__4371\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22379\
        );

    \I__4370\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22376\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22372\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22369\
        );

    \I__4367\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22365\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__22372\,
            I => \N__22362\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__22369\,
            I => \N__22359\
        );

    \I__4364\ : InMux
    port map (
            O => \N__22368\,
            I => \N__22355\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__22365\,
            I => \N__22352\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__22362\,
            I => \N__22349\
        );

    \I__4361\ : Span4Mux_h
    port map (
            O => \N__22359\,
            I => \N__22346\
        );

    \I__4360\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22343\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__22355\,
            I => data_in_field_49
        );

    \I__4358\ : Odrv12
    port map (
            O => \N__22352\,
            I => data_in_field_49
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__22349\,
            I => data_in_field_49
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__22346\,
            I => data_in_field_49
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__22343\,
            I => data_in_field_49
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__22332\,
            I => \c0.n8887_cascade_\
        );

    \I__4353\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22323\
        );

    \I__4352\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22320\
        );

    \I__4351\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22317\
        );

    \I__4350\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22314\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__22323\,
            I => data_in_field_120
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__22320\,
            I => data_in_field_120
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__22317\,
            I => data_in_field_120
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__22314\,
            I => data_in_field_120
        );

    \I__4345\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22301\
        );

    \I__4344\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22298\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__22301\,
            I => \N__22295\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22291\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__22295\,
            I => \N__22288\
        );

    \I__4340\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22285\
        );

    \I__4339\ : Span4Mux_v
    port map (
            O => \N__22291\,
            I => \N__22279\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__22288\,
            I => \N__22279\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__22285\,
            I => \N__22276\
        );

    \I__4336\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22273\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__22279\,
            I => \N__22270\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__22276\,
            I => rand_data_30
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__22273\,
            I => rand_data_30
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__22270\,
            I => rand_data_30
        );

    \I__4331\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22256\
        );

    \I__4330\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22256\
        );

    \I__4329\ : InMux
    port map (
            O => \N__22261\,
            I => \N__22253\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__22256\,
            I => \N__22250\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__22253\,
            I => \c0.n8785\
        );

    \I__4326\ : Odrv12
    port map (
            O => \N__22250\,
            I => \c0.n8785\
        );

    \I__4325\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__4323\ : Span4Mux_h
    port map (
            O => \N__22239\,
            I => \N__22235\
        );

    \I__4322\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22232\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__22235\,
            I => \c0.n8887\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__22232\,
            I => \c0.n8887\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__22227\,
            I => \c0.n4240_cascade_\
        );

    \I__4318\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22220\
        );

    \I__4317\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22217\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__22220\,
            I => \N__22214\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__22217\,
            I => \N__22209\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__22214\,
            I => \N__22209\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__22209\,
            I => \N__22204\
        );

    \I__4312\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22201\
        );

    \I__4311\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22196\
        );

    \I__4310\ : Sp12to4
    port map (
            O => \N__22204\,
            I => \N__22191\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__22201\,
            I => \N__22191\
        );

    \I__4308\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22186\
        );

    \I__4307\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22186\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__22196\,
            I => \c0.data_in_field_13\
        );

    \I__4305\ : Odrv12
    port map (
            O => \N__22191\,
            I => \c0.data_in_field_13\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__22186\,
            I => \c0.data_in_field_13\
        );

    \I__4303\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22176\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__22176\,
            I => \N__22173\
        );

    \I__4301\ : Span4Mux_s2_h
    port map (
            O => \N__22173\,
            I => \N__22170\
        );

    \I__4300\ : Span4Mux_h
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__22167\,
            I => \c0.n44_adj_1609\
        );

    \I__4298\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22161\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__22161\,
            I => \c0.n4553\
        );

    \I__4296\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22152\
        );

    \I__4295\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22152\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22148\
        );

    \I__4293\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22143\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__22148\,
            I => \N__22140\
        );

    \I__4291\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22135\
        );

    \I__4290\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22135\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__22143\,
            I => data_in_field_53
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__22140\,
            I => data_in_field_53
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__22135\,
            I => data_in_field_53
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__4285\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__4283\ : Odrv12
    port map (
            O => \N__22119\,
            I => \c0.n8964\
        );

    \I__4282\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22113\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__4280\ : IoSpan4Mux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__4279\ : IoSpan4Mux
    port map (
            O => \N__22107\,
            I => \N__22104\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__22104\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__22101\,
            I => \N__22098\
        );

    \I__4276\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22094\
        );

    \I__4275\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22091\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__22094\,
            I => \N__22088\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__22091\,
            I => \N__22085\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__22088\,
            I => \N__22082\
        );

    \I__4271\ : Span4Mux_v
    port map (
            O => \N__22085\,
            I => \N__22079\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__22082\,
            I => \N__22076\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__22079\,
            I => \N__22073\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__22076\,
            I => \c0.n8942\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__22073\,
            I => \c0.n8942\
        );

    \I__4266\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__22065\,
            I => \N__22062\
        );

    \I__4264\ : Span4Mux_s2_h
    port map (
            O => \N__22062\,
            I => \N__22059\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__22059\,
            I => \N__22053\
        );

    \I__4262\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22050\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__22057\,
            I => \N__22047\
        );

    \I__4260\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22044\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__22053\,
            I => \N__22039\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__22050\,
            I => \N__22039\
        );

    \I__4257\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22036\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__22044\,
            I => \N__22031\
        );

    \I__4255\ : Span4Mux_s3_v
    port map (
            O => \N__22039\,
            I => \N__22031\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22028\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__22031\,
            I => data_in_field_57
        );

    \I__4252\ : Odrv12
    port map (
            O => \N__22028\,
            I => data_in_field_57
        );

    \I__4251\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22019\
        );

    \I__4250\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22013\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22010\
        );

    \I__4248\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22007\
        );

    \I__4247\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22004\
        );

    \I__4246\ : InMux
    port map (
            O => \N__22016\,
            I => \N__22001\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__21997\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__22010\,
            I => \N__21994\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__22007\,
            I => \N__21991\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__22004\,
            I => \N__21986\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21986\
        );

    \I__4240\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21983\
        );

    \I__4239\ : Span4Mux_s2_v
    port map (
            O => \N__21997\,
            I => \N__21980\
        );

    \I__4238\ : Span4Mux_h
    port map (
            O => \N__21994\,
            I => \N__21973\
        );

    \I__4237\ : Span4Mux_s3_h
    port map (
            O => \N__21991\,
            I => \N__21973\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__21986\,
            I => \N__21973\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__21983\,
            I => data_in_field_93
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__21980\,
            I => data_in_field_93
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__21973\,
            I => data_in_field_93
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__21966\,
            I => \N__21963\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__21954\,
            I => \c0.n4390\
        );

    \I__4227\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21946\
        );

    \I__4226\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21943\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__21949\,
            I => \N__21939\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__21946\,
            I => \N__21936\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__21943\,
            I => \N__21933\
        );

    \I__4222\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21930\
        );

    \I__4221\ : InMux
    port map (
            O => \N__21939\,
            I => \N__21925\
        );

    \I__4220\ : Span4Mux_s3_v
    port map (
            O => \N__21936\,
            I => \N__21922\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__21933\,
            I => \N__21917\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21917\
        );

    \I__4217\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21914\
        );

    \I__4216\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21911\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__21925\,
            I => \N__21908\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__21922\,
            I => \N__21903\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__21917\,
            I => \N__21903\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__21914\,
            I => data_in_field_87
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__21911\,
            I => data_in_field_87
        );

    \I__4210\ : Odrv12
    port map (
            O => \N__21908\,
            I => data_in_field_87
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__21903\,
            I => data_in_field_87
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__21894\,
            I => \N__21888\
        );

    \I__4207\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21885\
        );

    \I__4206\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21882\
        );

    \I__4205\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21877\
        );

    \I__4204\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21874\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__21885\,
            I => \N__21870\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21867\
        );

    \I__4201\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21864\
        );

    \I__4200\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21861\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__21877\,
            I => \N__21858\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__21874\,
            I => \N__21855\
        );

    \I__4197\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21852\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__21870\,
            I => \N__21849\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__21867\,
            I => \N__21844\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__21864\,
            I => \N__21844\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21837\
        );

    \I__4192\ : Span4Mux_s2_v
    port map (
            O => \N__21858\,
            I => \N__21837\
        );

    \I__4191\ : Span4Mux_h
    port map (
            O => \N__21855\,
            I => \N__21837\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__21852\,
            I => data_in_field_91
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__21849\,
            I => data_in_field_91
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__21844\,
            I => data_in_field_91
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__21837\,
            I => data_in_field_91
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__21828\,
            I => \N__21825\
        );

    \I__4185\ : InMux
    port map (
            O => \N__21825\,
            I => \N__21822\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__21822\,
            I => \N__21818\
        );

    \I__4183\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21815\
        );

    \I__4182\ : Span4Mux_h
    port map (
            O => \N__21818\,
            I => \N__21812\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__21815\,
            I => \c0.n8909\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__21812\,
            I => \c0.n8909\
        );

    \I__4179\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21801\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__21801\,
            I => \N__21798\
        );

    \I__4176\ : Odrv4
    port map (
            O => \N__21798\,
            I => \c0.n4197\
        );

    \I__4175\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21788\
        );

    \I__4174\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21788\
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__21793\,
            I => \N__21784\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21781\
        );

    \I__4171\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21778\
        );

    \I__4170\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21775\
        );

    \I__4169\ : Span4Mux_v
    port map (
            O => \N__21781\,
            I => \N__21771\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__21778\,
            I => \N__21766\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21766\
        );

    \I__4166\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21763\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__21771\,
            I => \N__21758\
        );

    \I__4164\ : Span4Mux_v
    port map (
            O => \N__21766\,
            I => \N__21758\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__21763\,
            I => data_in_field_60
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__21758\,
            I => data_in_field_60
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__21753\,
            I => \c0.n4197_cascade_\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__21750\,
            I => \N__21747\
        );

    \I__4159\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21744\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__21744\,
            I => \N__21741\
        );

    \I__4157\ : Span4Mux_h
    port map (
            O => \N__21741\,
            I => \N__21738\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__21738\,
            I => \c0.n4399\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__4154\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21727\
        );

    \I__4153\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21722\
        );

    \I__4152\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21722\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21719\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__21722\,
            I => \N__21714\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__21719\,
            I => \N__21711\
        );

    \I__4148\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21708\
        );

    \I__4147\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21705\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__21714\,
            I => \N__21698\
        );

    \I__4145\ : Span4Mux_v
    port map (
            O => \N__21711\,
            I => \N__21698\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__21708\,
            I => \N__21698\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__21705\,
            I => data_in_field_61
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__21698\,
            I => data_in_field_61
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__21693\,
            I => \c0.n4399_cascade_\
        );

    \I__4140\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21687\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21683\
        );

    \I__4138\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21680\
        );

    \I__4137\ : Odrv12
    port map (
            O => \N__21683\,
            I => \c0.n4288\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__21680\,
            I => \c0.n4288\
        );

    \I__4135\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21672\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__21672\,
            I => \c0.n10\
        );

    \I__4133\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21666\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__21666\,
            I => \N__21663\
        );

    \I__4131\ : Span4Mux_v
    port map (
            O => \N__21663\,
            I => \N__21658\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__21662\,
            I => \N__21655\
        );

    \I__4129\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21651\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__21658\,
            I => \N__21647\
        );

    \I__4127\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21642\
        );

    \I__4126\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21642\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__21651\,
            I => \N__21639\
        );

    \I__4124\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21636\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__21647\,
            I => rand_data_9
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__21642\,
            I => rand_data_9
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__21639\,
            I => rand_data_9
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__21636\,
            I => rand_data_9
        );

    \I__4119\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21619\
        );

    \I__4117\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21616\
        );

    \I__4116\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21613\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__21619\,
            I => \N__21608\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__21616\,
            I => \N__21603\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__21613\,
            I => \N__21603\
        );

    \I__4112\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21598\
        );

    \I__4111\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21598\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__21608\,
            I => data_in_field_121
        );

    \I__4109\ : Odrv12
    port map (
            O => \N__21603\,
            I => data_in_field_121
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__21598\,
            I => data_in_field_121
        );

    \I__4107\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21585\
        );

    \I__4106\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21585\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__21585\,
            I => \N__21581\
        );

    \I__4104\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21578\
        );

    \I__4103\ : Span12Mux_s4_v
    port map (
            O => \N__21581\,
            I => \N__21573\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__21578\,
            I => \N__21570\
        );

    \I__4101\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21567\
        );

    \I__4100\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21564\
        );

    \I__4099\ : Odrv12
    port map (
            O => \N__21573\,
            I => rand_data_15
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__21570\,
            I => rand_data_15
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__21567\,
            I => rand_data_15
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__21564\,
            I => rand_data_15
        );

    \I__4095\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21551\
        );

    \I__4094\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21546\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21543\
        );

    \I__4092\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21538\
        );

    \I__4091\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21538\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__21546\,
            I => \N__21532\
        );

    \I__4089\ : Span4Mux_s1_v
    port map (
            O => \N__21543\,
            I => \N__21532\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__21538\,
            I => \N__21529\
        );

    \I__4087\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21525\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__21532\,
            I => \N__21522\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__21529\,
            I => \N__21519\
        );

    \I__4084\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21516\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__21525\,
            I => data_in_field_143
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__21522\,
            I => data_in_field_143
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__21519\,
            I => data_in_field_143
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__21516\,
            I => data_in_field_143
        );

    \I__4079\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21502\
        );

    \I__4078\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21499\
        );

    \I__4077\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21496\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21493\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__21499\,
            I => \N__21490\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21487\
        );

    \I__4073\ : Span4Mux_h
    port map (
            O => \N__21493\,
            I => \N__21483\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__21490\,
            I => \N__21478\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__21487\,
            I => \N__21478\
        );

    \I__4070\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21475\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__21483\,
            I => \N__21472\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__21478\,
            I => rand_data_28
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__21475\,
            I => rand_data_28
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__21472\,
            I => rand_data_28
        );

    \I__4065\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21460\
        );

    \I__4064\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21455\
        );

    \I__4063\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21452\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__21460\,
            I => \N__21449\
        );

    \I__4061\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21446\
        );

    \I__4060\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21443\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__21455\,
            I => rand_data_13
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__21452\,
            I => rand_data_13
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__21449\,
            I => rand_data_13
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__21446\,
            I => rand_data_13
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__21443\,
            I => rand_data_13
        );

    \I__4054\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21426\
        );

    \I__4053\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21423\
        );

    \I__4052\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21420\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__21429\,
            I => \N__21417\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21414\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21411\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21406\
        );

    \I__4047\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21403\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__21414\,
            I => \N__21400\
        );

    \I__4045\ : Span4Mux_v
    port map (
            O => \N__21411\,
            I => \N__21397\
        );

    \I__4044\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21394\
        );

    \I__4043\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21391\
        );

    \I__4042\ : Span4Mux_h
    port map (
            O => \N__21406\,
            I => \N__21388\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__21403\,
            I => \c0.data_in_field_29\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__21400\,
            I => \c0.data_in_field_29\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__21397\,
            I => \c0.data_in_field_29\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__21394\,
            I => \c0.data_in_field_29\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__21391\,
            I => \c0.data_in_field_29\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__21388\,
            I => \c0.data_in_field_29\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__21375\,
            I => \N__21371\
        );

    \I__4034\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__4033\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21364\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__21368\,
            I => \N__21361\
        );

    \I__4031\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21358\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21354\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__21361\,
            I => \N__21351\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__21358\,
            I => \N__21348\
        );

    \I__4027\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21345\
        );

    \I__4026\ : Span4Mux_s3_h
    port map (
            O => \N__21354\,
            I => \N__21342\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__21351\,
            I => \N__21337\
        );

    \I__4024\ : Span4Mux_s3_h
    port map (
            O => \N__21348\,
            I => \N__21337\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__21345\,
            I => \c0.data_in_field_21\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__21342\,
            I => \c0.data_in_field_21\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__21337\,
            I => \c0.data_in_field_21\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__21330\,
            I => \c0.n9608_cascade_\
        );

    \I__4019\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21323\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__21326\,
            I => \N__21319\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21316\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__21322\,
            I => \N__21312\
        );

    \I__4015\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21309\
        );

    \I__4014\ : Span4Mux_v
    port map (
            O => \N__21316\,
            I => \N__21306\
        );

    \I__4013\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21303\
        );

    \I__4012\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21300\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__21309\,
            I => \c0.data_in_field_5\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__21306\,
            I => \c0.data_in_field_5\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__21303\,
            I => \c0.data_in_field_5\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__21300\,
            I => \c0.data_in_field_5\
        );

    \I__4007\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21288\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__21288\,
            I => \N__21285\
        );

    \I__4005\ : Span4Mux_s2_v
    port map (
            O => \N__21285\,
            I => \N__21282\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__21282\,
            I => \c0.n9147\
        );

    \I__4003\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21275\
        );

    \I__4002\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21271\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__21275\,
            I => \N__21268\
        );

    \I__4000\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21265\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21262\
        );

    \I__3998\ : Span4Mux_h
    port map (
            O => \N__21268\,
            I => \N__21259\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__21265\,
            I => \N__21255\
        );

    \I__3996\ : Span12Mux_v
    port map (
            O => \N__21262\,
            I => \N__21252\
        );

    \I__3995\ : Span4Mux_h
    port map (
            O => \N__21259\,
            I => \N__21249\
        );

    \I__3994\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21246\
        );

    \I__3993\ : Span12Mux_v
    port map (
            O => \N__21255\,
            I => \N__21243\
        );

    \I__3992\ : Odrv12
    port map (
            O => \N__21252\,
            I => rand_data_29
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__21249\,
            I => rand_data_29
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__21246\,
            I => rand_data_29
        );

    \I__3989\ : Odrv12
    port map (
            O => \N__21243\,
            I => rand_data_29
        );

    \I__3988\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21229\
        );

    \I__3987\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21226\
        );

    \I__3986\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21222\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21219\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21215\
        );

    \I__3983\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21212\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21209\
        );

    \I__3981\ : Span4Mux_h
    port map (
            O => \N__21219\,
            I => \N__21206\
        );

    \I__3980\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21203\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__21215\,
            I => \N__21200\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__21212\,
            I => \N__21197\
        );

    \I__3977\ : Span4Mux_s2_v
    port map (
            O => \N__21209\,
            I => \N__21192\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__21206\,
            I => \N__21192\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__21203\,
            I => data_in_field_109
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__21200\,
            I => data_in_field_109
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__21197\,
            I => data_in_field_109
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__21192\,
            I => data_in_field_109
        );

    \I__3971\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21176\
        );

    \I__3970\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21173\
        );

    \I__3969\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21168\
        );

    \I__3968\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21168\
        );

    \I__3967\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21165\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__21176\,
            I => rand_data_4
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__21173\,
            I => rand_data_4
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__21168\,
            I => rand_data_4
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__21165\,
            I => rand_data_4
        );

    \I__3962\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21150\
        );

    \I__3961\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21145\
        );

    \I__3960\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21145\
        );

    \I__3959\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21141\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__21150\,
            I => \N__21136\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__21145\,
            I => \N__21136\
        );

    \I__3956\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21133\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__21141\,
            I => rand_data_3
        );

    \I__3954\ : Odrv12
    port map (
            O => \N__21136\,
            I => rand_data_3
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__21133\,
            I => rand_data_3
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__21126\,
            I => \N__21122\
        );

    \I__3951\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21119\
        );

    \I__3950\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21116\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21113\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21108\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__21113\,
            I => \N__21108\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__21108\,
            I => \c0.n8992\
        );

    \I__3945\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__3943\ : Span4Mux_s2_h
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__3942\ : Span4Mux_h
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__21093\,
            I => \c0.n21_adj_1624\
        );

    \I__3940\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21086\
        );

    \I__3939\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21082\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__21086\,
            I => \N__21079\
        );

    \I__3937\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21076\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__21082\,
            I => \N__21072\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__21079\,
            I => \N__21067\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__21076\,
            I => \N__21067\
        );

    \I__3933\ : InMux
    port map (
            O => \N__21075\,
            I => \N__21064\
        );

    \I__3932\ : Span12Mux_v
    port map (
            O => \N__21072\,
            I => \N__21060\
        );

    \I__3931\ : Span4Mux_s3_h
    port map (
            O => \N__21067\,
            I => \N__21055\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21055\
        );

    \I__3929\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21052\
        );

    \I__3928\ : Odrv12
    port map (
            O => \N__21060\,
            I => rand_data_7
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__21055\,
            I => rand_data_7
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__21052\,
            I => rand_data_7
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__21045\,
            I => \N__21041\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__21044\,
            I => \N__21037\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21034\
        );

    \I__3922\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21031\
        );

    \I__3921\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21028\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__21023\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__21031\,
            I => \N__21023\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__21028\,
            I => \N__21020\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__21023\,
            I => \N__21015\
        );

    \I__3916\ : Span4Mux_v
    port map (
            O => \N__21020\,
            I => \N__21012\
        );

    \I__3915\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21009\
        );

    \I__3914\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21006\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__21015\,
            I => rand_data_1
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__21012\,
            I => rand_data_1
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__21009\,
            I => rand_data_1
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__21006\,
            I => rand_data_1
        );

    \I__3909\ : InMux
    port map (
            O => \N__20997\,
            I => \c0.n8116\
        );

    \I__3908\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20990\
        );

    \I__3907\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20987\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__20990\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__20987\,
            I => \c0.byte_transmit_counter2_5\
        );

    \I__3904\ : InMux
    port map (
            O => \N__20982\,
            I => \c0.n8117\
        );

    \I__3903\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20975\
        );

    \I__3902\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20972\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__20975\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__20972\,
            I => \c0.byte_transmit_counter2_6\
        );

    \I__3899\ : InMux
    port map (
            O => \N__20967\,
            I => \c0.n8118\
        );

    \I__3898\ : InMux
    port map (
            O => \N__20964\,
            I => \c0.n8119\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__20961\,
            I => \N__20957\
        );

    \I__3896\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20954\
        );

    \I__3895\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20951\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__20954\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__20951\,
            I => \c0.byte_transmit_counter2_7\
        );

    \I__3892\ : CEMux
    port map (
            O => \N__20946\,
            I => \N__20943\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__20937\,
            I => \c0.n4897\
        );

    \I__3888\ : SRMux
    port map (
            O => \N__20934\,
            I => \N__20931\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__20931\,
            I => \N__20928\
        );

    \I__3886\ : Span4Mux_h
    port map (
            O => \N__20928\,
            I => \N__20925\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__20925\,
            I => \c0.n5154\
        );

    \I__3884\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20917\
        );

    \I__3883\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20913\
        );

    \I__3882\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20910\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20907\
        );

    \I__3880\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20904\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__20913\,
            I => \N__20900\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__20910\,
            I => \N__20897\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__20907\,
            I => \N__20892\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20892\
        );

    \I__3875\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20889\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__20900\,
            I => rand_data_8
        );

    \I__3873\ : Odrv12
    port map (
            O => \N__20897\,
            I => rand_data_8
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__20892\,
            I => rand_data_8
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__20889\,
            I => rand_data_8
        );

    \I__3870\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20876\
        );

    \I__3869\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20872\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__20876\,
            I => \N__20869\
        );

    \I__3867\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20866\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__20872\,
            I => \N__20863\
        );

    \I__3865\ : Span4Mux_v
    port map (
            O => \N__20869\,
            I => \N__20858\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20858\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__20863\,
            I => \N__20855\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__20858\,
            I => \N__20852\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__20855\,
            I => \N__20849\
        );

    \I__3860\ : Span4Mux_h
    port map (
            O => \N__20852\,
            I => \N__20845\
        );

    \I__3859\ : Span4Mux_v
    port map (
            O => \N__20849\,
            I => \N__20842\
        );

    \I__3858\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20839\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__20845\,
            I => rand_data_22
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__20842\,
            I => rand_data_22
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__20839\,
            I => rand_data_22
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__20832\,
            I => \c0.n7194_cascade_\
        );

    \I__3853\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20826\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__20826\,
            I => \N__20823\
        );

    \I__3851\ : Span4Mux_h
    port map (
            O => \N__20823\,
            I => \N__20819\
        );

    \I__3850\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20816\
        );

    \I__3849\ : Span4Mux_s3_h
    port map (
            O => \N__20819\,
            I => \N__20811\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__20816\,
            I => \N__20811\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__20811\,
            I => \c0.n8449\
        );

    \I__3846\ : CEMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__20802\,
            I => \N__20799\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__20796\,
            I => n4839
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__20793\,
            I => \n4839_cascade_\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20786\
        );

    \I__3839\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20783\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20780\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__20783\,
            I => \N__20777\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__20780\,
            I => \N__20771\
        );

    \I__3835\ : Span4Mux_h
    port map (
            O => \N__20777\,
            I => \N__20768\
        );

    \I__3834\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20765\
        );

    \I__3833\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20760\
        );

    \I__3832\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20760\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__20771\,
            I => n31
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__20768\,
            I => n31
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__20765\,
            I => n31
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__20760\,
            I => n31
        );

    \I__3827\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20746\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__20750\,
            I => \N__20743\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__20749\,
            I => \N__20740\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20736\
        );

    \I__3823\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20733\
        );

    \I__3822\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20730\
        );

    \I__3821\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20727\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__20736\,
            I => \N__20724\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__20733\,
            I => \N__20719\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20719\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20711\
        );

    \I__3816\ : Span4Mux_h
    port map (
            O => \N__20724\,
            I => \N__20711\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__20719\,
            I => \N__20711\
        );

    \I__3814\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20708\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__20711\,
            I => \N__20705\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__20708\,
            I => data_in_field_65
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__20705\,
            I => data_in_field_65
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__20700\,
            I => \N__20697\
        );

    \I__3809\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20693\
        );

    \I__3808\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20690\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__20693\,
            I => \c0.tx2_transmit_N_1444\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__20690\,
            I => \c0.tx2_transmit_N_1444\
        );

    \I__3805\ : InMux
    port map (
            O => \N__20685\,
            I => \c0.n8113\
        );

    \I__3804\ : InMux
    port map (
            O => \N__20682\,
            I => \c0.n8114\
        );

    \I__3803\ : InMux
    port map (
            O => \N__20679\,
            I => \c0.n8115\
        );

    \I__3802\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20672\
        );

    \I__3801\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20668\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20665\
        );

    \I__3799\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20661\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20658\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__20665\,
            I => \N__20655\
        );

    \I__3796\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20652\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__20661\,
            I => rand_data_24
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__20658\,
            I => rand_data_24
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__20655\,
            I => rand_data_24
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__20652\,
            I => rand_data_24
        );

    \I__3791\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20640\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__20634\,
            I => n1903
        );

    \I__3787\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20626\
        );

    \I__3786\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20623\
        );

    \I__3785\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20620\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__20626\,
            I => \N__20617\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__20623\,
            I => \N__20614\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__20620\,
            I => \N__20609\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__20617\,
            I => \N__20609\
        );

    \I__3780\ : Span4Mux_s3_h
    port map (
            O => \N__20614\,
            I => \N__20606\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__20609\,
            I => \N__20601\
        );

    \I__3778\ : Span4Mux_h
    port map (
            O => \N__20606\,
            I => \N__20598\
        );

    \I__3777\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20593\
        );

    \I__3776\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20593\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20590\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__20598\,
            I => data_in_field_129
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__20593\,
            I => data_in_field_129
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__20590\,
            I => data_in_field_129
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__20583\,
            I => \N__20580\
        );

    \I__3770\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20574\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__20574\,
            I => \N__20571\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__20571\,
            I => \N__20568\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__20568\,
            I => \N__20565\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__20565\,
            I => \c0.n8791\
        );

    \I__3764\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20558\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__20561\,
            I => \N__20555\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__20558\,
            I => \N__20552\
        );

    \I__3761\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20549\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__20552\,
            I => \N__20546\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20542\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__20546\,
            I => \N__20539\
        );

    \I__3757\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20536\
        );

    \I__3756\ : Span4Mux_v
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__20539\,
            I => data_in_6_0
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__20536\,
            I => data_in_6_0
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__20533\,
            I => data_in_6_0
        );

    \I__3752\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__20520\,
            I => \N__20515\
        );

    \I__3749\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20510\
        );

    \I__3748\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20510\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__20515\,
            I => data_in_5_0
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__20510\,
            I => data_in_5_0
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__20505\,
            I => \c0.n19_adj_1665_cascade_\
        );

    \I__3744\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20496\
        );

    \I__3743\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20496\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20492\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__20495\,
            I => \N__20489\
        );

    \I__3740\ : Span4Mux_h
    port map (
            O => \N__20492\,
            I => \N__20486\
        );

    \I__3739\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20483\
        );

    \I__3738\ : Span4Mux_v
    port map (
            O => \N__20486\,
            I => \N__20480\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__20483\,
            I => tx2_active
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__20480\,
            I => tx2_active
        );

    \I__3735\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20468\
        );

    \I__3734\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20468\
        );

    \I__3733\ : InMux
    port map (
            O => \N__20473\,
            I => \N__20465\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20460\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20460\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__20460\,
            I => \N__20457\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__20457\,
            I => \N__20453\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__20456\,
            I => \N__20450\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__20453\,
            I => \N__20446\
        );

    \I__3726\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20441\
        );

    \I__3725\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20441\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__20446\,
            I => \c0.r_SM_Main_2_N_1483_0\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__20441\,
            I => \c0.r_SM_Main_2_N_1483_0\
        );

    \I__3722\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__20433\,
            I => \c0.n19_adj_1665\
        );

    \I__3720\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20426\
        );

    \I__3719\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20423\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__20426\,
            I => rx_data_6
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__20423\,
            I => rx_data_6
        );

    \I__3716\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20415\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__20415\,
            I => \N__20411\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20408\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__20411\,
            I => \N__20405\
        );

    \I__3712\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20402\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__20405\,
            I => rx_data_4
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__20402\,
            I => rx_data_4
        );

    \I__3709\ : InMux
    port map (
            O => \N__20397\,
            I => \N__20391\
        );

    \I__3708\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20391\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__20391\,
            I => rx_data_7
        );

    \I__3706\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20382\
        );

    \I__3705\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20382\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__20382\,
            I => data_in_20_7
        );

    \I__3703\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20375\
        );

    \I__3702\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20372\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__20375\,
            I => data_in_19_7
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__20372\,
            I => data_in_19_7
        );

    \I__3699\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20362\
        );

    \I__3698\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20357\
        );

    \I__3697\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20357\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__20362\,
            I => n4044
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__20357\,
            I => n4044
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__20352\,
            I => \N__20348\
        );

    \I__3693\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20345\
        );

    \I__3692\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20342\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__20345\,
            I => rx_data_5
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__20342\,
            I => rx_data_5
        );

    \I__3689\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20331\
        );

    \I__3688\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20328\
        );

    \I__3687\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20323\
        );

    \I__3686\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20323\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__20331\,
            I => \N__20320\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20317\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__20323\,
            I => n4049
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__20320\,
            I => n4049
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__20317\,
            I => n4049
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__3679\ : InMux
    port map (
            O => \N__20307\,
            I => \N__20304\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__3677\ : Span4Mux_s2_h
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__3676\ : Span4Mux_h
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__20292\,
            I => \c0.n9476\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__20289\,
            I => \N__20286\
        );

    \I__3672\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20283\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__20283\,
            I => \N__20279\
        );

    \I__3670\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20276\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__20279\,
            I => n4
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__20276\,
            I => n4
        );

    \I__3667\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20267\
        );

    \I__3666\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20264\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__20267\,
            I => rx_data_3
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__20264\,
            I => rx_data_3
        );

    \I__3663\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20255\
        );

    \I__3662\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20252\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__20255\,
            I => data_in_19_6
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__20252\,
            I => data_in_19_6
        );

    \I__3659\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20243\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__20246\,
            I => \N__20240\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20237\
        );

    \I__3656\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20234\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__20237\,
            I => \N__20231\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__20234\,
            I => rx_data_0
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__20231\,
            I => rx_data_0
        );

    \I__3652\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20223\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20220\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__20220\,
            I => \N__20216\
        );

    \I__3649\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20213\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__20216\,
            I => data_in_18_7
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__20213\,
            I => data_in_18_7
        );

    \I__3646\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20202\
        );

    \I__3645\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20202\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__20202\,
            I => data_in_20_6
        );

    \I__3643\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__20196\,
            I => n4_adj_1725
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__20193\,
            I => \n4_adj_1725_cascade_\
        );

    \I__3640\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20186\
        );

    \I__3639\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20183\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__20186\,
            I => rx_data_1
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__20183\,
            I => rx_data_1
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__20178\,
            I => \n4044_cascade_\
        );

    \I__3635\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20169\
        );

    \I__3634\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20169\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__20169\,
            I => data_in_16_5
        );

    \I__3632\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20162\
        );

    \I__3631\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20159\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__20162\,
            I => data_in_18_5
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__20159\,
            I => data_in_18_5
        );

    \I__3628\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20148\
        );

    \I__3627\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20148\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__20148\,
            I => data_in_17_5
        );

    \I__3625\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20141\
        );

    \I__3624\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20138\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__20141\,
            I => data_in_18_6
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__20138\,
            I => data_in_18_6
        );

    \I__3621\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20130\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__20130\,
            I => \N__20127\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__20127\,
            I => \N__20123\
        );

    \I__3618\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20120\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__20123\,
            I => data_in_18_1
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__20120\,
            I => data_in_18_1
        );

    \I__3615\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20109\
        );

    \I__3614\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20109\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__20109\,
            I => data_in_19_1
        );

    \I__3612\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20100\
        );

    \I__3611\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20100\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__20100\,
            I => data_in_20_1
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__20097\,
            I => \N__20094\
        );

    \I__3608\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20088\
        );

    \I__3607\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20088\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__20088\,
            I => rx_data_2
        );

    \I__3605\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20082\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__20082\,
            I => \N__20078\
        );

    \I__3603\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20075\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__20078\,
            I => data_in_12_3
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__20075\,
            I => data_in_12_3
        );

    \I__3600\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20067\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__20067\,
            I => \N__20063\
        );

    \I__3598\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20060\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__20063\,
            I => data_in_11_3
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__20060\,
            I => data_in_11_3
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__20055\,
            I => \c0.n9590_cascade_\
        );

    \I__3594\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__20049\,
            I => \c0.n9153\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__20046\,
            I => \c0.n9156_cascade_\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__20043\,
            I => \c0.n9584_cascade_\
        );

    \I__3590\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__3588\ : Span12Mux_s3_v
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__3587\ : Odrv12
    port map (
            O => \N__20031\,
            I => \c0.n9150\
        );

    \I__3586\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20025\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__20016\,
            I => \c0.n22_adj_1678\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__20013\,
            I => \c0.n9587_cascade_\
        );

    \I__3580\ : InMux
    port map (
            O => \N__20010\,
            I => \N__20007\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__20004\,
            I => \c0.tx2.r_Tx_Data_5\
        );

    \I__3577\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19998\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19995\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__19995\,
            I => \N__19991\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19988\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__19991\,
            I => data_in_10_5
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__19988\,
            I => data_in_10_5
        );

    \I__3571\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19977\
        );

    \I__3570\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19977\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__19977\,
            I => data_in_11_5
        );

    \I__3568\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19970\
        );

    \I__3567\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19967\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__19970\,
            I => data_in_13_5
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__19967\,
            I => data_in_13_5
        );

    \I__3564\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19956\
        );

    \I__3563\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19956\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__19956\,
            I => data_in_12_5
        );

    \I__3561\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19949\
        );

    \I__3560\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19946\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__19949\,
            I => data_in_14_5
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__19946\,
            I => data_in_14_5
        );

    \I__3557\ : InMux
    port map (
            O => \N__19941\,
            I => \N__19935\
        );

    \I__3556\ : InMux
    port map (
            O => \N__19940\,
            I => \N__19935\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__19935\,
            I => data_in_15_5
        );

    \I__3554\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19924\
        );

    \I__3552\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19921\
        );

    \I__3551\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19917\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__19924\,
            I => \N__19914\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__19921\,
            I => \N__19911\
        );

    \I__3548\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19907\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__19917\,
            I => \N__19902\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__19914\,
            I => \N__19902\
        );

    \I__3545\ : Span4Mux_s2_v
    port map (
            O => \N__19911\,
            I => \N__19899\
        );

    \I__3544\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19896\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__19907\,
            I => data_in_field_141
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__19902\,
            I => data_in_field_141
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__19899\,
            I => data_in_field_141
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__19896\,
            I => data_in_field_141
        );

    \I__3539\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19883\
        );

    \I__3538\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19879\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__19883\,
            I => \N__19876\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19872\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19867\
        );

    \I__3534\ : Span12Mux_v
    port map (
            O => \N__19876\,
            I => \N__19867\
        );

    \I__3533\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19864\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__19872\,
            I => rand_data_21
        );

    \I__3531\ : Odrv12
    port map (
            O => \N__19867\,
            I => rand_data_21
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__19864\,
            I => rand_data_21
        );

    \I__3529\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19853\
        );

    \I__3528\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19849\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__19853\,
            I => \N__19846\
        );

    \I__3526\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19843\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__19849\,
            I => \N__19840\
        );

    \I__3524\ : Span4Mux_h
    port map (
            O => \N__19846\,
            I => \N__19836\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19833\
        );

    \I__3522\ : Span12Mux_v
    port map (
            O => \N__19840\,
            I => \N__19830\
        );

    \I__3521\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19827\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__19836\,
            I => rand_data_17
        );

    \I__3519\ : Odrv12
    port map (
            O => \N__19833\,
            I => rand_data_17
        );

    \I__3518\ : Odrv12
    port map (
            O => \N__19830\,
            I => rand_data_17
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__19827\,
            I => rand_data_17
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__19818\,
            I => \N__19814\
        );

    \I__3515\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19811\
        );

    \I__3514\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19808\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__19811\,
            I => \N__19805\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19802\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__19805\,
            I => \N__19795\
        );

    \I__3510\ : Span4Mux_s2_h
    port map (
            O => \N__19802\,
            I => \N__19795\
        );

    \I__3509\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19790\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19790\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__19795\,
            I => \N__19787\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__19790\,
            I => data_in_field_113
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__19787\,
            I => data_in_field_113
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__19782\,
            I => \N__19778\
        );

    \I__3503\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19775\
        );

    \I__3502\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19772\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__19775\,
            I => \N__19766\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19763\
        );

    \I__3499\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19760\
        );

    \I__3498\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19757\
        );

    \I__3497\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19754\
        );

    \I__3496\ : Sp12to4
    port map (
            O => \N__19766\,
            I => \N__19747\
        );

    \I__3495\ : Sp12to4
    port map (
            O => \N__19763\,
            I => \N__19747\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19747\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19744\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__19754\,
            I => data_in_field_149
        );

    \I__3491\ : Odrv12
    port map (
            O => \N__19747\,
            I => data_in_field_149
        );

    \I__3490\ : Odrv12
    port map (
            O => \N__19744\,
            I => data_in_field_149
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__3488\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19731\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__3486\ : Span4Mux_v
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__19725\,
            I => \c0.n1893_adj_1635\
        );

    \I__3484\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__19716\,
            I => \N__19711\
        );

    \I__3481\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19708\
        );

    \I__3480\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19705\
        );

    \I__3479\ : Sp12to4
    port map (
            O => \N__19711\,
            I => \N__19699\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__19708\,
            I => \N__19699\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__19705\,
            I => \N__19696\
        );

    \I__3476\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19693\
        );

    \I__3475\ : Odrv12
    port map (
            O => \N__19699\,
            I => rand_data_23
        );

    \I__3474\ : Odrv12
    port map (
            O => \N__19696\,
            I => rand_data_23
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__19693\,
            I => rand_data_23
        );

    \I__3472\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19681\
        );

    \I__3471\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19678\
        );

    \I__3470\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19673\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19670\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19667\
        );

    \I__3467\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19664\
        );

    \I__3466\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19661\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19658\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__19670\,
            I => \N__19655\
        );

    \I__3463\ : Span4Mux_s1_v
    port map (
            O => \N__19667\,
            I => \N__19650\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19650\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19645\
        );

    \I__3460\ : Span4Mux_v
    port map (
            O => \N__19658\,
            I => \N__19645\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__19655\,
            I => data_in_field_85
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__19650\,
            I => data_in_field_85
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__19645\,
            I => data_in_field_85
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__19638\,
            I => \c0.n9596_cascade_\
        );

    \I__3455\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19628\
        );

    \I__3453\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19624\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__19628\,
            I => \N__19621\
        );

    \I__3451\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19618\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__19624\,
            I => data_in_field_117
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__19621\,
            I => data_in_field_117
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__19618\,
            I => data_in_field_117
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__19611\,
            I => \N__19607\
        );

    \I__3446\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19602\
        );

    \I__3445\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19602\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__19602\,
            I => \N__19598\
        );

    \I__3443\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19595\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__19598\,
            I => \N__19592\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__19595\,
            I => \N__19589\
        );

    \I__3440\ : Span4Mux_s2_v
    port map (
            O => \N__19592\,
            I => \N__19585\
        );

    \I__3439\ : Span12Mux_v
    port map (
            O => \N__19589\,
            I => \N__19582\
        );

    \I__3438\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19579\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__19585\,
            I => rand_data_25
        );

    \I__3436\ : Odrv12
    port map (
            O => \N__19582\,
            I => rand_data_25
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__19579\,
            I => rand_data_25
        );

    \I__3434\ : InMux
    port map (
            O => \N__19572\,
            I => n8179
        );

    \I__3433\ : InMux
    port map (
            O => \N__19569\,
            I => n8180
        );

    \I__3432\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19562\
        );

    \I__3431\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19559\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__19562\,
            I => \N__19556\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__19559\,
            I => \N__19553\
        );

    \I__3428\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19549\
        );

    \I__3427\ : Span4Mux_v
    port map (
            O => \N__19553\,
            I => \N__19546\
        );

    \I__3426\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19543\
        );

    \I__3425\ : Sp12to4
    port map (
            O => \N__19549\,
            I => \N__19540\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__19546\,
            I => \N__19534\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__19543\,
            I => \N__19534\
        );

    \I__3422\ : Span12Mux_s5_h
    port map (
            O => \N__19540\,
            I => \N__19531\
        );

    \I__3421\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19528\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__19534\,
            I => rand_data_27
        );

    \I__3419\ : Odrv12
    port map (
            O => \N__19531\,
            I => rand_data_27
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__19528\,
            I => rand_data_27
        );

    \I__3417\ : InMux
    port map (
            O => \N__19521\,
            I => n8181
        );

    \I__3416\ : InMux
    port map (
            O => \N__19518\,
            I => n8182
        );

    \I__3415\ : InMux
    port map (
            O => \N__19515\,
            I => n8183
        );

    \I__3414\ : InMux
    port map (
            O => \N__19512\,
            I => n8184
        );

    \I__3413\ : InMux
    port map (
            O => \N__19509\,
            I => n8185
        );

    \I__3412\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19503\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__19503\,
            I => \N__19497\
        );

    \I__3410\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19494\
        );

    \I__3409\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19489\
        );

    \I__3408\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19489\
        );

    \I__3407\ : Span4Mux_v
    port map (
            O => \N__19497\,
            I => \N__19486\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__19494\,
            I => rand_data_31
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__19489\,
            I => rand_data_31
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__19486\,
            I => rand_data_31
        );

    \I__3403\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19470\
        );

    \I__3401\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19467\
        );

    \I__3400\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19462\
        );

    \I__3399\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19462\
        );

    \I__3398\ : Span4Mux_s2_v
    port map (
            O => \N__19470\,
            I => \N__19459\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__19467\,
            I => data_in_field_104
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__19462\,
            I => data_in_field_104
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__19459\,
            I => data_in_field_104
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__19452\,
            I => \c0.n9734_cascade_\
        );

    \I__3393\ : InMux
    port map (
            O => \N__19449\,
            I => \bfn_6_29_0_\
        );

    \I__3392\ : InMux
    port map (
            O => \N__19446\,
            I => n8171
        );

    \I__3391\ : InMux
    port map (
            O => \N__19443\,
            I => n8172
        );

    \I__3390\ : InMux
    port map (
            O => \N__19440\,
            I => \N__19435\
        );

    \I__3389\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19432\
        );

    \I__3388\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19429\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__19435\,
            I => \N__19424\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__19432\,
            I => \N__19424\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__19429\,
            I => \N__19421\
        );

    \I__3384\ : Span4Mux_h
    port map (
            O => \N__19424\,
            I => \N__19417\
        );

    \I__3383\ : Span12Mux_s5_h
    port map (
            O => \N__19421\,
            I => \N__19414\
        );

    \I__3382\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19411\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__19417\,
            I => rand_data_19
        );

    \I__3380\ : Odrv12
    port map (
            O => \N__19414\,
            I => rand_data_19
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__19411\,
            I => rand_data_19
        );

    \I__3378\ : InMux
    port map (
            O => \N__19404\,
            I => n8173
        );

    \I__3377\ : InMux
    port map (
            O => \N__19401\,
            I => n8174
        );

    \I__3376\ : InMux
    port map (
            O => \N__19398\,
            I => n8175
        );

    \I__3375\ : InMux
    port map (
            O => \N__19395\,
            I => n8176
        );

    \I__3374\ : InMux
    port map (
            O => \N__19392\,
            I => n8177
        );

    \I__3373\ : InMux
    port map (
            O => \N__19389\,
            I => \bfn_6_30_0_\
        );

    \I__3372\ : InMux
    port map (
            O => \N__19386\,
            I => n8161
        );

    \I__3371\ : InMux
    port map (
            O => \N__19383\,
            I => \bfn_6_28_0_\
        );

    \I__3370\ : InMux
    port map (
            O => \N__19380\,
            I => n8163
        );

    \I__3369\ : InMux
    port map (
            O => \N__19377\,
            I => n8164
        );

    \I__3368\ : InMux
    port map (
            O => \N__19374\,
            I => n8165
        );

    \I__3367\ : InMux
    port map (
            O => \N__19371\,
            I => n8166
        );

    \I__3366\ : InMux
    port map (
            O => \N__19368\,
            I => n8167
        );

    \I__3365\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19362\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__19362\,
            I => \N__19358\
        );

    \I__3363\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19355\
        );

    \I__3362\ : Sp12to4
    port map (
            O => \N__19358\,
            I => \N__19347\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__19355\,
            I => \N__19347\
        );

    \I__3360\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19344\
        );

    \I__3359\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19341\
        );

    \I__3358\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19338\
        );

    \I__3357\ : Odrv12
    port map (
            O => \N__19347\,
            I => rand_data_14
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__19344\,
            I => rand_data_14
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__19341\,
            I => rand_data_14
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__19338\,
            I => rand_data_14
        );

    \I__3353\ : InMux
    port map (
            O => \N__19329\,
            I => n8168
        );

    \I__3352\ : InMux
    port map (
            O => \N__19326\,
            I => n8169
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__19323\,
            I => \c0.n4897_cascade_\
        );

    \I__3350\ : InMux
    port map (
            O => \N__19320\,
            I => \bfn_6_27_0_\
        );

    \I__3349\ : InMux
    port map (
            O => \N__19317\,
            I => n8155
        );

    \I__3348\ : InMux
    port map (
            O => \N__19314\,
            I => n8156
        );

    \I__3347\ : InMux
    port map (
            O => \N__19311\,
            I => n8157
        );

    \I__3346\ : InMux
    port map (
            O => \N__19308\,
            I => n8158
        );

    \I__3345\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19300\
        );

    \I__3344\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19296\
        );

    \I__3343\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19293\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__19300\,
            I => \N__19290\
        );

    \I__3341\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19287\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__19296\,
            I => \N__19284\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__19293\,
            I => \N__19281\
        );

    \I__3338\ : Span4Mux_v
    port map (
            O => \N__19290\,
            I => \N__19278\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__19287\,
            I => \N__19273\
        );

    \I__3336\ : Sp12to4
    port map (
            O => \N__19284\,
            I => \N__19273\
        );

    \I__3335\ : Span12Mux_s4_h
    port map (
            O => \N__19281\,
            I => \N__19265\
        );

    \I__3334\ : Sp12to4
    port map (
            O => \N__19278\,
            I => \N__19265\
        );

    \I__3333\ : Span12Mux_s5_v
    port map (
            O => \N__19273\,
            I => \N__19265\
        );

    \I__3332\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19262\
        );

    \I__3331\ : Odrv12
    port map (
            O => \N__19265\,
            I => rand_data_5
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__19262\,
            I => rand_data_5
        );

    \I__3329\ : InMux
    port map (
            O => \N__19257\,
            I => n8159
        );

    \I__3328\ : InMux
    port map (
            O => \N__19254\,
            I => n8160
        );

    \I__3327\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__19248\,
            I => n9091
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__19245\,
            I => \n9092_cascade_\
        );

    \I__3324\ : IoInMux
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__3322\ : Span4Mux_s2_v
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__3321\ : Span4Mux_v
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__19230\,
            I => \LED_c\
        );

    \I__3319\ : SRMux
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__3317\ : Span12Mux_v
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__3316\ : Odrv12
    port map (
            O => \N__19218\,
            I => n8761
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \N__19210\
        );

    \I__3314\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19207\
        );

    \I__3313\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19203\
        );

    \I__3312\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19200\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19197\
        );

    \I__3310\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19194\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__19203\,
            I => data_in_field_48
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__19200\,
            I => data_in_field_48
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__19197\,
            I => data_in_field_48
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__19194\,
            I => data_in_field_48
        );

    \I__3305\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__19182\,
            I => \N__19176\
        );

    \I__3303\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19173\
        );

    \I__3302\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19168\
        );

    \I__3301\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19168\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__19176\,
            I => \N__19165\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__19173\,
            I => data_in_1_4
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__19168\,
            I => data_in_1_4
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__19165\,
            I => data_in_1_4
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__3295\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19143\
        );

    \I__3294\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19138\
        );

    \I__3293\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19138\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__19152\,
            I => \N__19135\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__19151\,
            I => \N__19121\
        );

    \I__3290\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19114\
        );

    \I__3289\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19109\
        );

    \I__3288\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19105\
        );

    \I__3287\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19102\
        );

    \I__3286\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19099\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__19143\,
            I => \N__19096\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__19138\,
            I => \N__19093\
        );

    \I__3283\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19090\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__19134\,
            I => \N__19081\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19078\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__19132\,
            I => \N__19075\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__19131\,
            I => \N__19071\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__19130\,
            I => \N__19068\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__19129\,
            I => \N__19050\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__19128\,
            I => \N__19047\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__19127\,
            I => \N__19042\
        );

    \I__3274\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19036\
        );

    \I__3273\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19027\
        );

    \I__3272\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19027\
        );

    \I__3271\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19027\
        );

    \I__3270\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19027\
        );

    \I__3269\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19020\
        );

    \I__3268\ : InMux
    port map (
            O => \N__19118\,
            I => \N__19020\
        );

    \I__3267\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19020\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19017\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19012\
        );

    \I__3264\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19012\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19009\
        );

    \I__3262\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19006\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19003\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__19102\,
            I => \N__18992\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__18992\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__19096\,
            I => \N__18992\
        );

    \I__3257\ : Span4Mux_s1_h
    port map (
            O => \N__19093\,
            I => \N__18992\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__19090\,
            I => \N__18992\
        );

    \I__3255\ : InMux
    port map (
            O => \N__19089\,
            I => \N__18987\
        );

    \I__3254\ : InMux
    port map (
            O => \N__19088\,
            I => \N__18987\
        );

    \I__3253\ : InMux
    port map (
            O => \N__19087\,
            I => \N__18982\
        );

    \I__3252\ : InMux
    port map (
            O => \N__19086\,
            I => \N__18982\
        );

    \I__3251\ : InMux
    port map (
            O => \N__19085\,
            I => \N__18971\
        );

    \I__3250\ : InMux
    port map (
            O => \N__19084\,
            I => \N__18971\
        );

    \I__3249\ : InMux
    port map (
            O => \N__19081\,
            I => \N__18971\
        );

    \I__3248\ : InMux
    port map (
            O => \N__19078\,
            I => \N__18971\
        );

    \I__3247\ : InMux
    port map (
            O => \N__19075\,
            I => \N__18971\
        );

    \I__3246\ : InMux
    port map (
            O => \N__19074\,
            I => \N__18964\
        );

    \I__3245\ : InMux
    port map (
            O => \N__19071\,
            I => \N__18964\
        );

    \I__3244\ : InMux
    port map (
            O => \N__19068\,
            I => \N__18964\
        );

    \I__3243\ : InMux
    port map (
            O => \N__19067\,
            I => \N__18959\
        );

    \I__3242\ : InMux
    port map (
            O => \N__19066\,
            I => \N__18959\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19065\,
            I => \N__18956\
        );

    \I__3240\ : InMux
    port map (
            O => \N__19064\,
            I => \N__18949\
        );

    \I__3239\ : InMux
    port map (
            O => \N__19063\,
            I => \N__18949\
        );

    \I__3238\ : InMux
    port map (
            O => \N__19062\,
            I => \N__18949\
        );

    \I__3237\ : InMux
    port map (
            O => \N__19061\,
            I => \N__18934\
        );

    \I__3236\ : InMux
    port map (
            O => \N__19060\,
            I => \N__18934\
        );

    \I__3235\ : InMux
    port map (
            O => \N__19059\,
            I => \N__18934\
        );

    \I__3234\ : InMux
    port map (
            O => \N__19058\,
            I => \N__18934\
        );

    \I__3233\ : InMux
    port map (
            O => \N__19057\,
            I => \N__18934\
        );

    \I__3232\ : InMux
    port map (
            O => \N__19056\,
            I => \N__18934\
        );

    \I__3231\ : InMux
    port map (
            O => \N__19055\,
            I => \N__18934\
        );

    \I__3230\ : InMux
    port map (
            O => \N__19054\,
            I => \N__18923\
        );

    \I__3229\ : InMux
    port map (
            O => \N__19053\,
            I => \N__18923\
        );

    \I__3228\ : InMux
    port map (
            O => \N__19050\,
            I => \N__18923\
        );

    \I__3227\ : InMux
    port map (
            O => \N__19047\,
            I => \N__18923\
        );

    \I__3226\ : InMux
    port map (
            O => \N__19046\,
            I => \N__18923\
        );

    \I__3225\ : InMux
    port map (
            O => \N__19045\,
            I => \N__18912\
        );

    \I__3224\ : InMux
    port map (
            O => \N__19042\,
            I => \N__18912\
        );

    \I__3223\ : InMux
    port map (
            O => \N__19041\,
            I => \N__18912\
        );

    \I__3222\ : InMux
    port map (
            O => \N__19040\,
            I => \N__18912\
        );

    \I__3221\ : InMux
    port map (
            O => \N__19039\,
            I => \N__18912\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__19036\,
            I => \N__18907\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__19027\,
            I => \N__18907\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__19020\,
            I => \N__18904\
        );

    \I__3217\ : Span12Mux_s3_h
    port map (
            O => \N__19017\,
            I => \N__18901\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__19012\,
            I => \N__18896\
        );

    \I__3215\ : Span4Mux_v
    port map (
            O => \N__19009\,
            I => \N__18896\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__19006\,
            I => \N__18889\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__19003\,
            I => \N__18889\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__18992\,
            I => \N__18889\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__18987\,
            I => n9069
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__18982\,
            I => n9069
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__18971\,
            I => n9069
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__18964\,
            I => n9069
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__18959\,
            I => n9069
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__18956\,
            I => n9069
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__18949\,
            I => n9069
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__18934\,
            I => n9069
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__18923\,
            I => n9069
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__18912\,
            I => n9069
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__18907\,
            I => n9069
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__18904\,
            I => n9069
        );

    \I__3199\ : Odrv12
    port map (
            O => \N__18901\,
            I => n9069
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__18896\,
            I => n9069
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__18889\,
            I => n9069
        );

    \I__3196\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18854\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__18857\,
            I => \N__18851\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18846\
        );

    \I__3193\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18843\
        );

    \I__3192\ : InMux
    port map (
            O => \N__18850\,
            I => \N__18840\
        );

    \I__3191\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18837\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__18846\,
            I => \N__18834\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__18843\,
            I => \N__18831\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__18840\,
            I => data_in_field_45
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__18837\,
            I => data_in_field_45
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__18834\,
            I => data_in_field_45
        );

    \I__3185\ : Odrv12
    port map (
            O => \N__18831\,
            I => data_in_field_45
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__3183\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18816\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__18816\,
            I => \c0.n9602\
        );

    \I__3181\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18809\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \N__18806\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18803\
        );

    \I__3178\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18798\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__18803\,
            I => \N__18795\
        );

    \I__3176\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18792\
        );

    \I__3175\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18789\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__18798\,
            I => \c0.data_in_field_12\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__18795\,
            I => \c0.data_in_field_12\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__18792\,
            I => \c0.data_in_field_12\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__18789\,
            I => \c0.data_in_field_12\
        );

    \I__3170\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18777\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18774\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__18774\,
            I => \N__18770\
        );

    \I__3167\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18767\
        );

    \I__3166\ : Sp12to4
    port map (
            O => \N__18770\,
            I => \N__18762\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__18767\,
            I => \N__18762\
        );

    \I__3164\ : Odrv12
    port map (
            O => \N__18762\,
            I => \c0.n9019\
        );

    \I__3163\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18754\
        );

    \I__3162\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18751\
        );

    \I__3161\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18748\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__18754\,
            I => \N__18745\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__18751\,
            I => \N__18740\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__18748\,
            I => \N__18737\
        );

    \I__3157\ : Span4Mux_h
    port map (
            O => \N__18745\,
            I => \N__18734\
        );

    \I__3156\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18729\
        );

    \I__3155\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18729\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__18740\,
            I => \c0.data_in_field_28\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__18737\,
            I => \c0.data_in_field_28\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__18734\,
            I => \c0.data_in_field_28\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__18729\,
            I => \c0.data_in_field_28\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__18720\,
            I => \c0.n9746_cascade_\
        );

    \I__3149\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18712\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18708\
        );

    \I__3147\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18704\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__18712\,
            I => \N__18701\
        );

    \I__3145\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18698\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__18708\,
            I => \N__18695\
        );

    \I__3143\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18692\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__18704\,
            I => \c0.data_in_field_32\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__18701\,
            I => \c0.data_in_field_32\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__18698\,
            I => \c0.data_in_field_32\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__18695\,
            I => \c0.data_in_field_32\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__18692\,
            I => \c0.data_in_field_32\
        );

    \I__3137\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__18678\,
            I => \N__18672\
        );

    \I__3135\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18669\
        );

    \I__3134\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18665\
        );

    \I__3133\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18662\
        );

    \I__3132\ : Span4Mux_h
    port map (
            O => \N__18672\,
            I => \N__18659\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__18669\,
            I => \N__18656\
        );

    \I__3130\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18653\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__18665\,
            I => data_in_field_42
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__18662\,
            I => data_in_field_42
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__18659\,
            I => data_in_field_42
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__18656\,
            I => data_in_field_42
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__18653\,
            I => data_in_field_42
        );

    \I__3124\ : InMux
    port map (
            O => \N__18642\,
            I => \N__18637\
        );

    \I__3123\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18631\
        );

    \I__3122\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18628\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18625\
        );

    \I__3120\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18622\
        );

    \I__3119\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18617\
        );

    \I__3118\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18617\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__18631\,
            I => data_in_field_40
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__18628\,
            I => data_in_field_40
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__18625\,
            I => data_in_field_40
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__18622\,
            I => data_in_field_40
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__18617\,
            I => data_in_field_40
        );

    \I__3112\ : InMux
    port map (
            O => \N__18606\,
            I => \N__18603\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__18603\,
            I => \N__18598\
        );

    \I__3110\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18593\
        );

    \I__3109\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18593\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__18598\,
            I => \N__18590\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18587\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__18590\,
            I => \c0.n4208\
        );

    \I__3105\ : Odrv12
    port map (
            O => \N__18587\,
            I => \c0.n4208\
        );

    \I__3104\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18579\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__18579\,
            I => \N__18574\
        );

    \I__3102\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18570\
        );

    \I__3101\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18567\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__18574\,
            I => \N__18564\
        );

    \I__3099\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18561\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__18570\,
            I => data_in_3_4
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__18567\,
            I => data_in_3_4
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__18564\,
            I => data_in_3_4
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__18561\,
            I => data_in_3_4
        );

    \I__3094\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18548\
        );

    \I__3093\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18545\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__18548\,
            I => \N__18540\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18537\
        );

    \I__3090\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18534\
        );

    \I__3089\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18531\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__18540\,
            I => \N__18528\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__18537\,
            I => data_in_3_2
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__18534\,
            I => data_in_3_2
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__18531\,
            I => data_in_3_2
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__18528\,
            I => data_in_3_2
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__18519\,
            I => \N__18516\
        );

    \I__3082\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18512\
        );

    \I__3081\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18509\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__18512\,
            I => \N__18504\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18501\
        );

    \I__3078\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18496\
        );

    \I__3077\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18496\
        );

    \I__3076\ : Span4Mux_h
    port map (
            O => \N__18504\,
            I => \N__18493\
        );

    \I__3075\ : Span4Mux_h
    port map (
            O => \N__18501\,
            I => \N__18490\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__18496\,
            I => data_in_2_4
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__18493\,
            I => data_in_2_4
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__18490\,
            I => data_in_2_4
        );

    \I__3071\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18479\
        );

    \I__3070\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18476\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__18479\,
            I => data_in_17_0
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__18476\,
            I => data_in_17_0
        );

    \I__3067\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18467\
        );

    \I__3066\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18464\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__18467\,
            I => \N__18459\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18459\
        );

    \I__3063\ : Span4Mux_h
    port map (
            O => \N__18459\,
            I => \N__18456\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__18456\,
            I => \N__18453\
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__18453\,
            I => \c0.n8960\
        );

    \I__3060\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18446\
        );

    \I__3059\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18443\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18440\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__18443\,
            I => \N__18436\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__18440\,
            I => \N__18433\
        );

    \I__3055\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18430\
        );

    \I__3054\ : Span4Mux_h
    port map (
            O => \N__18436\,
            I => \N__18427\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__18433\,
            I => data_in_0_4
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__18430\,
            I => data_in_0_4
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__18427\,
            I => data_in_0_4
        );

    \I__3050\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18417\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__18417\,
            I => \N__18414\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__18414\,
            I => n1890
        );

    \I__3047\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18408\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__18408\,
            I => \N__18405\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__18405\,
            I => \N__18401\
        );

    \I__3044\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18398\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__18401\,
            I => data_in_14_0
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__18398\,
            I => data_in_14_0
        );

    \I__3041\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18387\
        );

    \I__3040\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18387\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__18387\,
            I => data_in_15_0
        );

    \I__3038\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18376\
        );

    \I__3036\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18370\
        );

    \I__3035\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18370\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__18376\,
            I => \N__18367\
        );

    \I__3033\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18364\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18361\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__18367\,
            I => data_in_2_2
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__18364\,
            I => data_in_2_2
        );

    \I__3029\ : Odrv12
    port map (
            O => \N__18361\,
            I => data_in_2_2
        );

    \I__3028\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18348\
        );

    \I__3027\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18348\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__18348\,
            I => data_in_16_0
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__3024\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18336\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18336\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__18336\,
            I => data_in_20_0
        );

    \I__3021\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__18330\,
            I => \N__18327\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__18327\,
            I => n1898
        );

    \I__3018\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18320\
        );

    \I__3017\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18317\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__18320\,
            I => data_in_20_5
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__18317\,
            I => data_in_20_5
        );

    \I__3014\ : InMux
    port map (
            O => \N__18312\,
            I => \N__18303\
        );

    \I__3013\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18303\
        );

    \I__3012\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18303\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__18303\,
            I => data_in_5_5
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__18300\,
            I => \N__18297\
        );

    \I__3009\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__18294\,
            I => \N__18291\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__18291\,
            I => \N__18286\
        );

    \I__3006\ : InMux
    port map (
            O => \N__18290\,
            I => \N__18283\
        );

    \I__3005\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18280\
        );

    \I__3004\ : Span4Mux_h
    port map (
            O => \N__18286\,
            I => \N__18277\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__18283\,
            I => data_in_4_5
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__18280\,
            I => data_in_4_5
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__18277\,
            I => data_in_4_5
        );

    \I__3000\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18261\
        );

    \I__2999\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18261\
        );

    \I__2998\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18261\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__18261\,
            I => data_in_6_5
        );

    \I__2996\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18252\
        );

    \I__2995\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18252\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__18252\,
            I => data_in_7_5
        );

    \I__2993\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18243\
        );

    \I__2992\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18243\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__18243\,
            I => data_in_8_5
        );

    \I__2990\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18234\
        );

    \I__2989\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18234\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__18234\,
            I => data_in_9_5
        );

    \I__2987\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18227\
        );

    \I__2986\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18224\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__18227\,
            I => data_in_16_3
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__18224\,
            I => data_in_16_3
        );

    \I__2983\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18213\
        );

    \I__2982\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18213\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__18213\,
            I => data_in_15_3
        );

    \I__2980\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18206\
        );

    \I__2979\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18203\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__18206\,
            I => data_in_17_3
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__18203\,
            I => data_in_17_3
        );

    \I__2976\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18194\
        );

    \I__2975\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18191\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__18194\,
            I => data_in_18_3
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__18191\,
            I => data_in_18_3
        );

    \I__2972\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18180\
        );

    \I__2971\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18180\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__18180\,
            I => data_in_19_3
        );

    \I__2969\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18171\
        );

    \I__2968\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18171\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__18171\,
            I => data_in_20_3
        );

    \I__2966\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18162\
        );

    \I__2965\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18162\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__18162\,
            I => data_in_19_5
        );

    \I__2963\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18156\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__18156\,
            I => \N__18152\
        );

    \I__2961\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18149\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__18152\,
            I => data_in_17_6
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__18149\,
            I => data_in_17_6
        );

    \I__2958\ : InMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__18141\,
            I => \N__18137\
        );

    \I__2956\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18134\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__18137\,
            I => data_in_10_3
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__18134\,
            I => data_in_10_3
        );

    \I__2953\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__18126\,
            I => \N__18122\
        );

    \I__2951\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18119\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__18122\,
            I => data_in_9_3
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__18119\,
            I => data_in_9_3
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \c0.n3056_cascade_\
        );

    \I__2947\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__2945\ : Span4Mux_h
    port map (
            O => \N__18105\,
            I => \N__18102\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__18102\,
            I => \c0.n22_adj_1676\
        );

    \I__2943\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18096\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__18096\,
            I => \c0.n38_adj_1616\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__2940\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18087\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__18084\,
            I => \c0.n36\
        );

    \I__2937\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18078\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__18078\,
            I => \c0.n37\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__2934\ : InMux
    port map (
            O => \N__18072\,
            I => \N__18069\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__18069\,
            I => \c0.data_in_frame_19_7\
        );

    \I__2932\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18063\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__18063\,
            I => \N__18058\
        );

    \I__2930\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18052\
        );

    \I__2929\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18052\
        );

    \I__2928\ : Span4Mux_s2_v
    port map (
            O => \N__18058\,
            I => \N__18049\
        );

    \I__2927\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18046\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__18052\,
            I => data_in_field_135
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__18049\,
            I => data_in_field_135
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__18046\,
            I => data_in_field_135
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__18039\,
            I => \c0.n9662_cascade_\
        );

    \I__2922\ : InMux
    port map (
            O => \N__18036\,
            I => \N__18033\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18033\,
            I => \c0.n9665\
        );

    \I__2920\ : InMux
    port map (
            O => \N__18030\,
            I => \N__18024\
        );

    \I__2919\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18024\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__18024\,
            I => data_in_13_3
        );

    \I__2917\ : InMux
    port map (
            O => \N__18021\,
            I => \N__18015\
        );

    \I__2916\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18015\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__18015\,
            I => data_in_14_3
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__18012\,
            I => \c0.n6_adj_1604_cascade_\
        );

    \I__2913\ : InMux
    port map (
            O => \N__18009\,
            I => \N__18006\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__18006\,
            I => \N__18003\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__18003\,
            I => \N__18000\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__18000\,
            I => \c0.n8983\
        );

    \I__2909\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17994\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17991\
        );

    \I__2907\ : Span12Mux_s5_v
    port map (
            O => \N__17991\,
            I => \N__17988\
        );

    \I__2906\ : Odrv12
    port map (
            O => \N__17988\,
            I => \c0.n8948\
        );

    \I__2905\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17982\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__17979\,
            I => \c0.n8945\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__17976\,
            I => \c0.n8983_cascade_\
        );

    \I__2901\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17970\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__2899\ : Span12Mux_s3_v
    port map (
            O => \N__17967\,
            I => \N__17963\
        );

    \I__2898\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17960\
        );

    \I__2897\ : Odrv12
    port map (
            O => \N__17963\,
            I => \c0.n9004\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__17960\,
            I => \c0.n9004\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \N__17951\
        );

    \I__2894\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17948\
        );

    \I__2893\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17945\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__17948\,
            I => \N__17939\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__17945\,
            I => \N__17936\
        );

    \I__2890\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17933\
        );

    \I__2889\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17928\
        );

    \I__2888\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17928\
        );

    \I__2887\ : Span12Mux_h
    port map (
            O => \N__17939\,
            I => \N__17925\
        );

    \I__2886\ : Span4Mux_s2_h
    port map (
            O => \N__17936\,
            I => \N__17922\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__17933\,
            I => data_in_field_89
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__17928\,
            I => data_in_field_89
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__17925\,
            I => data_in_field_89
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__17922\,
            I => data_in_field_89
        );

    \I__2881\ : InMux
    port map (
            O => \N__17913\,
            I => \N__17909\
        );

    \I__2880\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17906\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__17909\,
            I => \N__17903\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__17906\,
            I => \c0.n4203\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__17903\,
            I => \c0.n4203\
        );

    \I__2876\ : InMux
    port map (
            O => \N__17898\,
            I => \N__17895\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17895\,
            I => \N__17892\
        );

    \I__2874\ : Span4Mux_s2_v
    port map (
            O => \N__17892\,
            I => \N__17889\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__17889\,
            I => \c0.n8890\
        );

    \I__2872\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17882\
        );

    \I__2871\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17879\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__17882\,
            I => \c0.n8874\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__17879\,
            I => \c0.n8874\
        );

    \I__2868\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17871\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__2866\ : Span4Mux_s2_v
    port map (
            O => \N__17868\,
            I => \N__17865\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__17865\,
            I => \c0.n24_adj_1607\
        );

    \I__2864\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17859\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__17859\,
            I => \c0.n23\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__17856\,
            I => \c0.n25_cascade_\
        );

    \I__2861\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17850\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__17850\,
            I => \c0.n26_adj_1606\
        );

    \I__2859\ : InMux
    port map (
            O => \N__17847\,
            I => \N__17844\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__17844\,
            I => \N__17841\
        );

    \I__2857\ : Span4Mux_v
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__2856\ : Span4Mux_h
    port map (
            O => \N__17838\,
            I => \N__17835\
        );

    \I__2855\ : Odrv4
    port map (
            O => \N__17835\,
            I => \c0.data_in_frame_20_3\
        );

    \I__2854\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17829\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__17829\,
            I => \N__17825\
        );

    \I__2852\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17822\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__17825\,
            I => \N__17819\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17816\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__17819\,
            I => \N__17811\
        );

    \I__2848\ : Span4Mux_s1_v
    port map (
            O => \N__17816\,
            I => \N__17811\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__17811\,
            I => \N__17808\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__17808\,
            I => \c0.n8974\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__2844\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17799\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__2842\ : Span4Mux_s2_v
    port map (
            O => \N__17796\,
            I => \N__17793\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__17793\,
            I => \c0.n22_adj_1617\
        );

    \I__2840\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17787\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__17787\,
            I => \N__17784\
        );

    \I__2838\ : Span4Mux_s3_v
    port map (
            O => \N__17784\,
            I => \N__17781\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__17781\,
            I => \c0.n8933\
        );

    \I__2836\ : InMux
    port map (
            O => \N__17778\,
            I => \N__17775\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__17775\,
            I => \N__17772\
        );

    \I__2834\ : Span4Mux_s2_v
    port map (
            O => \N__17772\,
            I => \N__17769\
        );

    \I__2833\ : Span4Mux_v
    port map (
            O => \N__17769\,
            I => \N__17766\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__17766\,
            I => \c0.data_in_frame_20_7\
        );

    \I__2831\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17757\
        );

    \I__2830\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17757\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__17757\,
            I => \N__17752\
        );

    \I__2828\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17749\
        );

    \I__2827\ : InMux
    port map (
            O => \N__17755\,
            I => \N__17746\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__17752\,
            I => \N__17741\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17741\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__17746\,
            I => data_in_field_111
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__17741\,
            I => data_in_field_111
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__17736\,
            I => \c0.n4525_cascade_\
        );

    \I__2821\ : InMux
    port map (
            O => \N__17733\,
            I => \N__17729\
        );

    \I__2820\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17725\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__17729\,
            I => \N__17722\
        );

    \I__2818\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17719\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__17725\,
            I => \N__17714\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__17722\,
            I => \N__17714\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__17719\,
            I => data_in_field_107
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__17714\,
            I => data_in_field_107
        );

    \I__2813\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17706\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__17706\,
            I => \N__17700\
        );

    \I__2811\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17697\
        );

    \I__2810\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17692\
        );

    \I__2809\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17692\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__17700\,
            I => \N__17687\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__17697\,
            I => \N__17687\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__17692\,
            I => data_in_field_137
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__17687\,
            I => data_in_field_137
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__17682\,
            I => \c0.n8874_cascade_\
        );

    \I__2803\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17675\
        );

    \I__2802\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17672\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__17675\,
            I => \N__17668\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__17672\,
            I => \N__17665\
        );

    \I__2799\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17661\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__17668\,
            I => \N__17658\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__17665\,
            I => \N__17655\
        );

    \I__2796\ : InMux
    port map (
            O => \N__17664\,
            I => \N__17652\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__17661\,
            I => data_in_field_55
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__17658\,
            I => data_in_field_55
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__17655\,
            I => data_in_field_55
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__17652\,
            I => data_in_field_55
        );

    \I__2791\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17640\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__17640\,
            I => \c0.n6_adj_1636\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__17637\,
            I => \N__17633\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \N__17630\
        );

    \I__2787\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17627\
        );

    \I__2786\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17624\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__17627\,
            I => \N__17621\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17618\
        );

    \I__2783\ : Span4Mux_h
    port map (
            O => \N__17621\,
            I => \N__17615\
        );

    \I__2782\ : Span12Mux_v
    port map (
            O => \N__17618\,
            I => \N__17612\
        );

    \I__2781\ : Span4Mux_h
    port map (
            O => \N__17615\,
            I => \N__17609\
        );

    \I__2780\ : Odrv12
    port map (
            O => \N__17612\,
            I => \c0.n8989\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__17609\,
            I => \c0.n8989\
        );

    \I__2778\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17599\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__17603\,
            I => \N__17596\
        );

    \I__2776\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17590\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__17599\,
            I => \N__17586\
        );

    \I__2774\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17583\
        );

    \I__2773\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17580\
        );

    \I__2772\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17577\
        );

    \I__2771\ : InMux
    port map (
            O => \N__17593\,
            I => \N__17574\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__17590\,
            I => \N__17571\
        );

    \I__2769\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17568\
        );

    \I__2768\ : Span4Mux_s2_v
    port map (
            O => \N__17586\,
            I => \N__17563\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__17583\,
            I => \N__17563\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__17580\,
            I => data_in_field_63
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__17577\,
            I => data_in_field_63
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__17574\,
            I => data_in_field_63
        );

    \I__2763\ : Odrv12
    port map (
            O => \N__17571\,
            I => data_in_field_63
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__17568\,
            I => data_in_field_63
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__17563\,
            I => data_in_field_63
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__17550\,
            I => \N__17546\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__17549\,
            I => \N__17543\
        );

    \I__2758\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17537\
        );

    \I__2757\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17534\
        );

    \I__2756\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17527\
        );

    \I__2755\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17527\
        );

    \I__2754\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17527\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17524\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__17534\,
            I => \N__17521\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__17527\,
            I => \N__17514\
        );

    \I__2750\ : Span4Mux_h
    port map (
            O => \N__17524\,
            I => \N__17514\
        );

    \I__2749\ : Span4Mux_s3_h
    port map (
            O => \N__17521\,
            I => \N__17514\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__17514\,
            I => data_in_field_59
        );

    \I__2747\ : InMux
    port map (
            O => \N__17511\,
            I => \N__17507\
        );

    \I__2746\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17504\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__17507\,
            I => \N__17498\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__17504\,
            I => \N__17495\
        );

    \I__2743\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17490\
        );

    \I__2742\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17490\
        );

    \I__2741\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17487\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__17498\,
            I => \N__17484\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__17495\,
            I => \N__17479\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17479\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__17487\,
            I => data_in_field_51
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__17484\,
            I => data_in_field_51
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__17479\,
            I => data_in_field_51
        );

    \I__2734\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17469\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17465\
        );

    \I__2732\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17462\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__17465\,
            I => \N__17457\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17457\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__17454\,
            I => \c0.n4302\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__17451\,
            I => \N__17447\
        );

    \I__2726\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17443\
        );

    \I__2725\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17440\
        );

    \I__2724\ : InMux
    port map (
            O => \N__17446\,
            I => \N__17437\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__17443\,
            I => \N__17432\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__17440\,
            I => \N__17429\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17426\
        );

    \I__2720\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17423\
        );

    \I__2719\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17420\
        );

    \I__2718\ : Span4Mux_v
    port map (
            O => \N__17432\,
            I => \N__17413\
        );

    \I__2717\ : Span4Mux_s3_v
    port map (
            O => \N__17429\,
            I => \N__17413\
        );

    \I__2716\ : Span4Mux_s3_v
    port map (
            O => \N__17426\,
            I => \N__17413\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__17423\,
            I => data_in_field_79
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__17420\,
            I => data_in_field_79
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__17413\,
            I => data_in_field_79
        );

    \I__2712\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17403\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__17403\,
            I => \N__17399\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17395\
        );

    \I__2709\ : Span4Mux_v
    port map (
            O => \N__17399\,
            I => \N__17390\
        );

    \I__2708\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17387\
        );

    \I__2707\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17384\
        );

    \I__2706\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17381\
        );

    \I__2705\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17378\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__17390\,
            I => \N__17375\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17372\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__17384\,
            I => \N__17369\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__17381\,
            I => data_in_field_139
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__17378\,
            I => data_in_field_139
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__17375\,
            I => data_in_field_139
        );

    \I__2698\ : Odrv12
    port map (
            O => \N__17372\,
            I => data_in_field_139
        );

    \I__2697\ : Odrv12
    port map (
            O => \N__17369\,
            I => data_in_field_139
        );

    \I__2696\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17354\
        );

    \I__2695\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17351\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17348\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__17351\,
            I => \N__17343\
        );

    \I__2692\ : Span4Mux_h
    port map (
            O => \N__17348\,
            I => \N__17343\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__17343\,
            I => \c0.n8825\
        );

    \I__2690\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17337\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__17337\,
            I => \N__17334\
        );

    \I__2688\ : Odrv12
    port map (
            O => \N__17334\,
            I => \c0.n6_adj_1654\
        );

    \I__2687\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__17328\,
            I => \c0.n4253\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__17325\,
            I => \N__17322\
        );

    \I__2684\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17316\
        );

    \I__2682\ : Odrv12
    port map (
            O => \N__17316\,
            I => \c0.n4151\
        );

    \I__2681\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17306\
        );

    \I__2680\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17306\
        );

    \I__2679\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17301\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__17306\,
            I => \N__17298\
        );

    \I__2677\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17295\
        );

    \I__2676\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17292\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__17301\,
            I => \N__17289\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__17298\,
            I => \N__17286\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__17295\,
            I => \N__17283\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__17292\,
            I => \c0.data_in_field_17\
        );

    \I__2671\ : Odrv12
    port map (
            O => \N__17289\,
            I => \c0.data_in_field_17\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__17286\,
            I => \c0.data_in_field_17\
        );

    \I__2669\ : Odrv12
    port map (
            O => \N__17283\,
            I => \c0.data_in_field_17\
        );

    \I__2668\ : InMux
    port map (
            O => \N__17274\,
            I => \N__17271\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__17271\,
            I => \N__17268\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__17268\,
            I => \c0.n45\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__17265\,
            I => \N__17262\
        );

    \I__2664\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17258\
        );

    \I__2663\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17255\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__17258\,
            I => \N__17251\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17248\
        );

    \I__2660\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17245\
        );

    \I__2659\ : Span4Mux_v
    port map (
            O => \N__17251\,
            I => \N__17242\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__17248\,
            I => \c0.n4183\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__17245\,
            I => \c0.n4183\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__17242\,
            I => \c0.n4183\
        );

    \I__2655\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17232\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__17232\,
            I => \N__17229\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__17229\,
            I => \N__17225\
        );

    \I__2652\ : InMux
    port map (
            O => \N__17228\,
            I => \N__17222\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__17225\,
            I => \c0.n8864\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__17222\,
            I => \c0.n8864\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__17217\,
            I => \N__17214\
        );

    \I__2648\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17211\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__17211\,
            I => \N__17208\
        );

    \I__2646\ : Odrv12
    port map (
            O => \N__17208\,
            I => \c0.n8843\
        );

    \I__2645\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17201\
        );

    \I__2644\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17198\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__17201\,
            I => \N__17195\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__17198\,
            I => \c0.n8930\
        );

    \I__2641\ : Odrv12
    port map (
            O => \N__17195\,
            I => \c0.n8930\
        );

    \I__2640\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17187\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__17187\,
            I => \N__17184\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__17184\,
            I => \N__17181\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__17181\,
            I => \c0.n20\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__17178\,
            I => \c0.n21_cascade_\
        );

    \I__2635\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17172\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__17172\,
            I => \N__17169\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__17169\,
            I => \N__17166\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__17166\,
            I => \c0.n19\
        );

    \I__2631\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17160\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__17160\,
            I => \c0.n18\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__17157\,
            I => \c0.n8421_cascade_\
        );

    \I__2628\ : InMux
    port map (
            O => \N__17154\,
            I => \N__17150\
        );

    \I__2627\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17147\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__17150\,
            I => \N__17144\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__17147\,
            I => \N__17141\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__17144\,
            I => \c0.tx2_transmit_N_1334\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__17141\,
            I => \c0.tx2_transmit_N_1334\
        );

    \I__2622\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17133\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__17133\,
            I => \c0.n24_adj_1605\
        );

    \I__2620\ : InMux
    port map (
            O => \N__17130\,
            I => \N__17127\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__17127\,
            I => \N__17121\
        );

    \I__2618\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17118\
        );

    \I__2617\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17113\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17113\
        );

    \I__2615\ : Span12Mux_s5_v
    port map (
            O => \N__17121\,
            I => \N__17110\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__17118\,
            I => data_in_field_75
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__17113\,
            I => data_in_field_75
        );

    \I__2612\ : Odrv12
    port map (
            O => \N__17110\,
            I => data_in_field_75
        );

    \I__2611\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17100\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__17100\,
            I => \N__17094\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17089\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17089\
        );

    \I__2607\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17086\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__17094\,
            I => \N__17083\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__17089\,
            I => \N__17080\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__17086\,
            I => data_in_field_67
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__17083\,
            I => data_in_field_67
        );

    \I__2602\ : Odrv12
    port map (
            O => \N__17080\,
            I => data_in_field_67
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__17073\,
            I => \c0.n9506_cascade_\
        );

    \I__2600\ : InMux
    port map (
            O => \N__17070\,
            I => \N__17064\
        );

    \I__2599\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17061\
        );

    \I__2598\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17058\
        );

    \I__2597\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17054\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__17064\,
            I => \N__17051\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__17061\,
            I => \N__17046\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__17058\,
            I => \N__17046\
        );

    \I__2593\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17043\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__17054\,
            I => \c0.data_in_field_34\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__17051\,
            I => \c0.data_in_field_34\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__17046\,
            I => \c0.data_in_field_34\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__17043\,
            I => \c0.data_in_field_34\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__17034\,
            I => \c0.n4_adj_1592_cascade_\
        );

    \I__2587\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17028\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__17028\,
            I => \N__17025\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__17025\,
            I => \N__17022\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__17022\,
            I => \c0.n4324\
        );

    \I__2583\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17016\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__17016\,
            I => \c0.n21_adj_1599\
        );

    \I__2581\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17010\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__17010\,
            I => \N__17007\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__17007\,
            I => \N__17003\
        );

    \I__2578\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17000\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__17003\,
            I => \c0.n4200\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__17000\,
            I => \c0.n4200\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__16995\,
            I => \N__16992\
        );

    \I__2574\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16989\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__16989\,
            I => \c0.n28\
        );

    \I__2572\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16983\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__16983\,
            I => \c0.n23_adj_1608\
        );

    \I__2570\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16977\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__16977\,
            I => \N__16974\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__16974\,
            I => \N__16968\
        );

    \I__2567\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16963\
        );

    \I__2566\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16963\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16960\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__16968\,
            I => data_in_1_7
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__16963\,
            I => data_in_1_7
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__16960\,
            I => data_in_1_7
        );

    \I__2561\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16950\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__16950\,
            I => \N__16947\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__16947\,
            I => \N__16942\
        );

    \I__2558\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16937\
        );

    \I__2557\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16937\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__16942\,
            I => \c0.data_in_field_15\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__16937\,
            I => \c0.data_in_field_15\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__16932\,
            I => \n1895_cascade_\
        );

    \I__2553\ : InMux
    port map (
            O => \N__16929\,
            I => \N__16926\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__16926\,
            I => \N__16923\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__16923\,
            I => n1889
        );

    \I__2550\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16917\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16914\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__16914\,
            I => \N__16911\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__16911\,
            I => n1897
        );

    \I__2546\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16904\
        );

    \I__2545\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16901\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__16904\,
            I => \N__16897\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__16901\,
            I => \N__16894\
        );

    \I__2542\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16891\
        );

    \I__2541\ : Odrv12
    port map (
            O => \N__16897\,
            I => data_in_4_4
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__16894\,
            I => data_in_4_4
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__16891\,
            I => data_in_4_4
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__16884\,
            I => \N__16880\
        );

    \I__2537\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16875\
        );

    \I__2536\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16872\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__16879\,
            I => \N__16869\
        );

    \I__2534\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16866\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__16875\,
            I => \N__16863\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__16872\,
            I => \N__16860\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16857\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__16866\,
            I => data_in_2_0
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__16863\,
            I => data_in_2_0
        );

    \I__2528\ : Odrv12
    port map (
            O => \N__16860\,
            I => data_in_2_0
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__16857\,
            I => data_in_2_0
        );

    \I__2526\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16843\
        );

    \I__2525\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16840\
        );

    \I__2524\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16836\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__16843\,
            I => \N__16833\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__16840\,
            I => \N__16830\
        );

    \I__2521\ : InMux
    port map (
            O => \N__16839\,
            I => \N__16827\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__16836\,
            I => \c0.data_in_field_26\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__16833\,
            I => \c0.data_in_field_26\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__16830\,
            I => \c0.data_in_field_26\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__16827\,
            I => \c0.data_in_field_26\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__16818\,
            I => \N__16813\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__16817\,
            I => \N__16810\
        );

    \I__2514\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16807\
        );

    \I__2513\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16802\
        );

    \I__2512\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16799\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16807\,
            I => \N__16796\
        );

    \I__2510\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16793\
        );

    \I__2509\ : InMux
    port map (
            O => \N__16805\,
            I => \N__16790\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__16802\,
            I => \c0.data_in_field_18\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__16799\,
            I => \c0.data_in_field_18\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__16796\,
            I => \c0.data_in_field_18\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__16793\,
            I => \c0.data_in_field_18\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__16790\,
            I => \c0.data_in_field_18\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__16779\,
            I => \N__16776\
        );

    \I__2502\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16773\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__16773\,
            I => \N__16770\
        );

    \I__2500\ : Span12Mux_s4_h
    port map (
            O => \N__16770\,
            I => \N__16767\
        );

    \I__2499\ : Odrv12
    port map (
            O => \N__16767\,
            I => \c0.n9512\
        );

    \I__2498\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16761\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__16761\,
            I => \N__16757\
        );

    \I__2496\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16754\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__16757\,
            I => \N__16751\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__16754\,
            I => \N__16746\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__16751\,
            I => \N__16743\
        );

    \I__2492\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16738\
        );

    \I__2491\ : InMux
    port map (
            O => \N__16749\,
            I => \N__16738\
        );

    \I__2490\ : Span4Mux_h
    port map (
            O => \N__16746\,
            I => \N__16735\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__16743\,
            I => data_in_2_1
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__16738\,
            I => data_in_2_1
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__16735\,
            I => data_in_2_1
        );

    \I__2486\ : InMux
    port map (
            O => \N__16728\,
            I => \N__16725\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__16725\,
            I => \N__16722\
        );

    \I__2484\ : Span4Mux_h
    port map (
            O => \N__16722\,
            I => \N__16719\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__16719\,
            I => \c0.n4492\
        );

    \I__2482\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16713\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__16713\,
            I => \N__16709\
        );

    \I__2480\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16706\
        );

    \I__2479\ : Span4Mux_h
    port map (
            O => \N__16709\,
            I => \N__16703\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__16706\,
            I => \c0.n24\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__16703\,
            I => \c0.n24\
        );

    \I__2476\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16694\
        );

    \I__2475\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16691\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__16694\,
            I => \c0.n8902\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__16691\,
            I => \c0.n8902\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__16686\,
            I => \c0.n4492_cascade_\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__16683\,
            I => \c0.n8948_cascade_\
        );

    \I__2470\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16677\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__16677\,
            I => \N__16673\
        );

    \I__2468\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16670\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__16673\,
            I => \N__16667\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__16670\,
            I => \N__16664\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__16667\,
            I => \c0.n8858\
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__16664\,
            I => \c0.n8858\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__16659\,
            I => \N__16656\
        );

    \I__2462\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16653\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__16653\,
            I => \c0.n19_adj_1602\
        );

    \I__2460\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16647\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__16647\,
            I => \N__16643\
        );

    \I__2458\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16639\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__16643\,
            I => \N__16636\
        );

    \I__2456\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16633\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__16639\,
            I => data_in_0_1
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__16636\,
            I => data_in_0_1
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__16633\,
            I => data_in_0_1
        );

    \I__2452\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16623\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__16623\,
            I => \N__16620\
        );

    \I__2450\ : Span4Mux_h
    port map (
            O => \N__16620\,
            I => \N__16617\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__16617\,
            I => \N__16611\
        );

    \I__2448\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16608\
        );

    \I__2447\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16603\
        );

    \I__2446\ : InMux
    port map (
            O => \N__16614\,
            I => \N__16603\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__16611\,
            I => \c0.data_in_field_1\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__16608\,
            I => \c0.data_in_field_1\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__16603\,
            I => \c0.data_in_field_1\
        );

    \I__2442\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16587\
        );

    \I__2441\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16587\
        );

    \I__2440\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16587\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__16587\,
            I => data_in_6_6
        );

    \I__2438\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16581\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__16581\,
            I => \N__16577\
        );

    \I__2436\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16574\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__16577\,
            I => \N__16571\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__16574\,
            I => data_in_8_6
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__16571\,
            I => data_in_8_6
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__16566\,
            I => \N__16563\
        );

    \I__2431\ : InMux
    port map (
            O => \N__16563\,
            I => \N__16557\
        );

    \I__2430\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16557\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__16557\,
            I => data_in_7_6
        );

    \I__2428\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__16545\,
            I => \N__16539\
        );

    \I__2424\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16534\
        );

    \I__2423\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16534\
        );

    \I__2422\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16531\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__16539\,
            I => data_in_3_5
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__16534\,
            I => data_in_3_5
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__16531\,
            I => data_in_3_5
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__16524\,
            I => \N__16521\
        );

    \I__2417\ : InMux
    port map (
            O => \N__16521\,
            I => \N__16515\
        );

    \I__2416\ : InMux
    port map (
            O => \N__16520\,
            I => \N__16508\
        );

    \I__2415\ : InMux
    port map (
            O => \N__16519\,
            I => \N__16508\
        );

    \I__2414\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16508\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__16515\,
            I => data_in_3_6
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__16508\,
            I => data_in_3_6
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__16503\,
            I => \c0.n8843_cascade_\
        );

    \I__2410\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16497\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__16497\,
            I => \N__16493\
        );

    \I__2408\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16490\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__16493\,
            I => \N__16484\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__16490\,
            I => \N__16481\
        );

    \I__2405\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16478\
        );

    \I__2404\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16473\
        );

    \I__2403\ : InMux
    port map (
            O => \N__16487\,
            I => \N__16473\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__16484\,
            I => \c0.data_in_field_31\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__16481\,
            I => \c0.data_in_field_31\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__16478\,
            I => \c0.data_in_field_31\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__16473\,
            I => \c0.data_in_field_31\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__16464\,
            I => \c0.n4151_cascade_\
        );

    \I__2397\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16451\
        );

    \I__2396\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16451\
        );

    \I__2395\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16451\
        );

    \I__2394\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16448\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__16451\,
            I => \c0.data_in_field_30\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__16448\,
            I => \c0.data_in_field_30\
        );

    \I__2391\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16440\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__16440\,
            I => \N__16436\
        );

    \I__2389\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16431\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__16436\,
            I => \N__16428\
        );

    \I__2387\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16425\
        );

    \I__2386\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16422\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__16431\,
            I => \c0.data_in_field_22\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__16428\,
            I => \c0.data_in_field_22\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__16425\,
            I => \c0.data_in_field_22\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__16422\,
            I => \c0.data_in_field_22\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__16413\,
            I => \N__16408\
        );

    \I__2380\ : InMux
    port map (
            O => \N__16412\,
            I => \N__16405\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__16411\,
            I => \N__16401\
        );

    \I__2378\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16398\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__16405\,
            I => \N__16395\
        );

    \I__2376\ : InMux
    port map (
            O => \N__16404\,
            I => \N__16390\
        );

    \I__2375\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16390\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__16398\,
            I => \c0.data_in_field_14\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__16395\,
            I => \c0.data_in_field_14\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__16390\,
            I => \c0.data_in_field_14\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__16383\,
            I => \c0.n9638_cascade_\
        );

    \I__2370\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16375\
        );

    \I__2369\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16372\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__16378\,
            I => \N__16368\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__16375\,
            I => \N__16365\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16362\
        );

    \I__2365\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16359\
        );

    \I__2364\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16355\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__16365\,
            I => \N__16352\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__16362\,
            I => \N__16347\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__16359\,
            I => \N__16347\
        );

    \I__2360\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16344\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__16355\,
            I => \c0.data_in_field_6\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__16352\,
            I => \c0.data_in_field_6\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__16347\,
            I => \c0.data_in_field_6\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__16344\,
            I => \c0.data_in_field_6\
        );

    \I__2355\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16332\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__16332\,
            I => \N__16329\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__16329\,
            I => \N__16325\
        );

    \I__2352\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16322\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__16325\,
            I => data_in_15_4
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__16322\,
            I => data_in_15_4
        );

    \I__2349\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16313\
        );

    \I__2348\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16310\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__16313\,
            I => data_in_17_4
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__16310\,
            I => data_in_17_4
        );

    \I__2345\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16299\
        );

    \I__2344\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16299\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__16299\,
            I => data_in_16_4
        );

    \I__2342\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16290\
        );

    \I__2341\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16290\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__16290\,
            I => data_in_17_7
        );

    \I__2339\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16283\
        );

    \I__2338\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16280\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__16283\,
            I => data_in_19_4
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__16280\,
            I => data_in_19_4
        );

    \I__2335\ : InMux
    port map (
            O => \N__16275\,
            I => \N__16271\
        );

    \I__2334\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16268\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__16271\,
            I => data_in_18_4
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__16268\,
            I => data_in_18_4
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__16263\,
            I => \N__16259\
        );

    \I__2330\ : InMux
    port map (
            O => \N__16262\,
            I => \N__16256\
        );

    \I__2329\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16251\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__16256\,
            I => \N__16248\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__16255\,
            I => \N__16245\
        );

    \I__2326\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16242\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__16251\,
            I => \N__16239\
        );

    \I__2324\ : Span4Mux_h
    port map (
            O => \N__16248\,
            I => \N__16236\
        );

    \I__2323\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16233\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__16242\,
            I => data_in_2_5
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__16239\,
            I => data_in_2_5
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__16236\,
            I => data_in_2_5
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__16233\,
            I => data_in_2_5
        );

    \I__2318\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16221\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__16221\,
            I => \N__16216\
        );

    \I__2316\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16211\
        );

    \I__2315\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16211\
        );

    \I__2314\ : Span4Mux_h
    port map (
            O => \N__16216\,
            I => \N__16208\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__16211\,
            I => data_in_5_6
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__16208\,
            I => data_in_5_6
        );

    \I__2311\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16200\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__16200\,
            I => \N__16197\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__16197\,
            I => \N__16192\
        );

    \I__2308\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16189\
        );

    \I__2307\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16186\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__16192\,
            I => data_in_4_6
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__16189\,
            I => data_in_4_6
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__16186\,
            I => data_in_4_6
        );

    \I__2303\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16174\
        );

    \I__2302\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16166\
        );

    \I__2301\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16166\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16163\
        );

    \I__2299\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16158\
        );

    \I__2298\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16158\
        );

    \I__2297\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16155\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__16166\,
            I => \r_Bit_Index_0_adj_1743\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__16163\,
            I => \r_Bit_Index_0_adj_1743\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__16158\,
            I => \r_Bit_Index_0_adj_1743\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__16155\,
            I => \r_Bit_Index_0_adj_1743\
        );

    \I__2292\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16139\
        );

    \I__2291\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16139\
        );

    \I__2290\ : InMux
    port map (
            O => \N__16144\,
            I => \N__16136\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__16139\,
            I => \N__16133\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__16136\,
            I => n9075
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__16133\,
            I => n9075
        );

    \I__2286\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16122\
        );

    \I__2285\ : InMux
    port map (
            O => \N__16127\,
            I => \N__16122\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16118\
        );

    \I__2283\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16115\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__16118\,
            I => n5346
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__16115\,
            I => n5346
        );

    \I__2280\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16104\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__16109\,
            I => \N__16099\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__16108\,
            I => \N__16096\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__16107\,
            I => \N__16092\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__16104\,
            I => \N__16089\
        );

    \I__2275\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16082\
        );

    \I__2274\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16082\
        );

    \I__2273\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16082\
        );

    \I__2272\ : InMux
    port map (
            O => \N__16096\,
            I => \N__16075\
        );

    \I__2271\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16075\
        );

    \I__2270\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16075\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__16089\,
            I => \r_Bit_Index_1_adj_1742\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__16082\,
            I => \r_Bit_Index_1_adj_1742\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__16075\,
            I => \r_Bit_Index_1_adj_1742\
        );

    \I__2266\ : InMux
    port map (
            O => \N__16068\,
            I => \N__16065\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__16065\,
            I => \N__16062\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__16062\,
            I => \N__16058\
        );

    \I__2263\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16055\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__16058\,
            I => data_in_15_1
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__16055\,
            I => data_in_15_1
        );

    \I__2260\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16046\
        );

    \I__2259\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16043\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__16046\,
            I => \N__16040\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__16043\,
            I => \N__16037\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__16040\,
            I => \N__16033\
        );

    \I__2255\ : Span4Mux_h
    port map (
            O => \N__16037\,
            I => \N__16030\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16036\,
            I => \N__16027\
        );

    \I__2253\ : Span4Mux_v
    port map (
            O => \N__16033\,
            I => \N__16024\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__16030\,
            I => data_in_5_4
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__16027\,
            I => data_in_5_4
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__16024\,
            I => data_in_5_4
        );

    \I__2249\ : InMux
    port map (
            O => \N__16017\,
            I => \N__16013\
        );

    \I__2248\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16010\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__16013\,
            I => data_in_17_1
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__16010\,
            I => data_in_17_1
        );

    \I__2245\ : InMux
    port map (
            O => \N__16005\,
            I => \N__16001\
        );

    \I__2244\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15998\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__16001\,
            I => data_in_16_1
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__15998\,
            I => data_in_16_1
        );

    \I__2241\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15989\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15986\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__15989\,
            I => data_in_14_7
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__15986\,
            I => data_in_14_7
        );

    \I__2237\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15975\
        );

    \I__2236\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15975\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__15975\,
            I => data_in_15_7
        );

    \I__2234\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15966\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15966\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__15966\,
            I => data_in_16_7
        );

    \I__2231\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15960\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__15960\,
            I => \c0.n24_adj_1615\
        );

    \I__2229\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15954\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__15954\,
            I => \c0.n34\
        );

    \I__2227\ : InMux
    port map (
            O => \N__15951\,
            I => \N__15947\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__15950\,
            I => \N__15944\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15934\
        );

    \I__2224\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15925\
        );

    \I__2223\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15925\
        );

    \I__2222\ : InMux
    port map (
            O => \N__15942\,
            I => \N__15925\
        );

    \I__2221\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15925\
        );

    \I__2220\ : InMux
    port map (
            O => \N__15940\,
            I => \N__15922\
        );

    \I__2219\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15915\
        );

    \I__2218\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15915\
        );

    \I__2217\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15915\
        );

    \I__2216\ : Odrv12
    port map (
            O => \N__15934\,
            I => \r_SM_Main_1_adj_1739\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__15925\,
            I => \r_SM_Main_1_adj_1739\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__15922\,
            I => \r_SM_Main_1_adj_1739\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__15915\,
            I => \r_SM_Main_1_adj_1739\
        );

    \I__2212\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15903\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__15903\,
            I => n8747
        );

    \I__2210\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15897\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__15897\,
            I => \c0.tx2.r_Tx_Data_7\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__15894\,
            I => \c0.tx2.n9716_cascade_\
        );

    \I__2207\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15888\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__15888\,
            I => \c0.tx2.n9719\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__15885\,
            I => \n4691_cascade_\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__15882\,
            I => \c0.n4574_cascade_\
        );

    \I__2203\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15873\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15873\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__15873\,
            I => \N__15866\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15861\
        );

    \I__2199\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15861\
        );

    \I__2198\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15858\
        );

    \I__2197\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15855\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__15866\,
            I => data_in_field_81
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__15861\,
            I => data_in_field_81
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__15858\,
            I => data_in_field_81
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__15855\,
            I => data_in_field_81
        );

    \I__2192\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15842\
        );

    \I__2191\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15838\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__15842\,
            I => \N__15834\
        );

    \I__2189\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15831\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__15838\,
            I => \N__15828\
        );

    \I__2187\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15823\
        );

    \I__2186\ : Span12Mux_h
    port map (
            O => \N__15834\,
            I => \N__15818\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__15831\,
            I => \N__15818\
        );

    \I__2184\ : Span4Mux_s2_h
    port map (
            O => \N__15828\,
            I => \N__15815\
        );

    \I__2183\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15810\
        );

    \I__2182\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15810\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__15823\,
            I => data_in_field_47
        );

    \I__2180\ : Odrv12
    port map (
            O => \N__15818\,
            I => data_in_field_47
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__15815\,
            I => data_in_field_47
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__15810\,
            I => data_in_field_47
        );

    \I__2177\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15798\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__15798\,
            I => \c0.n4333\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__15795\,
            I => \c0.n4333_cascade_\
        );

    \I__2174\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15789\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__15789\,
            I => n3_adj_1749
        );

    \I__2172\ : IoInMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__15783\,
            I => \N__15779\
        );

    \I__2170\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15776\
        );

    \I__2169\ : IoSpan4Mux
    port map (
            O => \N__15779\,
            I => \N__15773\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__15776\,
            I => \N__15770\
        );

    \I__2167\ : Span4Mux_s3_h
    port map (
            O => \N__15773\,
            I => \N__15764\
        );

    \I__2166\ : Span4Mux_s3_h
    port map (
            O => \N__15770\,
            I => \N__15764\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15761\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__15764\,
            I => tx2_o
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__15761\,
            I => tx2_o
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__15756\,
            I => \c0.n8788_cascade_\
        );

    \I__2161\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15750\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__15750\,
            I => \c0.n14_adj_1648\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__2158\ : InMux
    port map (
            O => \N__15744\,
            I => \N__15741\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__15741\,
            I => \N__15737\
        );

    \I__2156\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15734\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__15737\,
            I => \c0.n8936\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__15734\,
            I => \c0.n8936\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__15729\,
            I => \c0.n24_adj_1600_cascade_\
        );

    \I__2152\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15723\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__15723\,
            I => \c0.n18_adj_1603\
        );

    \I__2150\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15716\
        );

    \I__2149\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15713\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15710\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__15713\,
            I => \N__15707\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__15710\,
            I => \c0.n4107\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__15707\,
            I => \c0.n4107\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__15702\,
            I => \c0.tx2_transmit_N_1334_cascade_\
        );

    \I__2143\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15696\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__15696\,
            I => \N__15693\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__15693\,
            I => \c0.n8980\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__15690\,
            I => \c0.n22_adj_1601_cascade_\
        );

    \I__2139\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__15684\,
            I => \c0.n26\
        );

    \I__2137\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15678\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__15678\,
            I => \N__15675\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__15675\,
            I => \N__15672\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__15672\,
            I => \c0.n16\
        );

    \I__2133\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15663\
        );

    \I__2132\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15660\
        );

    \I__2131\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15655\
        );

    \I__2130\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15655\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__15663\,
            I => \N__15652\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__15660\,
            I => data_in_field_115
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__15655\,
            I => data_in_field_115
        );

    \I__2126\ : Odrv12
    port map (
            O => \N__15652\,
            I => data_in_field_115
        );

    \I__2125\ : InMux
    port map (
            O => \N__15645\,
            I => \N__15642\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__15642\,
            I => \c0.n4452\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__15639\,
            I => \c0.n4253_cascade_\
        );

    \I__2122\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15632\
        );

    \I__2121\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15629\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__15632\,
            I => \N__15626\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15621\
        );

    \I__2118\ : Span4Mux_s2_v
    port map (
            O => \N__15626\,
            I => \N__15618\
        );

    \I__2117\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15613\
        );

    \I__2116\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15613\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__15621\,
            I => data_in_field_71
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__15618\,
            I => data_in_field_71
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__15613\,
            I => data_in_field_71
        );

    \I__2112\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15599\
        );

    \I__2111\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15599\
        );

    \I__2110\ : InMux
    port map (
            O => \N__15604\,
            I => \N__15596\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__15599\,
            I => \N__15591\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__15596\,
            I => \N__15588\
        );

    \I__2107\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15585\
        );

    \I__2106\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15582\
        );

    \I__2105\ : Span4Mux_v
    port map (
            O => \N__15591\,
            I => \N__15575\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__15588\,
            I => \N__15575\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__15585\,
            I => \N__15575\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__15582\,
            I => data_in_field_147
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__15575\,
            I => data_in_field_147
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__15570\,
            I => \N__15565\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__15569\,
            I => \N__15562\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__15568\,
            I => \N__15559\
        );

    \I__2097\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15555\
        );

    \I__2096\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15550\
        );

    \I__2095\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15550\
        );

    \I__2094\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15547\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15542\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__15550\,
            I => \N__15542\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__15547\,
            I => data_in_field_127
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__15542\,
            I => data_in_field_127
        );

    \I__2089\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15534\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__15534\,
            I => \c0.n9650\
        );

    \I__2087\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15528\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__2085\ : Span4Mux_s3_h
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__15522\,
            I => \c0.n16_adj_1598\
        );

    \I__2083\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15515\
        );

    \I__2082\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15512\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__15515\,
            I => \N__15509\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__15512\,
            I => \N__15506\
        );

    \I__2079\ : Span4Mux_s2_h
    port map (
            O => \N__15509\,
            I => \N__15501\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__15506\,
            I => \N__15501\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__15501\,
            I => \c0.n9016\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__15498\,
            I => \c0.n6_adj_1645_cascade_\
        );

    \I__2075\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15492\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__15492\,
            I => \N__15488\
        );

    \I__2073\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15485\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__15488\,
            I => \N__15480\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__15485\,
            I => \N__15480\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__15480\,
            I => \c0.n4154\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__15477\,
            I => \c0.n10_adj_1640_cascade_\
        );

    \I__2068\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15471\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__15468\,
            I => \N__15465\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__15465\,
            I => \c0.n4434\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__15462\,
            I => \c0.n8933_cascade_\
        );

    \I__2063\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15455\
        );

    \I__2062\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15452\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__15455\,
            I => \N__15449\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__15452\,
            I => \c0.n8822\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__15449\,
            I => \c0.n8822\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__15444\,
            I => \c0.n8314_cascade_\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__15441\,
            I => \N__15437\
        );

    \I__2056\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15431\
        );

    \I__2055\ : InMux
    port map (
            O => \N__15437\,
            I => \N__15431\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__15436\,
            I => \N__15428\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__15431\,
            I => \N__15425\
        );

    \I__2052\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15422\
        );

    \I__2051\ : Span4Mux_h
    port map (
            O => \N__15425\,
            I => \N__15416\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__15422\,
            I => \N__15416\
        );

    \I__2049\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15411\
        );

    \I__2048\ : Span4Mux_v
    port map (
            O => \N__15416\,
            I => \N__15408\
        );

    \I__2047\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15403\
        );

    \I__2046\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15403\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__15411\,
            I => \N__15400\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__15408\,
            I => data_in_field_145
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__15403\,
            I => data_in_field_145
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__15400\,
            I => data_in_field_145
        );

    \I__2041\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15390\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15387\
        );

    \I__2039\ : Span4Mux_s3_h
    port map (
            O => \N__15387\,
            I => \N__15383\
        );

    \I__2038\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15380\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__15383\,
            I => \c0.n4556\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__15380\,
            I => \c0.n4556\
        );

    \I__2035\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15372\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__15372\,
            I => \N__15368\
        );

    \I__2033\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15365\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__15368\,
            I => \c0.n8861\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__15365\,
            I => \c0.n8861\
        );

    \I__2030\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15357\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__15357\,
            I => \c0.n6\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__15354\,
            I => \c0.n4452_cascade_\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__15351\,
            I => \N__15347\
        );

    \I__2026\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15344\
        );

    \I__2025\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15341\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__15344\,
            I => \N__15338\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__15341\,
            I => \N__15335\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__15338\,
            I => \N__15330\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__15335\,
            I => \N__15330\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__15330\,
            I => \c0.n8906\
        );

    \I__2019\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15324\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__15321\,
            I => \N__15318\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__15318\,
            I => n1892
        );

    \I__2015\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15312\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__15312\,
            I => \N__15309\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__15309\,
            I => \N__15306\
        );

    \I__2012\ : Span4Mux_s0_h
    port map (
            O => \N__15306\,
            I => \N__15303\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__15303\,
            I => n1891
        );

    \I__2010\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15297\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__15297\,
            I => \c0.n8831\
        );

    \I__2008\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15288\
        );

    \I__2007\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15285\
        );

    \I__2006\ : InMux
    port map (
            O => \N__15292\,
            I => \N__15282\
        );

    \I__2005\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15279\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__15288\,
            I => \c0.data_in_field_9\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__15285\,
            I => \c0.data_in_field_9\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__15282\,
            I => \c0.data_in_field_9\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__15279\,
            I => \c0.data_in_field_9\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__15270\,
            I => \c0.n8831_cascade_\
        );

    \I__1999\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15264\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__1997\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15255\
        );

    \I__1996\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15252\
        );

    \I__1995\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15249\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__15258\,
            I => \N__15244\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__15255\,
            I => \N__15244\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__15252\,
            I => \N__15239\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__15249\,
            I => \N__15239\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__15244\,
            I => \N__15236\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__15239\,
            I => data_in_1_0
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__15236\,
            I => data_in_1_0
        );

    \I__1987\ : InMux
    port map (
            O => \N__15231\,
            I => \N__15228\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__15228\,
            I => \N__15225\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__15225\,
            I => \N__15222\
        );

    \I__1984\ : Span4Mux_s1_h
    port map (
            O => \N__15222\,
            I => \N__15219\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__15219\,
            I => n1888
        );

    \I__1982\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15212\
        );

    \I__1981\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15208\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__15212\,
            I => \N__15205\
        );

    \I__1979\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15202\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__15208\,
            I => \N__15199\
        );

    \I__1977\ : Odrv12
    port map (
            O => \N__15205\,
            I => data_in_5_3
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__15202\,
            I => data_in_5_3
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__15199\,
            I => data_in_5_3
        );

    \I__1974\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15189\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__15189\,
            I => \N__15186\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__15186\,
            I => \N__15182\
        );

    \I__1971\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15179\
        );

    \I__1970\ : Span4Mux_s2_h
    port map (
            O => \N__15182\,
            I => \N__15175\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__15179\,
            I => \N__15172\
        );

    \I__1968\ : InMux
    port map (
            O => \N__15178\,
            I => \N__15169\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__15175\,
            I => data_in_4_3
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__15172\,
            I => data_in_4_3
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__15169\,
            I => data_in_4_3
        );

    \I__1964\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15157\
        );

    \I__1963\ : InMux
    port map (
            O => \N__15161\,
            I => \N__15154\
        );

    \I__1962\ : InMux
    port map (
            O => \N__15160\,
            I => \N__15151\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__15157\,
            I => \c0.n4131\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__15154\,
            I => \c0.n4131\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__15151\,
            I => \c0.n4131\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__15144\,
            I => \N__15141\
        );

    \I__1957\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15138\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__15138\,
            I => \N__15133\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15130\
        );

    \I__1954\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15127\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__15133\,
            I => \N__15124\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__15130\,
            I => \c0.n4224\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__15127\,
            I => \c0.n4224\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__15124\,
            I => \c0.n4224\
        );

    \I__1949\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15114\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__15114\,
            I => \N__15111\
        );

    \I__1947\ : Odrv12
    port map (
            O => \N__15111\,
            I => \c0.n4127\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__15108\,
            I => \N__15105\
        );

    \I__1945\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15102\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__15102\,
            I => \N__15097\
        );

    \I__1943\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15092\
        );

    \I__1942\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15092\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__15097\,
            I => data_in_0_3
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__15092\,
            I => data_in_0_3
        );

    \I__1939\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15081\
        );

    \I__1938\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15078\
        );

    \I__1937\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15075\
        );

    \I__1936\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15072\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__15081\,
            I => \N__15069\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__15078\,
            I => \N__15064\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__15075\,
            I => \N__15064\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__15072\,
            I => \N__15058\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__15069\,
            I => \N__15058\
        );

    \I__1930\ : Span4Mux_s3_h
    port map (
            O => \N__15064\,
            I => \N__15055\
        );

    \I__1929\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15052\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__15058\,
            I => \c0.data_in_field_3\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__15055\,
            I => \c0.data_in_field_3\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__15052\,
            I => \c0.data_in_field_3\
        );

    \I__1925\ : InMux
    port map (
            O => \N__15045\,
            I => \N__15042\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__15042\,
            I => \N__15039\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__15039\,
            I => \c0.n20_adj_1597\
        );

    \I__1922\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15033\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__15033\,
            I => \N__15030\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__15030\,
            I => \c0.n22_adj_1595\
        );

    \I__1919\ : InMux
    port map (
            O => \N__15027\,
            I => \N__15023\
        );

    \I__1918\ : InMux
    port map (
            O => \N__15026\,
            I => \N__15019\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__15023\,
            I => \N__15015\
        );

    \I__1916\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15012\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__15019\,
            I => \N__15009\
        );

    \I__1914\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15006\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__15015\,
            I => data_in_2_6
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__15012\,
            I => data_in_2_6
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__15009\,
            I => data_in_2_6
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__15006\,
            I => data_in_2_6
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__14997\,
            I => \n9069_cascade_\
        );

    \I__1908\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14990\
        );

    \I__1907\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14986\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__14990\,
            I => \N__14982\
        );

    \I__1905\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14979\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__14986\,
            I => \N__14976\
        );

    \I__1903\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14973\
        );

    \I__1902\ : Span4Mux_s3_h
    port map (
            O => \N__14982\,
            I => \N__14970\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14965\
        );

    \I__1900\ : Span4Mux_s3_h
    port map (
            O => \N__14976\,
            I => \N__14965\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__14973\,
            I => data_in_3_3
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__14970\,
            I => data_in_3_3
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__14965\,
            I => data_in_3_3
        );

    \I__1896\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14955\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14952\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__14952\,
            I => \c0.n8849\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__14949\,
            I => \n4_adj_1750_cascade_\
        );

    \I__1892\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14943\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__14943\,
            I => \N__14938\
        );

    \I__1890\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14935\
        );

    \I__1889\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14931\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__14938\,
            I => \N__14928\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14925\
        );

    \I__1886\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14922\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__14931\,
            I => \c0.data_in_field_2\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__14928\,
            I => \c0.data_in_field_2\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__14925\,
            I => \c0.data_in_field_2\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__14922\,
            I => \c0.data_in_field_2\
        );

    \I__1881\ : InMux
    port map (
            O => \N__14913\,
            I => \N__14909\
        );

    \I__1880\ : InMux
    port map (
            O => \N__14912\,
            I => \N__14906\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__14909\,
            I => \N__14902\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__14906\,
            I => \N__14899\
        );

    \I__1877\ : InMux
    port map (
            O => \N__14905\,
            I => \N__14894\
        );

    \I__1876\ : Span4Mux_s3_h
    port map (
            O => \N__14902\,
            I => \N__14889\
        );

    \I__1875\ : Span4Mux_s3_h
    port map (
            O => \N__14899\,
            I => \N__14889\
        );

    \I__1874\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14886\
        );

    \I__1873\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14883\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__14894\,
            I => \c0.data_in_field_33\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__14889\,
            I => \c0.data_in_field_33\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__14886\,
            I => \c0.data_in_field_33\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__14883\,
            I => \c0.data_in_field_33\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__14874\,
            I => \c0.n6_adj_1632_cascade_\
        );

    \I__1867\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14868\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__14868\,
            I => \c0.n8804\
        );

    \I__1865\ : InMux
    port map (
            O => \N__14865\,
            I => \N__14862\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__14862\,
            I => \N__14858\
        );

    \I__1863\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14853\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__14858\,
            I => \N__14850\
        );

    \I__1861\ : InMux
    port map (
            O => \N__14857\,
            I => \N__14847\
        );

    \I__1860\ : InMux
    port map (
            O => \N__14856\,
            I => \N__14844\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__14853\,
            I => data_in_1_6
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__14850\,
            I => data_in_1_6
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__14847\,
            I => data_in_1_6
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__14844\,
            I => data_in_1_6
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__14835\,
            I => \N__14832\
        );

    \I__1854\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14827\
        );

    \I__1853\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14824\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__14830\,
            I => \N__14821\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__14827\,
            I => \N__14817\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__14824\,
            I => \N__14814\
        );

    \I__1849\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14809\
        );

    \I__1848\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14809\
        );

    \I__1847\ : Span4Mux_h
    port map (
            O => \N__14817\,
            I => \N__14806\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__14814\,
            I => \N__14803\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__14809\,
            I => data_in_3_7
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__14806\,
            I => data_in_3_7
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__14803\,
            I => data_in_3_7
        );

    \I__1842\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14793\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__14793\,
            I => \N__14789\
        );

    \I__1840\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14786\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__14789\,
            I => data_in_13_0
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__14786\,
            I => data_in_13_0
        );

    \I__1837\ : InMux
    port map (
            O => \N__14781\,
            I => \N__14778\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__14778\,
            I => \N__14773\
        );

    \I__1835\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14770\
        );

    \I__1834\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14767\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__14773\,
            I => data_in_4_0
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__14770\,
            I => data_in_4_0
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__14767\,
            I => data_in_4_0
        );

    \I__1830\ : InMux
    port map (
            O => \N__14760\,
            I => \N__14757\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__14757\,
            I => \c0.n13_adj_1671\
        );

    \I__1828\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14751\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__14751\,
            I => \c0.n13_adj_1672\
        );

    \I__1826\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14744\
        );

    \I__1825\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14741\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__14744\,
            I => \N__14737\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14734\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__14740\,
            I => \N__14730\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__14737\,
            I => \N__14727\
        );

    \I__1820\ : Span4Mux_s3_h
    port map (
            O => \N__14734\,
            I => \N__14724\
        );

    \I__1819\ : InMux
    port map (
            O => \N__14733\,
            I => \N__14721\
        );

    \I__1818\ : InMux
    port map (
            O => \N__14730\,
            I => \N__14718\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__14727\,
            I => data_in_1_2
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__14724\,
            I => data_in_1_2
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__14721\,
            I => data_in_1_2
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__14718\,
            I => data_in_1_2
        );

    \I__1813\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14706\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__14706\,
            I => \N__14701\
        );

    \I__1811\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14696\
        );

    \I__1810\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14696\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__14701\,
            I => data_in_6_3
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__14696\,
            I => data_in_6_3
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__14691\,
            I => \N__14688\
        );

    \I__1806\ : InMux
    port map (
            O => \N__14688\,
            I => \N__14685\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__14685\,
            I => \N__14682\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__14682\,
            I => \N__14676\
        );

    \I__1803\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14669\
        );

    \I__1802\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14669\
        );

    \I__1801\ : InMux
    port map (
            O => \N__14679\,
            I => \N__14669\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__14676\,
            I => data_in_1_3
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__14669\,
            I => data_in_1_3
        );

    \I__1798\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14661\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__14661\,
            I => \N__14657\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__14660\,
            I => \N__14654\
        );

    \I__1795\ : Span4Mux_s3_h
    port map (
            O => \N__14657\,
            I => \N__14649\
        );

    \I__1794\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14642\
        );

    \I__1793\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14642\
        );

    \I__1792\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14642\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__14649\,
            I => data_in_2_3
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__14642\,
            I => data_in_2_3
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__14637\,
            I => \N__14634\
        );

    \I__1788\ : InMux
    port map (
            O => \N__14634\,
            I => \N__14631\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__14631\,
            I => \N__14628\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__14628\,
            I => \c0.n4495\
        );

    \I__1785\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14621\
        );

    \I__1784\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14618\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__14621\,
            I => data_in_15_6
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__14618\,
            I => data_in_15_6
        );

    \I__1781\ : InMux
    port map (
            O => \N__14613\,
            I => \N__14609\
        );

    \I__1780\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14606\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__14609\,
            I => data_in_14_6
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__14606\,
            I => data_in_14_6
        );

    \I__1777\ : InMux
    port map (
            O => \N__14601\,
            I => \N__14597\
        );

    \I__1776\ : InMux
    port map (
            O => \N__14600\,
            I => \N__14594\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__14597\,
            I => data_in_20_4
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__14594\,
            I => data_in_20_4
        );

    \I__1773\ : InMux
    port map (
            O => \N__14589\,
            I => \N__14585\
        );

    \I__1772\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14580\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__14585\,
            I => \N__14577\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__14584\,
            I => \N__14574\
        );

    \I__1769\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14571\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__14580\,
            I => \N__14566\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__14577\,
            I => \N__14566\
        );

    \I__1766\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14563\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__14571\,
            I => data_in_3_0
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__14566\,
            I => data_in_3_0
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__14563\,
            I => data_in_3_0
        );

    \I__1762\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14552\
        );

    \I__1761\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14548\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__14552\,
            I => \N__14545\
        );

    \I__1759\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14542\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__14548\,
            I => data_in_0_5
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__14545\,
            I => data_in_0_5
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__14542\,
            I => data_in_0_5
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__14535\,
            I => \c0.n28_adj_1668_cascade_\
        );

    \I__1754\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14529\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__14529\,
            I => \c0.n30_adj_1674\
        );

    \I__1752\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14523\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__14523\,
            I => \c0.n22_adj_1667\
        );

    \I__1750\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14517\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__14517\,
            I => \N__14514\
        );

    \I__1748\ : Span4Mux_s3_h
    port map (
            O => \N__14514\,
            I => \N__14509\
        );

    \I__1747\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14504\
        );

    \I__1746\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14504\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__14509\,
            I => data_in_0_0
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__14504\,
            I => data_in_0_0
        );

    \I__1743\ : InMux
    port map (
            O => \N__14499\,
            I => \N__14496\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__14496\,
            I => \N__14493\
        );

    \I__1741\ : Span4Mux_s3_h
    port map (
            O => \N__14493\,
            I => \N__14489\
        );

    \I__1740\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14486\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__14489\,
            I => data_in_13_7
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__14486\,
            I => data_in_13_7
        );

    \I__1737\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14475\
        );

    \I__1736\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14475\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__14475\,
            I => data_in_16_6
        );

    \I__1734\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14468\
        );

    \I__1733\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14465\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__14468\,
            I => data_in_9_6
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__14465\,
            I => data_in_9_6
        );

    \I__1730\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14454\
        );

    \I__1729\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14454\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__14454\,
            I => data_in_10_6
        );

    \I__1727\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14445\
        );

    \I__1726\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14445\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__14445\,
            I => data_in_11_6
        );

    \I__1724\ : InMux
    port map (
            O => \N__14442\,
            I => \N__14438\
        );

    \I__1723\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14435\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__14438\,
            I => data_in_13_6
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__14435\,
            I => data_in_13_6
        );

    \I__1720\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14424\
        );

    \I__1719\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14424\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__14424\,
            I => data_in_12_6
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__14421\,
            I => \c0.n9752_cascade_\
        );

    \I__1716\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14414\
        );

    \I__1715\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14410\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__14414\,
            I => \N__14406\
        );

    \I__1713\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14403\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__14410\,
            I => \N__14400\
        );

    \I__1711\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14396\
        );

    \I__1710\ : Span12Mux_s3_v
    port map (
            O => \N__14406\,
            I => \N__14393\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__14403\,
            I => \N__14388\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__14400\,
            I => \N__14388\
        );

    \I__1707\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14385\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__14396\,
            I => \c0.data_in_field_39\
        );

    \I__1705\ : Odrv12
    port map (
            O => \N__14393\,
            I => \c0.data_in_field_39\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__14388\,
            I => \c0.data_in_field_39\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__14385\,
            I => \c0.data_in_field_39\
        );

    \I__1702\ : InMux
    port map (
            O => \N__14376\,
            I => \N__14373\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__14373\,
            I => \c0.n9120\
        );

    \I__1700\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14367\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__14367\,
            I => \N__14364\
        );

    \I__1698\ : Span4Mux_s2_v
    port map (
            O => \N__14364\,
            I => \N__14361\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__14361\,
            I => \c0.tx2.r_Tx_Data_3\
        );

    \I__1696\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14355\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__14355\,
            I => \N__14352\
        );

    \I__1694\ : Span4Mux_h
    port map (
            O => \N__14352\,
            I => \N__14349\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__14349\,
            I => \c0.tx2.r_Tx_Data_1\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__14346\,
            I => \c0.tx2.n9692_cascade_\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__14343\,
            I => \c0.tx2.n9695_cascade_\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__14340\,
            I => \c0.tx2.o_Tx_Serial_N_1511_cascade_\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__14337\,
            I => \n2207_cascade_\
        );

    \I__1688\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14327\
        );

    \I__1687\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14327\
        );

    \I__1686\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14324\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__14327\,
            I => \r_Bit_Index_2_adj_1741\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__14324\,
            I => \r_Bit_Index_2_adj_1741\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__14319\,
            I => \N__14311\
        );

    \I__1682\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14308\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__14317\,
            I => \N__14305\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__14316\,
            I => \N__14301\
        );

    \I__1679\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14292\
        );

    \I__1678\ : InMux
    port map (
            O => \N__14314\,
            I => \N__14292\
        );

    \I__1677\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14292\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__14308\,
            I => \N__14289\
        );

    \I__1675\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14284\
        );

    \I__1674\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14284\
        );

    \I__1673\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14277\
        );

    \I__1672\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14277\
        );

    \I__1671\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14277\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__14292\,
            I => \r_SM_Main_0_adj_1740\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__14289\,
            I => \r_SM_Main_0_adj_1740\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__14284\,
            I => \r_SM_Main_0_adj_1740\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__14277\,
            I => \r_SM_Main_0_adj_1740\
        );

    \I__1666\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14261\
        );

    \I__1665\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14252\
        );

    \I__1664\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14252\
        );

    \I__1663\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14252\
        );

    \I__1662\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14252\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__14261\,
            I => \r_SM_Main_2_N_1480_1_adj_1744\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__14252\,
            I => \r_SM_Main_2_N_1480_1_adj_1744\
        );

    \I__1659\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14241\
        );

    \I__1658\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14238\
        );

    \I__1657\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14233\
        );

    \I__1656\ : InMux
    port map (
            O => \N__14244\,
            I => \N__14233\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14230\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__14238\,
            I => data_in_field_83
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__14233\,
            I => data_in_field_83
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__14230\,
            I => data_in_field_83
        );

    \I__1651\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14220\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__14220\,
            I => \N__14217\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__14217\,
            I => \c0.n9126\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__14214\,
            I => \c0.n9123_cascade_\
        );

    \I__1647\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14208\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__14208\,
            I => \N__14205\
        );

    \I__1645\ : Span4Mux_s2_v
    port map (
            O => \N__14205\,
            I => \N__14202\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__14202\,
            I => \c0.n9240\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__14199\,
            I => \c0.n9644_cascade_\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__14196\,
            I => \c0.n9647_cascade_\
        );

    \I__1641\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14190\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__14190\,
            I => \c0.n9656\
        );

    \I__1639\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14184\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__14184\,
            I => n6164
        );

    \I__1637\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14178\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__14178\,
            I => \N__14173\
        );

    \I__1635\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14168\
        );

    \I__1634\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14168\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__14173\,
            I => data_in_field_105
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__14168\,
            I => data_in_field_105
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__14163\,
            I => \c0.n8890_cascade_\
        );

    \I__1630\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14157\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__14157\,
            I => \N__14154\
        );

    \I__1628\ : Span4Mux_h
    port map (
            O => \N__14154\,
            I => \N__14151\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__14151\,
            I => \N__14148\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__14148\,
            I => \c0.n14_adj_1638\
        );

    \I__1625\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14142\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__14142\,
            I => \N__14139\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__14139\,
            I => \c0.n4285\
        );

    \I__1622\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14132\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14129\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__14132\,
            I => \N__14126\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__14129\,
            I => \N__14123\
        );

    \I__1618\ : Odrv12
    port map (
            O => \N__14126\,
            I => \c0.n9007\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__14123\,
            I => \c0.n9007\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__14118\,
            I => \c0.n18_adj_1589_cascade_\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__14115\,
            I => \c0.n20_adj_1590_cascade_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14109\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__14109\,
            I => \N__14105\
        );

    \I__1612\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14102\
        );

    \I__1611\ : Sp12to4
    port map (
            O => \N__14105\,
            I => \N__14097\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__14102\,
            I => \N__14097\
        );

    \I__1609\ : Odrv12
    port map (
            O => \N__14097\,
            I => \c0.n29\
        );

    \I__1608\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14091\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__14091\,
            I => \N__14088\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__14088\,
            I => \c0.n4114\
        );

    \I__1605\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14082\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__14082\,
            I => \c0.n4448\
        );

    \I__1603\ : InMux
    port map (
            O => \N__14079\,
            I => \N__14076\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__14076\,
            I => \c0.n4445\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__14073\,
            I => \N__14070\
        );

    \I__1600\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14067\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__14067\,
            I => \N__14063\
        );

    \I__1598\ : InMux
    port map (
            O => \N__14066\,
            I => \N__14060\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__14063\,
            I => \c0.n8896\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__14060\,
            I => \c0.n8896\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__14055\,
            I => \c0.n10_adj_1647_cascade_\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__14052\,
            I => \N__14049\
        );

    \I__1593\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14046\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__14046\,
            I => \N__14043\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__14043\,
            I => \c0.data_in_frame_19_1\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__14040\,
            I => \c0.n9704_cascade_\
        );

    \I__1589\ : InMux
    port map (
            O => \N__14037\,
            I => \N__14034\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__14034\,
            I => \N__14031\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__14031\,
            I => \N__14028\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__14028\,
            I => \N__14025\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__14025\,
            I => \c0.data_in_frame_20_1\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__14022\,
            I => \c0.n9707_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14016\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__14016\,
            I => \N__14013\
        );

    \I__1581\ : Span4Mux_s3_h
    port map (
            O => \N__14013\,
            I => \N__14010\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__14010\,
            I => \c0.n22_adj_1682\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__14007\,
            I => \c0.n9722_cascade_\
        );

    \I__1578\ : InMux
    port map (
            O => \N__14004\,
            I => \N__14000\
        );

    \I__1577\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13995\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14000\,
            I => \N__13992\
        );

    \I__1575\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13987\
        );

    \I__1574\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13987\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__13995\,
            I => \c0.data_in_field_7\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__13992\,
            I => \c0.data_in_field_7\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__13987\,
            I => \c0.data_in_field_7\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__13980\,
            I => \N__13976\
        );

    \I__1569\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13973\
        );

    \I__1568\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13968\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__13973\,
            I => \N__13965\
        );

    \I__1566\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13960\
        );

    \I__1565\ : InMux
    port map (
            O => \N__13971\,
            I => \N__13960\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__13968\,
            I => \c0.data_in_field_23\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__13965\,
            I => \c0.data_in_field_23\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__13960\,
            I => \c0.data_in_field_23\
        );

    \I__1561\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13949\
        );

    \I__1560\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13946\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__13949\,
            I => \N__13943\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__13946\,
            I => \c0.n4514\
        );

    \I__1557\ : Odrv12
    port map (
            O => \N__13943\,
            I => \c0.n4514\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__1555\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13928\
        );

    \I__1554\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13921\
        );

    \I__1553\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13921\
        );

    \I__1552\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13921\
        );

    \I__1551\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13918\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__13928\,
            I => \N__13913\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__13921\,
            I => \N__13913\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__13918\,
            I => \c0.data_in_field_4\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__13913\,
            I => \c0.data_in_field_4\
        );

    \I__1546\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13905\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__13905\,
            I => \N__13900\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__13904\,
            I => \N__13897\
        );

    \I__1543\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13894\
        );

    \I__1542\ : Span4Mux_v
    port map (
            O => \N__13900\,
            I => \N__13891\
        );

    \I__1541\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13888\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__13894\,
            I => data_in_0_7
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__13891\,
            I => data_in_0_7
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__13888\,
            I => data_in_0_7
        );

    \I__1537\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13878\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__13878\,
            I => \N__13873\
        );

    \I__1535\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13868\
        );

    \I__1534\ : InMux
    port map (
            O => \N__13876\,
            I => \N__13868\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__13873\,
            I => \c0.n8776\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__13868\,
            I => \c0.n8776\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__13863\,
            I => \c0.n4131_cascade_\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__13860\,
            I => \c0.n8927_cascade_\
        );

    \I__1529\ : InMux
    port map (
            O => \N__13857\,
            I => \N__13854\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__13854\,
            I => \N__13851\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__13851\,
            I => \N__13848\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__13848\,
            I => n1896
        );

    \I__1525\ : InMux
    port map (
            O => \N__13845\,
            I => \N__13842\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13842\,
            I => \N__13839\
        );

    \I__1523\ : Span4Mux_h
    port map (
            O => \N__13839\,
            I => \N__13833\
        );

    \I__1522\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13828\
        );

    \I__1521\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13828\
        );

    \I__1520\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13825\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__13833\,
            I => data_in_2_7
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__13828\,
            I => data_in_2_7
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__13825\,
            I => data_in_2_7
        );

    \I__1516\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13814\
        );

    \I__1515\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13810\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__13814\,
            I => \N__13807\
        );

    \I__1513\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13804\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__13810\,
            I => data_in_0_6
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__13807\,
            I => data_in_0_6
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__13804\,
            I => data_in_0_6
        );

    \I__1509\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13793\
        );

    \I__1508\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13787\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__13793\,
            I => \N__13784\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13777\
        );

    \I__1505\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13777\
        );

    \I__1504\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13777\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__13787\,
            I => \c0.data_in_field_19\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__13784\,
            I => \c0.data_in_field_19\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__13777\,
            I => \c0.data_in_field_19\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13767\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__13767\,
            I => \c0.n14\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__13764\,
            I => \c0.n10_adj_1631_cascade_\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13757\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__13760\,
            I => \N__13754\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__13757\,
            I => \N__13749\
        );

    \I__1494\ : InMux
    port map (
            O => \N__13754\,
            I => \N__13742\
        );

    \I__1493\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13742\
        );

    \I__1492\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13742\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__13749\,
            I => data_in_1_1
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__13742\,
            I => data_in_1_1
        );

    \I__1489\ : InMux
    port map (
            O => \N__13737\,
            I => \N__13734\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__13734\,
            I => \N__13730\
        );

    \I__1487\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13727\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__13730\,
            I => \N__13724\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__13727\,
            I => \N__13721\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__13724\,
            I => \N__13717\
        );

    \I__1483\ : Sp12to4
    port map (
            O => \N__13721\,
            I => \N__13714\
        );

    \I__1482\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13711\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__13717\,
            I => data_in_4_7
        );

    \I__1480\ : Odrv12
    port map (
            O => \N__13714\,
            I => data_in_4_7
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__13711\,
            I => data_in_4_7
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__13704\,
            I => \N__13701\
        );

    \I__1477\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13698\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__13698\,
            I => \N__13695\
        );

    \I__1475\ : Span4Mux_s2_h
    port map (
            O => \N__13695\,
            I => \N__13692\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__13692\,
            I => \c0.n47\
        );

    \I__1473\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13686\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__13686\,
            I => \N__13681\
        );

    \I__1471\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13678\
        );

    \I__1470\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13675\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__13681\,
            I => data_in_0_2
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__13678\,
            I => data_in_0_2
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__13675\,
            I => data_in_0_2
        );

    \I__1466\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13665\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__13665\,
            I => \c0.n4381\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__13662\,
            I => \c0.n4381_cascade_\
        );

    \I__1463\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13648\
        );

    \I__1462\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13648\
        );

    \I__1461\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13648\
        );

    \I__1460\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13643\
        );

    \I__1459\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13643\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__13648\,
            I => \c0.data_in_field_20\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__13643\,
            I => \c0.data_in_field_20\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__13638\,
            I => \N__13635\
        );

    \I__1455\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13632\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13629\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__13629\,
            I => \N__13624\
        );

    \I__1452\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13619\
        );

    \I__1451\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13619\
        );

    \I__1450\ : IoSpan4Mux
    port map (
            O => \N__13624\,
            I => \N__13616\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__13619\,
            I => data_in_4_1
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__13616\,
            I => data_in_4_1
        );

    \I__1447\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13607\
        );

    \I__1446\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13601\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__13607\,
            I => \N__13598\
        );

    \I__1444\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13591\
        );

    \I__1443\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13591\
        );

    \I__1442\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13591\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__13601\,
            I => \c0.data_in_field_35\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__13598\,
            I => \c0.data_in_field_35\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__13591\,
            I => \c0.data_in_field_35\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__13584\,
            I => \c0.n4154_cascade_\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__13581\,
            I => \N__13578\
        );

    \I__1436\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13575\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__13575\,
            I => \c0.n9578\
        );

    \I__1434\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13569\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__13569\,
            I => \c0.n8794\
        );

    \I__1432\ : InMux
    port map (
            O => \N__13566\,
            I => \N__13562\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__13565\,
            I => \N__13558\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__13562\,
            I => \N__13554\
        );

    \I__1429\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13549\
        );

    \I__1428\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13549\
        );

    \I__1427\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13546\
        );

    \I__1426\ : Span4Mux_h
    port map (
            O => \N__13554\,
            I => \N__13543\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13540\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__13546\,
            I => data_in_3_1
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__13543\,
            I => data_in_3_1
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__13540\,
            I => data_in_3_1
        );

    \I__1421\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13529\
        );

    \I__1420\ : InMux
    port map (
            O => \N__13532\,
            I => \N__13526\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__13529\,
            I => data_in_9_0
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__13526\,
            I => data_in_9_0
        );

    \I__1417\ : InMux
    port map (
            O => \N__13521\,
            I => \N__13517\
        );

    \I__1416\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13514\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__13517\,
            I => data_in_8_0
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__13514\,
            I => data_in_8_0
        );

    \I__1413\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13503\
        );

    \I__1412\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13503\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__13503\,
            I => data_in_7_0
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__13500\,
            I => \N__13497\
        );

    \I__1409\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13493\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__13496\,
            I => \N__13488\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__13493\,
            I => \N__13485\
        );

    \I__1406\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13482\
        );

    \I__1405\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13477\
        );

    \I__1404\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13477\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__13485\,
            I => data_in_1_5
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__13482\,
            I => data_in_1_5
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__13477\,
            I => data_in_1_5
        );

    \I__1400\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13467\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__13467\,
            I => \N__13463\
        );

    \I__1398\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13460\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__13463\,
            I => data_in_12_0
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__13460\,
            I => data_in_12_0
        );

    \I__1395\ : InMux
    port map (
            O => \N__13455\,
            I => \N__13452\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__13452\,
            I => \N__13449\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__13449\,
            I => \N__13446\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__13446\,
            I => \c0.n14_adj_1670\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__13443\,
            I => \N__13440\
        );

    \I__1390\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13437\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__13437\,
            I => \c0.n14_adj_1669\
        );

    \I__1388\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13431\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__13431\,
            I => \N__13428\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__13428\,
            I => \N__13425\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__13425\,
            I => \c0.n26_adj_1673\
        );

    \I__1384\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13419\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__13419\,
            I => \c0.n25_adj_1675\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__13416\,
            I => \c0.n9033_cascade_\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__13413\,
            I => \n3220_cascade_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13406\
        );

    \I__1379\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13403\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__13406\,
            I => data_in_9_7
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__13403\,
            I => data_in_9_7
        );

    \I__1376\ : InMux
    port map (
            O => \N__13398\,
            I => \N__13394\
        );

    \I__1375\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13391\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__13394\,
            I => data_in_8_7
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__13391\,
            I => data_in_8_7
        );

    \I__1372\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13383\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__13383\,
            I => \N__13380\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__13380\,
            I => \N__13377\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__13377\,
            I => n1900
        );

    \I__1368\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13368\
        );

    \I__1367\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13368\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__13368\,
            I => data_in_7_3
        );

    \I__1365\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13359\
        );

    \I__1364\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13359\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__13359\,
            I => data_in_8_3
        );

    \I__1362\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13352\
        );

    \I__1361\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13349\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__13352\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__13349\,
            I => \c0.tx2.r_Clock_Count_5\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__13344\,
            I => \c0.tx2.n5_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13337\
        );

    \I__1356\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13334\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__13337\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__13334\,
            I => \c0.tx2.r_Clock_Count_7\
        );

    \I__1353\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13326\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__13326\,
            I => \c0.tx2.n4081\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__13323\,
            I => \c0.tx2.n4081_cascade_\
        );

    \I__1350\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13317\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__13317\,
            I => \c0.tx2.n7\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__13314\,
            I => \c0.tx2.n8196_cascade_\
        );

    \I__1347\ : SRMux
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__13308\,
            I => \N__13304\
        );

    \I__1345\ : SRMux
    port map (
            O => \N__13307\,
            I => \N__13301\
        );

    \I__1344\ : Span4Mux_s1_h
    port map (
            O => \N__13304\,
            I => \N__13298\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__13301\,
            I => \N__13295\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__13298\,
            I => \c0.tx2.n5146\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__13295\,
            I => \c0.tx2.n5146\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__13290\,
            I => \n9075_cascade_\
        );

    \I__1339\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13280\
        );

    \I__1338\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13277\
        );

    \I__1337\ : InMux
    port map (
            O => \N__13285\,
            I => \N__13270\
        );

    \I__1336\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13270\
        );

    \I__1335\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13270\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__13280\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__13277\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__13270\,
            I => \c0.tx2.r_Clock_Count_8\
        );

    \I__1331\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13253\
        );

    \I__1330\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13253\
        );

    \I__1329\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13253\
        );

    \I__1328\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13250\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__13253\,
            I => \c0.tx2.n7399\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__13250\,
            I => \c0.tx2.n7399\
        );

    \I__1325\ : InMux
    port map (
            O => \N__13245\,
            I => \N__13242\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__13242\,
            I => \c0.tx2.n7236\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__13239\,
            I => \c0.tx2.n7236_cascade_\
        );

    \I__1322\ : InMux
    port map (
            O => \N__13236\,
            I => \N__13233\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__13230\,
            I => \N__13227\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__13227\,
            I => \c0.n4577\
        );

    \I__1318\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13221\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__13221\,
            I => \c0.n4282\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__13218\,
            I => \c0.n4476_cascade_\
        );

    \I__1315\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13212\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__13212\,
            I => \N__13209\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__13209\,
            I => \N__13206\
        );

    \I__1312\ : Odrv4
    port map (
            O => \N__13206\,
            I => \c0.n19_adj_1623\
        );

    \I__1311\ : InMux
    port map (
            O => \N__13203\,
            I => \N__13199\
        );

    \I__1310\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13196\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__13199\,
            I => \N__13190\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__13196\,
            I => \N__13190\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13187\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__13190\,
            I => \N__13184\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__13187\,
            I => data_in_5_7
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__13184\,
            I => data_in_5_7
        );

    \I__1303\ : IoInMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__13176\,
            I => \N__13173\
        );

    \I__1301\ : Span4Mux_s1_h
    port map (
            O => \N__13173\,
            I => \N__13170\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__13170\,
            I => tx2_enable
        );

    \I__1299\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13163\
        );

    \I__1298\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13160\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__13163\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__13160\,
            I => \c0.tx2.r_Clock_Count_2\
        );

    \I__1295\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13151\
        );

    \I__1294\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13148\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__13151\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__13148\,
            I => \c0.tx2.r_Clock_Count_6\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__13143\,
            I => \N__13139\
        );

    \I__1290\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13136\
        );

    \I__1289\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13133\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__13136\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__13133\,
            I => \c0.tx2.r_Clock_Count_1\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13124\
        );

    \I__1285\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13121\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__13124\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__13121\,
            I => \c0.tx2.r_Clock_Count_3\
        );

    \I__1282\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13112\
        );

    \I__1281\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13109\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13112\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__13109\,
            I => \c0.tx2.r_Clock_Count_4\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__13104\,
            I => \c0.n4568_cascade_\
        );

    \I__1277\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13098\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__13098\,
            I => \c0.n46\
        );

    \I__1275\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13091\
        );

    \I__1274\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13088\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__13091\,
            I => \N__13084\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__13088\,
            I => \N__13081\
        );

    \I__1271\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13078\
        );

    \I__1270\ : Span12Mux_s1_h
    port map (
            O => \N__13084\,
            I => \N__13073\
        );

    \I__1269\ : Span12Mux_s5_v
    port map (
            O => \N__13081\,
            I => \N__13073\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__13078\,
            I => data_in_6_7
        );

    \I__1267\ : Odrv12
    port map (
            O => \N__13073\,
            I => data_in_6_7
        );

    \I__1266\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13065\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__13065\,
            I => \c0.n8816\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__13062\,
            I => \c0.n4282_cascade_\
        );

    \I__1263\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13056\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__13053\
        );

    \I__1261\ : Span4Mux_s2_h
    port map (
            O => \N__13053\,
            I => \N__13050\
        );

    \I__1260\ : Span4Mux_h
    port map (
            O => \N__13050\,
            I => \N__13047\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__13047\,
            I => \c0.data_in_frame_20_5\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__13044\,
            I => \c0.n4215_cascade_\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__13041\,
            I => \c0.n18_adj_1593_cascade_\
        );

    \I__1256\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13035\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__13035\,
            I => \c0.n20_adj_1596\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__13032\,
            I => \c0.n17_cascade_\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__13029\,
            I => \c0.n4324_cascade_\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13026\,
            I => \N__13023\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__13023\,
            I => \c0.n8951\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__13020\,
            I => \c0.n8951_cascade_\
        );

    \I__1249\ : InMux
    port map (
            O => \N__13017\,
            I => \N__13014\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__13014\,
            I => \N__13011\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__13011\,
            I => \c0.n48\
        );

    \I__1246\ : InMux
    port map (
            O => \N__13008\,
            I => \N__13005\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__13005\,
            I => \c0.n4406\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__13002\,
            I => \c0.n4406_cascade_\
        );

    \I__1243\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12996\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__12996\,
            I => \N__12993\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__12993\,
            I => \c0.n43_adj_1610\
        );

    \I__1240\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12987\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12984\
        );

    \I__1238\ : Span4Mux_h
    port map (
            O => \N__12984\,
            I => \N__12981\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__12981\,
            I => n1894
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__12978\,
            I => \c0.n9542_cascade_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12972\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__12972\,
            I => \N__12969\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__12969\,
            I => \N__12966\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__12966\,
            I => \c0.n9180\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \c0.n4114_cascade_\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__12960\,
            I => \c0.n8801_cascade_\
        );

    \I__1229\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12954\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__12954\,
            I => \N__12948\
        );

    \I__1227\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12941\
        );

    \I__1226\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12941\
        );

    \I__1225\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12941\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__12948\,
            I => \c0.data_in_field_11\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__12941\,
            I => \c0.data_in_field_11\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__12936\,
            I => \N__12933\
        );

    \I__1221\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12930\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__12930\,
            I => \c0.n4276\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__12927\,
            I => \c0.n4276_cascade_\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__12924\,
            I => \c0.n12_adj_1633_cascade_\
        );

    \I__1217\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12917\
        );

    \I__1216\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12914\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__12917\,
            I => \c0.n4327\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__12914\,
            I => \c0.n4327\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__12909\,
            I => \c0.n4434_cascade_\
        );

    \I__1212\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12903\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__12903\,
            I => \c0.n8766\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__12900\,
            I => \c0.n9482_cascade_\
        );

    \I__1209\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12894\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12894\,
            I => \N__12891\
        );

    \I__1207\ : Span4Mux_v
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__12888\,
            I => \c0.n9207\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \c0.n9548_cascade_\
        );

    \I__1204\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12879\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__12879\,
            I => \N__12876\
        );

    \I__1202\ : Span4Mux_s3_v
    port map (
            O => \N__12876\,
            I => \N__12873\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__12873\,
            I => \N__12870\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__12870\,
            I => \c0.n9177\
        );

    \I__1199\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12863\
        );

    \I__1198\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12858\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__12863\,
            I => \N__12855\
        );

    \I__1196\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12850\
        );

    \I__1195\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12850\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__12858\,
            I => \N__12847\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__12855\,
            I => \c0.data_in_field_10\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__12850\,
            I => \c0.data_in_field_10\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__12847\,
            I => \c0.data_in_field_10\
        );

    \I__1190\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12834\
        );

    \I__1189\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12834\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__12834\,
            I => data_in_12_7
        );

    \I__1187\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12827\
        );

    \I__1186\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12824\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__12827\,
            I => data_in_13_4
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__12824\,
            I => data_in_13_4
        );

    \I__1183\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12813\
        );

    \I__1182\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12813\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__12813\,
            I => data_in_14_4
        );

    \I__1180\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12804\
        );

    \I__1179\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12804\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__12804\,
            I => data_in_10_0
        );

    \I__1177\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__12798\,
            I => \N__12794\
        );

    \I__1175\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12791\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__12794\,
            I => data_in_11_0
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__12791\,
            I => data_in_11_0
        );

    \I__1172\ : InMux
    port map (
            O => \N__12786\,
            I => \c0.tx2.n8109\
        );

    \I__1171\ : InMux
    port map (
            O => \N__12783\,
            I => \c0.tx2.n8110\
        );

    \I__1170\ : InMux
    port map (
            O => \N__12780\,
            I => \c0.tx2.n8111\
        );

    \I__1169\ : InMux
    port map (
            O => \N__12777\,
            I => \bfn_1_32_0_\
        );

    \I__1168\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12768\
        );

    \I__1167\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12768\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__12768\,
            I => data_in_7_7
        );

    \I__1165\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12759\
        );

    \I__1164\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12759\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__12759\,
            I => data_in_10_7
        );

    \I__1162\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12750\
        );

    \I__1161\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12750\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__12750\,
            I => data_in_11_7
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__12747\,
            I => \c0.n9524_cascade_\
        );

    \I__1158\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__12741\,
            I => \c0.n9183\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__12738\,
            I => \c0.n9186_cascade_\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__12735\,
            I => \c0.n9518_cascade_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__12729\,
            I => \N__12726\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__12726\,
            I => \c0.n22_adj_1680\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__12723\,
            I => \c0.n9521_cascade_\
        );

    \I__1150\ : InMux
    port map (
            O => \N__12720\,
            I => \N__12717\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__12717\,
            I => \c0.tx2.r_Clock_Count_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__12714\,
            I => \bfn_1_31_0_\
        );

    \I__1147\ : InMux
    port map (
            O => \N__12711\,
            I => \c0.tx2.n8105\
        );

    \I__1146\ : InMux
    port map (
            O => \N__12708\,
            I => \c0.tx2.n8106\
        );

    \I__1145\ : InMux
    port map (
            O => \N__12705\,
            I => \c0.tx2.n8107\
        );

    \I__1144\ : InMux
    port map (
            O => \N__12702\,
            I => \c0.tx2.n8108\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__12699\,
            I => \c0.n9464_cascade_\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__12696\,
            I => \c0.n9470_cascade_\
        );

    \I__1141\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12690\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__12690\,
            I => \c0.n9216\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__12687\,
            I => \c0.n9213_cascade_\
        );

    \I__1138\ : InMux
    port map (
            O => \N__12684\,
            I => \N__12681\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__12681\,
            I => \N__12678\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__12678\,
            I => \c0.n9210\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__12675\,
            I => \c0.n9458_cascade_\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__12672\,
            I => \c0.n9461_cascade_\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__12669\,
            I => \c0.n9530_cascade_\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__12666\,
            I => \c0.n54_cascade_\
        );

    \I__1131\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12660\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__12660\,
            I => \c0.n49\
        );

    \I__1129\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12654\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__12654\,
            I => \c0.n9001\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__12651\,
            I => \c0.n9001_cascade_\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__12648\,
            I => \c0.n10_adj_1637_cascade_\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__12645\,
            I => \N__12642\
        );

    \I__1124\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12639\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__12639\,
            I => \c0.data_in_frame_19_3\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__12636\,
            I => \c0.n9686_cascade_\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__12633\,
            I => \c0.n9689_cascade_\
        );

    \I__1120\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12627\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__12624\,
            I => \c0.n10_adj_1646\
        );

    \I__1117\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12617\
        );

    \I__1116\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12614\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__12617\,
            I => \N__12611\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__12614\,
            I => \c0.n8779\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__12611\,
            I => \c0.n8779\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__12606\,
            I => \c0.n9674_cascade_\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__12603\,
            I => \c0.n9677_cascade_\
        );

    \I__1110\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12597\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__12597\,
            I => \N__12594\
        );

    \I__1108\ : Odrv12
    port map (
            O => \N__12594\,
            I => \c0.n4431\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__12591\,
            I => \c0.n8849_cascade_\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__12588\,
            I => \c0.n20_adj_1622_cascade_\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__12585\,
            I => \N__12582\
        );

    \I__1104\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12579\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__12579\,
            I => \c0.data_in_frame_19_5\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__12576\,
            I => \c0.n4431_cascade_\
        );

    \I__1101\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12570\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__12570\,
            I => n1902
        );

    \I__1099\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12564\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__12564\,
            I => \N__12559\
        );

    \I__1097\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12556\
        );

    \I__1096\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12553\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__12559\,
            I => \N__12550\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__12556\,
            I => data_in_6_4
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__12553\,
            I => data_in_6_4
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__12550\,
            I => data_in_6_4
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__12543\,
            I => \c0.n24_cascade_\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__12540\,
            I => \c0.n4_adj_1594_cascade_\
        );

    \I__1089\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12528\
        );

    \I__1088\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12528\
        );

    \I__1087\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12528\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__12528\,
            I => data_in_5_1
        );

    \I__1085\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12520\
        );

    \I__1084\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12515\
        );

    \I__1083\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12515\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__12520\,
            I => data_in_6_1
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__12515\,
            I => data_in_6_1
        );

    \I__1080\ : InMux
    port map (
            O => \N__12510\,
            I => \N__12504\
        );

    \I__1079\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12504\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__12504\,
            I => data_in_7_1
        );

    \I__1077\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12498\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__12498\,
            I => \N__12494\
        );

    \I__1075\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12491\
        );

    \I__1074\ : Odrv12
    port map (
            O => \N__12494\,
            I => data_in_9_1
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__12491\,
            I => data_in_9_1
        );

    \I__1072\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12480\
        );

    \I__1071\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12480\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__12480\,
            I => data_in_8_1
        );

    \I__1069\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12471\
        );

    \I__1068\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12471\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__12471\,
            I => data_in_13_1
        );

    \I__1066\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12462\
        );

    \I__1065\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12462\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__12462\,
            I => data_in_12_1
        );

    \I__1063\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12453\
        );

    \I__1062\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12453\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__12453\,
            I => data_in_7_4
        );

    \I__1060\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12444\
        );

    \I__1059\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12444\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__12444\,
            I => data_in_8_4
        );

    \I__1057\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12435\
        );

    \I__1056\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12435\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__12435\,
            I => data_in_9_4
        );

    \I__1054\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12426\
        );

    \I__1053\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12426\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__12426\,
            I => data_in_10_4
        );

    \I__1051\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12417\
        );

    \I__1050\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12417\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__12417\,
            I => data_in_11_4
        );

    \I__1048\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12408\
        );

    \I__1047\ : InMux
    port map (
            O => \N__12413\,
            I => \N__12408\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__12408\,
            I => data_in_12_4
        );

    \I__1045\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12399\
        );

    \I__1044\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12399\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__12399\,
            I => data_in_10_1
        );

    \I__1042\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12390\
        );

    \I__1041\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12390\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__12390\,
            I => data_in_11_1
        );

    \I__1039\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12381\
        );

    \I__1038\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12381\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__12381\,
            I => data_in_14_1
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__12378\,
            I => \N__12375\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__12375\,
            I => \N__12372\
        );

    \I__1034\ : IoSpan4Mux
    port map (
            O => \N__12372\,
            I => \N__12369\
        );

    \I__1033\ : IoSpan4Mux
    port map (
            O => \N__12369\,
            I => \N__12366\
        );

    \I__1032\ : IoSpan4Mux
    port map (
            O => \N__12366\,
            I => \N__12363\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__12363\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_6_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_27_0_\
        );

    \IN_MUX_bfv_6_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n8162,
            carryinitout => \bfn_6_28_0_\
        );

    \IN_MUX_bfv_6_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n8170,
            carryinitout => \bfn_6_29_0_\
        );

    \IN_MUX_bfv_6_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n8178,
            carryinitout => \bfn_6_30_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_1_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx2.n8112\,
            carryinitout => \bfn_1_32_0_\
        );

    \IN_MUX_bfv_15_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_30_0_\
        );

    \IN_MUX_bfv_15_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n8097\,
            carryinitout => \bfn_15_31_0_\
        );

    \IN_MUX_bfv_11_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_31_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_16_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n8127\,
            carryinitout => \bfn_16_26_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_11_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_27_0_\
        );

    \IN_MUX_bfv_11_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n8137,
            carryinitout => \bfn_11_28_0_\
        );

    \IN_MUX_bfv_11_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n8145,
            carryinitout => \bfn_11_29_0_\
        );

    \IN_MUX_bfv_11_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n8153,
            carryinitout => \bfn_11_30_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12378\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.data_in_0___i74_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12405\,
            in1 => \N__29627\,
            in2 => \_gnd_net_\,
            in3 => \N__12497\,
            lcout => data_in_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i82_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12396\,
            in1 => \_gnd_net_\,
            in2 => \N__29843\,
            in3 => \N__12404\,
            lcout => data_in_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i90_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29631\,
            in1 => \N__12468\,
            in2 => \_gnd_net_\,
            in3 => \N__12395\,
            lcout => data_in_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i106_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12387\,
            in1 => \N__29626\,
            in2 => \_gnd_net_\,
            in3 => \N__12476\,
            lcout => data_in_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i114_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29625\,
            in1 => \N__16068\,
            in2 => \_gnd_net_\,
            in3 => \N__12386\,
            lcout => data_in_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i98_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29632\,
            in1 => \N__12477\,
            in2 => \_gnd_net_\,
            in3 => \N__12467\,
            lcout => data_in_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i53_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12459\,
            in1 => \N__29779\,
            in2 => \_gnd_net_\,
            in3 => \N__12562\,
            lcout => data_in_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i61_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12450\,
            in1 => \N__29776\,
            in2 => \_gnd_net_\,
            in3 => \N__12458\,
            lcout => data_in_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i69_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12441\,
            in1 => \N__29780\,
            in2 => \_gnd_net_\,
            in3 => \N__12449\,
            lcout => data_in_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i77_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12432\,
            in1 => \N__29777\,
            in2 => \_gnd_net_\,
            in3 => \N__12440\,
            lcout => data_in_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i85_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12423\,
            in1 => \N__29781\,
            in2 => \_gnd_net_\,
            in3 => \N__12431\,
            lcout => data_in_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i93_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12414\,
            in1 => \N__29778\,
            in2 => \_gnd_net_\,
            in3 => \N__12422\,
            lcout => data_in_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i101_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29775\,
            in1 => \N__12831\,
            in2 => \_gnd_net_\,
            in3 => \N__12413\,
            lcout => data_in_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i45_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29929\,
            in1 => \N__12563\,
            in2 => \_gnd_net_\,
            in3 => \N__16036\,
            lcout => data_in_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_41_i1_3_lut_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12535\,
            in1 => \N__19601\,
            in2 => \_gnd_net_\,
            in3 => \N__23419\,
            lcout => n1902,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i42_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12525\,
            in1 => \N__12536\,
            in2 => \_gnd_net_\,
            in3 => \N__29931\,
            lcout => data_in_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i34_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12537\,
            in1 => \_gnd_net_\,
            in2 => \N__30018\,
            in3 => \N__13628\,
            lcout => data_in_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13627\,
            in1 => \N__29930\,
            in2 => \_gnd_net_\,
            in3 => \N__13557\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i50_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__12524\,
            in1 => \_gnd_net_\,
            in2 => \N__30019\,
            in3 => \N__12510\,
            lcout => data_in_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_49_i1_3_lut_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23418\,
            in1 => \N__12523\,
            in2 => \_gnd_net_\,
            in3 => \N__19856\,
            lcout => n1894,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i58_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12485\,
            in2 => \N__30020\,
            in3 => \N__12509\,
            lcout => data_in_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i66_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12486\,
            in1 => \N__12501\,
            in2 => \_gnd_net_\,
            in3 => \N__29932\,
            lcout => data_in_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_677_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24754\,
            in1 => \N__18601\,
            in2 => \N__28300\,
            in3 => \N__28240\,
            lcout => \c0.n4431\,
            ltout => \c0.n4431_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_511_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22358\,
            in1 => \N__16712\,
            in2 => \N__12576\,
            in3 => \N__22476\,
            lcout => \c0.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_667_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24755\,
            in1 => \N__16847\,
            in2 => \_gnd_net_\,
            in3 => \N__18602\,
            lcout => \c0.n8878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i42_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__24776\,
            in1 => \N__12573\,
            in2 => \N__19152\,
            in3 => \_gnd_net_\,
            lcout => data_in_field_41,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_52_i1_3_lut_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12567\,
            in1 => \N__24336\,
            in2 => \_gnd_net_\,
            in3 => \N__23420\,
            lcout => n1891,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_658_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17305\,
            in1 => \N__16496\,
            in2 => \_gnd_net_\,
            in3 => \N__18716\,
            lcout => \c0.n24\,
            ltout => \c0.n24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_706_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12921\,
            in1 => \N__14912\,
            in2 => \N__12543\,
            in3 => \N__15085\,
            lcout => \c0.n8858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22674\,
            in1 => \N__18759\,
            in2 => \N__22984\,
            in3 => \N__22200\,
            lcout => OPEN,
            ltout => \c0.n4_adj_1594_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_519_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__23027\,
            in1 => \N__22976\,
            in2 => \N__12540\,
            in3 => \N__12621\,
            lcout => \c0.n22_adj_1595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i44_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22977\,
            in1 => \N__19154\,
            in2 => \_gnd_net_\,
            in3 => \N__13386\,
            lcout => data_in_field_43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_741_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22199\,
            in1 => \N__22673\,
            in2 => \_gnd_net_\,
            in3 => \N__22972\,
            lcout => \c0.n8766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9512_bdd_4_lut_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__33151\,
            in1 => \N__12862\,
            in2 => \N__16779\,
            in3 => \N__14946\,
            lcout => \c0.n9192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i14_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__23516\,
            in1 => \N__22207\,
            in2 => \N__13500\,
            in3 => \N__19147\,
            lcout => \c0.data_in_field_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_636_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15117\,
            in1 => \N__12861\,
            in2 => \N__12936\,
            in3 => \N__22614\,
            lcout => \c0.n10_adj_1646\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i11_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__19153\,
            in1 => \N__14748\,
            in2 => \N__23558\,
            in3 => \N__12867\,
            lcout => \c0.data_in_field_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7970_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__19770\,
            in1 => \N__32985\,
            in2 => \N__12585\,
            in3 => \N__32014\,
            lcout => OPEN,
            ltout => \c0.n9674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9674_bdd_4_lut_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32986\,
            in1 => \N__32606\,
            in2 => \N__12606\,
            in3 => \N__19932\,
            lcout => OPEN,
            ltout => \c0.n9677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__13059\,
            in1 => \N__31377\,
            in2 => \N__12603\,
            in3 => \N__31204\,
            lcout => \c0.n22_adj_1678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_666_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12957\,
            in1 => \N__14413\,
            in2 => \_gnd_net_\,
            in3 => \N__12600\,
            lcout => \c0.n8849\,
            ltout => \c0.n8849_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_575_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27371\,
            in1 => \N__22068\,
            in2 => \N__12591\,
            in3 => \N__19686\,
            lcout => OPEN,
            ltout => \c0.n20_adj_1622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i158_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13215\,
            in2 => \N__12588\,
            in3 => \N__21105\,
            lcout => \c0.data_in_frame_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35316\,
            ce => \N__29066\,
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17472\,
            in2 => \_gnd_net_\,
            in3 => \N__12620\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1637_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i156_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26757\,
            in1 => \N__14160\,
            in2 => \N__12648\,
            in3 => \N__20630\,
            lcout => \c0.data_in_frame_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35323\,
            ce => \N__29004\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7984_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33208\,
            in1 => \N__15604\,
            in2 => \N__12645\,
            in3 => \N__32040\,
            lcout => OPEN,
            ltout => \c0.n9686_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9686_bdd_4_lut_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__17398\,
            in1 => \N__33209\,
            in2 => \N__12636\,
            in3 => \N__23782\,
            lcout => OPEN,
            ltout => \c0.n9689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17847\,
            in1 => \N__31376\,
            in2 => \N__12633\,
            in3 => \N__31231\,
            lcout => \c0.n22_adj_1680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12630\,
            in1 => \N__14417\,
            in2 => \_gnd_net_\,
            in3 => \N__13979\,
            lcout => \c0.n8779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16973\,
            in1 => \_gnd_net_\,
            in2 => \N__30036\,
            in3 => \N__13903\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13838\,
            in1 => \N__30021\,
            in2 => \_gnd_net_\,
            in3 => \N__16972\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_697_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22532\,
            in1 => \N__13008\,
            in2 => \_gnd_net_\,
            in3 => \N__22018\,
            lcout => \c0.n6_adj_1654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9476_bdd_4_lut_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__33173\,
            in1 => \N__24780\,
            in2 => \N__20310\,
            in3 => \N__14913\,
            lcout => \c0.n9210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13733\,
            in1 => \_gnd_net_\,
            in2 => \N__14830\,
            in3 => \N__30022\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30024\,
            in1 => \N__14820\,
            in2 => \_gnd_net_\,
            in3 => \N__13837\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i48_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13095\,
            in1 => \N__30023\,
            in2 => \_gnd_net_\,
            in3 => \N__13195\,
            lcout => data_in_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13101\,
            in1 => \N__17274\,
            in2 => \N__13704\,
            in3 => \N__13017\,
            lcout => OPEN,
            ltout => \c0.n54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i162_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12999\,
            in1 => \N__22179\,
            in2 => \N__12666\,
            in3 => \N__12663\,
            lcout => \c0.data_in_frame_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35337\,
            ce => \N__29067\,
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27186\,
            in1 => \N__12657\,
            in2 => \N__17637\,
            in3 => \N__18780\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_714_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24561\,
            in1 => \N__18470\,
            in2 => \N__24503\,
            in3 => \N__17468\,
            lcout => \c0.n9001\,
            ltout => \c0.n9001_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_546_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25083\,
            in1 => \N__17832\,
            in2 => \N__12651\,
            in3 => \N__15519\,
            lcout => \c0.n28_adj_1612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7795_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__33190\,
            in1 => \N__32041\,
            in2 => \N__19818\,
            in3 => \N__21622\,
            lcout => OPEN,
            ltout => \c0.n9464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9464_bdd_4_lut_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__27791\,
            in1 => \N__14181\,
            in2 => \N__12699\,
            in3 => \N__33191\,
            lcout => \c0.n9216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7800_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33192\,
            in1 => \N__15869\,
            in2 => \N__17955\,
            in3 => \N__32042\,
            lcout => OPEN,
            ltout => \c0.n9470_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9470_bdd_4_lut_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__24490\,
            in1 => \N__20751\,
            in2 => \N__12696\,
            in3 => \N__33193\,
            lcout => OPEN,
            ltout => \c0.n9213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_7810_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__31617\,
            in1 => \N__12693\,
            in2 => \N__12687\,
            in3 => \N__31229\,
            lcout => OPEN,
            ltout => \c0.n9458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9458_bdd_4_lut_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__12897\,
            in1 => \N__12684\,
            in2 => \N__12675\,
            in3 => \N__31618\,
            lcout => OPEN,
            ltout => \c0.n9461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i1_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31619\,
            in1 => \N__14019\,
            in2 => \N__12672\,
            in3 => \N__32377\,
            lcout => \c0.tx2.r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35344\,
            ce => \N__32273\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7850_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33199\,
            in1 => \N__14247\,
            in2 => \N__21894\,
            in3 => \N__32057\,
            lcout => OPEN,
            ltout => \c0.n9530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9530_bdd_4_lut_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__17130\,
            in1 => \N__17103\,
            in2 => \N__12669\,
            in3 => \N__33200\,
            lcout => \c0.n9183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7845_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33201\,
            in1 => \N__15669\,
            in2 => \N__26691\,
            in3 => \N__32058\,
            lcout => OPEN,
            ltout => \c0.n9524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9524_bdd_4_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__23852\,
            in1 => \N__33202\,
            in2 => \N__12747\,
            in3 => \N__17732\,
            lcout => OPEN,
            ltout => \c0.n9186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_7865_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__12744\,
            in1 => \N__31630\,
            in2 => \N__12738\,
            in3 => \N__31230\,
            lcout => OPEN,
            ltout => \c0.n9518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9518_bdd_4_lut_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31631\,
            in1 => \N__12882\,
            in2 => \N__12735\,
            in3 => \N__12975\,
            lcout => OPEN,
            ltout => \c0.n9521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i3_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__12732\,
            in1 => \N__31632\,
            in2 => \N__12723\,
            in3 => \N__32388\,
            lcout => \c0.tx2.r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35352\,
            ce => \N__32264\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count__i0_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12720\,
            in2 => \_gnd_net_\,
            in3 => \N__12714\,
            lcout => \c0.tx2.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_1_31_0_\,
            carryout => \c0.tx2.n8105\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i1_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13142\,
            in2 => \_gnd_net_\,
            in3 => \N__12711\,
            lcout => \c0.tx2.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.tx2.n8105\,
            carryout => \c0.tx2.n8106\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i2_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13167\,
            in2 => \_gnd_net_\,
            in3 => \N__12708\,
            lcout => \c0.tx2.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.tx2.n8106\,
            carryout => \c0.tx2.n8107\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i3_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13128\,
            in2 => \_gnd_net_\,
            in3 => \N__12705\,
            lcout => \c0.tx2.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.tx2.n8107\,
            carryout => \c0.tx2.n8108\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i4_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13116\,
            in2 => \_gnd_net_\,
            in3 => \N__12702\,
            lcout => \c0.tx2.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.tx2.n8108\,
            carryout => \c0.tx2.n8109\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i5_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13356\,
            in2 => \_gnd_net_\,
            in3 => \N__12786\,
            lcout => \c0.tx2.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.tx2.n8109\,
            carryout => \c0.tx2.n8110\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i6_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13155\,
            in2 => \_gnd_net_\,
            in3 => \N__12783\,
            lcout => \c0.tx2.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.tx2.n8110\,
            carryout => \c0.tx2.n8111\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i7_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13341\,
            in2 => \_gnd_net_\,
            in3 => \N__12780\,
            lcout => \c0.tx2.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \c0.tx2.n8111\,
            carryout => \c0.tx2.n8112\,
            clk => \N__35359\,
            ce => \N__26876\,
            sr => \N__13307\
        );

    \c0.tx2.r_Clock_Count__i8_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13287\,
            in2 => \_gnd_net_\,
            in3 => \N__12777\,
            lcout => \c0.tx2.r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35367\,
            ce => \N__26880\,
            sr => \N__13311\
        );

    \c0.data_in_0___i56_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12774\,
            in1 => \_gnd_net_\,
            in2 => \N__29844\,
            in3 => \N__13087\,
            lcout => data_in_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i64_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29642\,
            in1 => \N__13398\,
            in2 => \_gnd_net_\,
            in3 => \N__12773\,
            lcout => data_in_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i80_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12765\,
            in1 => \N__29634\,
            in2 => \_gnd_net_\,
            in3 => \N__13409\,
            lcout => data_in_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i88_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12756\,
            in1 => \_gnd_net_\,
            in2 => \N__29845\,
            in3 => \N__12764\,
            lcout => data_in_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i96_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12840\,
            in1 => \N__29635\,
            in2 => \_gnd_net_\,
            in3 => \N__12755\,
            lcout => data_in_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i104_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29633\,
            in1 => \N__12839\,
            in2 => \_gnd_net_\,
            in3 => \N__14499\,
            lcout => data_in_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i109_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29570\,
            in1 => \N__12830\,
            in2 => \_gnd_net_\,
            in3 => \N__12819\,
            lcout => data_in_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i73_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12810\,
            in1 => \N__29713\,
            in2 => \_gnd_net_\,
            in3 => \N__13532\,
            lcout => data_in_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i117_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29571\,
            in1 => \N__16335\,
            in2 => \_gnd_net_\,
            in3 => \N__12818\,
            lcout => data_in_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i81_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29712\,
            in1 => \N__12801\,
            in2 => \_gnd_net_\,
            in3 => \N__12809\,
            lcout => data_in_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29492\,
            in1 => \N__13685\,
            in2 => \_gnd_net_\,
            in3 => \N__14747\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_679_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18449\,
            in1 => \N__13752\,
            in2 => \N__13496\,
            in3 => \N__16642\,
            lcout => \c0.n14_adj_1669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29485\,
            in1 => \_gnd_net_\,
            in2 => \N__13760\,
            in3 => \N__16646\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16750\,
            in1 => \N__29486\,
            in2 => \_gnd_net_\,
            in3 => \N__13753\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i89_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__13470\,
            in1 => \_gnd_net_\,
            in2 => \N__29700\,
            in3 => \N__12797\,
            lcout => data_in_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13491\,
            in1 => \N__29487\,
            in2 => \_gnd_net_\,
            in3 => \N__16262\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29488\,
            in1 => \N__13561\,
            in2 => \_gnd_net_\,
            in3 => \N__16749\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_683_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14831\,
            in1 => \N__14856\,
            in2 => \N__13565\,
            in3 => \N__13684\,
            lcout => \c0.n26_adj_1673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_46_i1_3_lut_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22305\,
            in1 => \N__16224\,
            in2 => \_gnd_net_\,
            in3 => \N__23325\,
            lcout => n1897,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7870_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__32038\,
            in1 => \N__33034\,
            in2 => \N__28305\,
            in3 => \N__13792\,
            lcout => OPEN,
            ltout => \c0.n9548_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9548_bdd_4_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__12952\,
            in1 => \N__33064\,
            in2 => \N__12885\,
            in3 => \N__15086\,
            lcout => \c0.n9177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9578_bdd_4_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__13934\,
            in1 => \N__33033\,
            in2 => \N__13581\,
            in3 => \N__18813\,
            lcout => \c0.n9162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_712_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13790\,
            in1 => \N__13932\,
            in2 => \N__18857\,
            in3 => \N__17068\,
            lcout => \c0.n4327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_736_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12866\,
            in1 => \N__12951\,
            in2 => \_gnd_net_\,
            in3 => \N__16839\,
            lcout => \c0.n4224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_731_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13933\,
            lcout => OPEN,
            ltout => \c0.n8801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13572\,
            in1 => \N__15137\,
            in2 => \N__12960\,
            in3 => \N__16816\,
            lcout => \c0.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i12_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__12953\,
            in1 => \N__23429\,
            in2 => \N__14691\,
            in3 => \N__19146\,
            lcout => \c0.data_in_field_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35311\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_631_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28229\,
            in2 => \_gnd_net_\,
            in3 => \N__15291\,
            lcout => \c0.n4276\,
            ltout => \c0.n4276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_598_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27975\,
            in1 => \N__17312\,
            in2 => \N__12927\,
            in3 => \N__13668\,
            lcout => OPEN,
            ltout => \c0.n12_adj_1633_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_603_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21315\,
            in1 => \N__16728\,
            in2 => \N__12924\,
            in3 => \N__12920\,
            lcout => \c0.n4434\,
            ltout => \c0.n4434_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_593_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18773\,
            in1 => \N__15845\,
            in2 => \N__12909\,
            in3 => \N__12906\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7815_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__28230\,
            in1 => \N__32039\,
            in2 => \N__33174\,
            in3 => \N__17313\,
            lcout => OPEN,
            ltout => \c0.n9482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9482_bdd_4_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__15293\,
            in1 => \N__16626\,
            in2 => \N__12900\,
            in3 => \N__33115\,
            lcout => \c0.n9207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i50_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22368\,
            in1 => \N__12990\,
            in2 => \_gnd_net_\,
            in3 => \N__19108\,
            lcout => data_in_field_49,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7860_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__17503\,
            in1 => \N__32891\,
            in2 => \N__17549\,
            in3 => \N__31992\,
            lcout => OPEN,
            ltout => \c0.n9542_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9542_bdd_4_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__13605\,
            in1 => \N__32892\,
            in2 => \N__12978\,
            in3 => \N__22983\,
            lcout => \c0.n9180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i36_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__23484\,
            in1 => \N__15192\,
            in2 => \N__19158\,
            in3 => \N__13606\,
            lcout => \c0.data_in_field_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_711_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21409\,
            in1 => \N__17502\,
            in2 => \_gnd_net_\,
            in3 => \N__15827\,
            lcout => \c0.n8855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_579_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23781\,
            in2 => \_gnd_net_\,
            in3 => \N__26685\,
            lcout => \c0.n4577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29614\,
            in1 => \N__16883\,
            in2 => \_gnd_net_\,
            in3 => \N__15261\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_687_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17057\,
            in1 => \N__13604\,
            in2 => \N__21322\,
            in3 => \N__14898\,
            lcout => \c0.n4114\,
            ltout => \c0.n4114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_664_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15826\,
            in2 => \N__12963\,
            in3 => \N__21367\,
            lcout => \c0.n8864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25677\,
            in1 => \N__13026\,
            in2 => \N__15351\,
            in3 => \N__17511\,
            lcout => OPEN,
            ltout => \c0.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i168_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32457\,
            in1 => \N__15681\,
            in2 => \N__13032\,
            in3 => \N__14136\,
            lcout => \c0.data_in_frame_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35331\,
            ce => \N__29003\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_628_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17228\,
            in1 => \N__13797\,
            in2 => \_gnd_net_\,
            in3 => \N__16379\,
            lcout => \c0.n4324\,
            ltout => \c0.n4324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31733\,
            in1 => \N__27666\,
            in2 => \N__13029\,
            in3 => \N__17762\,
            lcout => \c0.n8951\,
            ltout => \c0.n8951_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26787\,
            in1 => \N__28206\,
            in2 => \N__13020\,
            in3 => \N__17204\,
            lcout => \c0.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_735_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31734\,
            in1 => \N__27667\,
            in2 => \_gnd_net_\,
            in3 => \N__17763\,
            lcout => \c0.n4479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_662_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14942\,
            in1 => \N__13952\,
            in2 => \N__17265\,
            in3 => \N__15087\,
            lcout => \c0.n8930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_680_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16971\,
            in1 => \N__13813\,
            in2 => \N__13904\,
            in3 => \N__13836\,
            lcout => \c0.n14_adj_1670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_703_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17099\,
            in1 => \_gnd_net_\,
            in2 => \N__17603\,
            in3 => \N__15595\,
            lcout => \c0.n4406\,
            ltout => \c0.n4406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17406\,
            in1 => \N__27792\,
            in2 => \N__13002\,
            in3 => \N__14112\,
            lcout => \c0.n43_adj_1610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i108_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19565\,
            in1 => \N__17728\,
            in2 => \_gnd_net_\,
            in3 => \N__29032\,
            lcout => data_in_field_107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i90_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21669\,
            in1 => \_gnd_net_\,
            in2 => \N__29069\,
            in3 => \N__17944\,
            lcout => data_in_field_89,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_580_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15624\,
            lcout => \c0.n8921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i72_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__15625\,
            in1 => \_gnd_net_\,
            in2 => \N__29068\,
            in3 => \N__21085\,
            lcout => data_in_field_71,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i102_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24158\,
            in1 => \N__19303\,
            in2 => \_gnd_net_\,
            in3 => \N__29031\,
            lcout => data_in_field_101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i166_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15531\,
            in1 => \N__15350\,
            in2 => \N__22101\,
            in3 => \N__13038\,
            lcout => \c0.data_in_frame_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35345\,
            ce => \N__29026\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_715_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20631\,
            in1 => \N__26081\,
            in2 => \_gnd_net_\,
            in3 => \N__14066\,
            lcout => \c0.n4215\,
            ltout => \c0.n4215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_518_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13068\,
            in1 => \N__17358\,
            in2 => \N__13044\,
            in3 => \N__16680\,
            lcout => OPEN,
            ltout => \c0.n18_adj_1593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_520_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14145\,
            in1 => \N__17966\,
            in2 => \N__13041\,
            in3 => \N__22375\,
            lcout => \c0.n20_adj_1596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_611_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26409\,
            in1 => \N__32172\,
            in2 => \_gnd_net_\,
            in3 => \N__26329\,
            lcout => OPEN,
            ltout => \c0.n4568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24605\,
            in1 => \N__15393\,
            in2 => \N__13104\,
            in3 => \N__24861\,
            lcout => \c0.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_47_i1_3_lut_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19506\,
            in1 => \N__13202\,
            in2 => \_gnd_net_\,
            in3 => \N__23266\,
            lcout => n1896,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state__i0_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23676\,
            in2 => \N__23326\,
            in3 => \N__23616\,
            lcout => \FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35353\,
            ce => \N__20808\,
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_55_i1_3_lut_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23262\,
            in1 => \N__13094\,
            in2 => \_gnd_net_\,
            in3 => \N__19714\,
            lcout => n1888,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4613_3_lut_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21507\,
            in1 => \N__16050\,
            in2 => \_gnd_net_\,
            in3 => \N__23267\,
            lcout => n6164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_527_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24488\,
            in2 => \_gnd_net_\,
            in3 => \N__28397\,
            lcout => \c0.n9004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_540_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21950\,
            in2 => \_gnd_net_\,
            in3 => \N__21893\,
            lcout => \c0.n8816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_642_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17589\,
            in2 => \_gnd_net_\,
            in3 => \N__15606\,
            lcout => \c0.n8807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_574_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15605\,
            in1 => \N__19635\,
            in2 => \N__15436\,
            in3 => \N__27729\,
            lcout => \c0.n4282\,
            ltout => \c0.n4282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13062\,
            in3 => \N__24560\,
            lcout => \c0.n9007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_629_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15871\,
            in2 => \_gnd_net_\,
            in3 => \N__14246\,
            lcout => OPEN,
            ltout => \c0.n4476_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_576_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13236\,
            in1 => \N__13224\,
            in2 => \N__13218\,
            in3 => \N__21951\,
            lcout => \c0.n19_adj_1623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i40_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13720\,
            in1 => \N__29396\,
            in2 => \_gnd_net_\,
            in3 => \N__13203\,
            lcout => data_in_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i82_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19857\,
            in1 => \N__15872\,
            in2 => \_gnd_net_\,
            in3 => \N__29070\,
            lcout => data_in_field_81,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15782\,
            lcout => tx2_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14304\,
            in2 => \_gnd_net_\,
            in3 => \N__13283\,
            lcout => \c0.tx2.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i2_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__13285\,
            in1 => \N__13329\,
            in2 => \N__14317\,
            in3 => \N__13263\,
            lcout => \r_SM_Main_2_adj_1738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_4_lut_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__13166\,
            in1 => \N__13154\,
            in2 => \N__13143\,
            in3 => \N__13127\,
            lcout => OPEN,
            ltout => \c0.tx2.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5854_4_lut_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__13115\,
            in1 => \N__13355\,
            in2 => \N__13344\,
            in3 => \N__13340\,
            lcout => \c0.tx2.n7399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1_2_lut_2_lut_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26917\,
            in2 => \_gnd_net_\,
            in3 => \N__15940\,
            lcout => \c0.tx2.n4081\,
            ltout => \c0.tx2.n4081_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_4_lut_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13284\,
            in1 => \N__14318\,
            in2 => \N__13323\,
            in3 => \N__13261\,
            lcout => OPEN,
            ltout => \c0.tx2.n8196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i7758_4_lut_4_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__13262\,
            in1 => \N__13320\,
            in2 => \N__13314\,
            in3 => \N__26918\,
            lcout => \c0.tx2.n5146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i7404_4_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__26919\,
            in1 => \N__15941\,
            in2 => \N__14319\,
            in3 => \N__14264\,
            lcout => n9075,
            ltout => \n9075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i7412_3_lut_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__15942\,
            in1 => \_gnd_net_\,
            in2 => \N__13290\,
            in3 => \N__13245\,
            lcout => n5346,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i5868_2_lut_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13286\,
            in2 => \_gnd_net_\,
            in3 => \N__13260\,
            lcout => \r_SM_Main_2_N_1480_1_adj_1744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16110\,
            in1 => \N__14332\,
            in2 => \_gnd_net_\,
            in3 => \N__16179\,
            lcout => \c0.tx2.n7236\,
            ltout => \c0.tx2.n7236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i1673_4_lut_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__20473\,
            in1 => \N__15943\,
            in2 => \N__13239\,
            in3 => \N__14265\,
            lcout => OPEN,
            ltout => \n3220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i0_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110100"
        )
    port map (
            in0 => \N__14267\,
            in1 => \N__14315\,
            in2 => \N__13413\,
            in3 => \N__26920\,
            lcout => \r_SM_Main_0_adj_1740\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_i1_LC_2_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__14266\,
            in1 => \N__14314\,
            in2 => \N__15950\,
            in3 => \N__26921\,
            lcout => \r_SM_Main_1_adj_1739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i72_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29650\,
            in1 => \N__13410\,
            in2 => \_gnd_net_\,
            in3 => \N__13397\,
            lcout => data_in_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_43_i1_3_lut_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19566\,
            in1 => \N__15215\,
            in2 => \_gnd_net_\,
            in3 => \N__23541\,
            lcout => n1900,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i71_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29861\,
            in1 => \N__14472\,
            in2 => \_gnd_net_\,
            in3 => \N__16580\,
            lcout => data_in_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i111_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14613\,
            in1 => \N__29862\,
            in2 => \_gnd_net_\,
            in3 => \N__14441\,
            lcout => data_in_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i52_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29859\,
            in1 => \N__13374\,
            in2 => \_gnd_net_\,
            in3 => \N__14705\,
            lcout => data_in_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_51_i1_3_lut_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14704\,
            in1 => \N__19438\,
            in2 => \_gnd_net_\,
            in3 => \N__23540\,
            lcout => n1892,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i60_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__13365\,
            in1 => \_gnd_net_\,
            in2 => \N__29986\,
            in3 => \N__13373\,
            lcout => data_in_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i68_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29759\,
            in1 => \N__18129\,
            in2 => \_gnd_net_\,
            in3 => \N__13364\,
            lcout => data_in_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i65_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29860\,
            in1 => \N__13533\,
            in2 => \_gnd_net_\,
            in3 => \N__13520\,
            lcout => data_in_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i49_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13509\,
            in1 => \N__29493\,
            in2 => \_gnd_net_\,
            in3 => \N__20545\,
            lcout => data_in_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i57_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__13521\,
            in1 => \_gnd_net_\,
            in2 => \N__29701\,
            in3 => \N__13508\,
            lcout => data_in_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14555\,
            in1 => \N__13492\,
            in2 => \_gnd_net_\,
            in3 => \N__29497\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i97_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29358\,
            in1 => \N__14796\,
            in2 => \_gnd_net_\,
            in3 => \N__13466\,
            lcout => data_in_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_704_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14993\,
            in1 => \N__18515\,
            in2 => \N__14740\,
            in3 => \N__18552\,
            lcout => \c0.n25_adj_1675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7366_4_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13455\,
            in1 => \N__14760\,
            in2 => \N__13443\,
            in3 => \N__14754\,
            lcout => OPEN,
            ltout => \c0.n9033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_723_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__13434\,
            in1 => \N__13422\,
            in2 => \N__13416\,
            in3 => \N__14532\,
            lcout => \c0.n8449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33313\,
            in1 => \N__26461\,
            in2 => \N__17636\,
            in3 => \N__27936\,
            lcout => \c0.n20_adj_1659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i152_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21089\,
            in1 => \N__25170\,
            in2 => \_gnd_net_\,
            in3 => \N__29064\,
            lcout => data_in_field_151,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i21_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__13659\,
            in1 => \N__23564\,
            in2 => \N__18519\,
            in3 => \N__19149\,
            lcout => \c0.data_in_field_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14588\,
            in1 => \N__29616\,
            in2 => \_gnd_net_\,
            in3 => \N__16878\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7895_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__13658\,
            in1 => \N__32000\,
            in2 => \N__33031\,
            in3 => \N__18758\,
            lcout => \c0.n9578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_732_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16371\,
            in2 => \_gnd_net_\,
            in3 => \N__13657\,
            lcout => \c0.n8794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15027\,
            in1 => \N__14857\,
            in2 => \_gnd_net_\,
            in3 => \N__29615\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i27_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__23479\,
            in1 => \N__18551\,
            in2 => \N__19132\,
            in3 => \N__16846\,
            lcout => \c0.data_in_field_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i26_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__13566\,
            in1 => \N__23482\,
            in2 => \N__28244\,
            in3 => \N__19084\,
            lcout => \c0.data_in_field_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i33_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__23480\,
            in1 => \N__18715\,
            in2 => \N__19133\,
            in3 => \N__14781\,
            lcout => \c0.data_in_field_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i28_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__14994\,
            in1 => \N__23483\,
            in2 => \N__28299\,
            in3 => \N__19085\,
            lcout => \c0.data_in_field_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i3_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__23481\,
            in1 => \N__13689\,
            in2 => \N__19134\,
            in3 => \N__14941\,
            lcout => \c0.data_in_field_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_694_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13655\,
            in1 => \N__16358\,
            in2 => \_gnd_net_\,
            in3 => \N__16435\,
            lcout => \c0.n4381\,
            ltout => \c0.n4381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_685_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17069\,
            in1 => \N__13611\,
            in2 => \N__13662\,
            in3 => \N__14004\,
            lcout => \c0.n8899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_583_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13656\,
            in1 => \N__16806\,
            in2 => \N__13938\,
            in3 => \N__18711\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i1_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__14520\,
            in1 => \N__27982\,
            in2 => \N__23546\,
            in3 => \N__19045\,
            lcout => \c0.data_in_field_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i7_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__19040\,
            in1 => \N__13818\,
            in2 => \N__16378\,
            in3 => \N__23478\,
            lcout => \c0.data_in_field_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i34_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__23472\,
            in1 => \N__19041\,
            in2 => \N__13638\,
            in3 => \N__14905\,
            lcout => \c0.data_in_field_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_607_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13610\,
            in1 => \N__15300\,
            in2 => \N__21375\,
            in3 => \N__13953\,
            lcout => \c0.n4154\,
            ltout => \c0.n4154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_591_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13584\,
            in3 => \N__24785\,
            lcout => \c0.n4200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i6_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__19039\,
            in1 => \N__14556\,
            in2 => \N__21326\,
            in3 => \N__23477\,
            lcout => \c0.data_in_field_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_641_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15136\,
            in2 => \_gnd_net_\,
            in3 => \N__18642\,
            lcout => \c0.n8776\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i20_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__14664\,
            in1 => \N__23473\,
            in2 => \N__19127\,
            in3 => \N__13796\,
            lcout => \c0.data_in_field_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13876\,
            in1 => \N__15162\,
            in2 => \_gnd_net_\,
            in3 => \N__17006\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_594_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28292\,
            in1 => \N__13770\,
            in2 => \N__13764\,
            in3 => \N__15720\,
            lcout => \c0.n8427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i25_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__19046\,
            in1 => \N__14589\,
            in2 => \N__28079\,
            in3 => \N__23493\,
            lcout => \c0.data_in_field_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i10_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__13761\,
            in1 => \N__15294\,
            in2 => \N__23547\,
            in3 => \N__19053\,
            lcout => \c0.data_in_field_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i40_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__13737\,
            in1 => \N__23486\,
            in2 => \N__19129\,
            in3 => \N__14409\,
            lcout => \c0.data_in_field_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15375\,
            in1 => \N__23733\,
            in2 => \N__14637\,
            in3 => \N__13877\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i35_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__26982\,
            in1 => \N__23485\,
            in2 => \N__19128\,
            in3 => \N__17067\,
            lcout => \c0.data_in_field_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i5_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__18450\,
            in1 => \N__13931\,
            in2 => \N__23548\,
            in3 => \N__19054\,
            lcout => \c0.data_in_field_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i30_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__16554\,
            in1 => \N__23527\,
            in2 => \N__21429\,
            in3 => \N__19125\,
            lcout => \c0.data_in_field_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i8_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__23525\,
            in1 => \N__13908\,
            in2 => \N__19151\,
            in3 => \N__14003\,
            lcout => \c0.data_in_field_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_655_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28069\,
            in2 => \_gnd_net_\,
            in3 => \N__14399\,
            lcout => \c0.n4131\,
            ltout => \c0.n4131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_700_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13881\,
            in2 => \N__13863\,
            in3 => \N__22615\,
            lcout => \c0.n8927\,
            ltout => \c0.n8927_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__15371\,
            in1 => \N__18681\,
            in2 => \N__13860\,
            in3 => \N__17254\,
            lcout => \c0.n20_adj_1597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i48_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19120\,
            in1 => \N__13857\,
            in2 => \_gnd_net_\,
            in3 => \N__15837\,
            lcout => data_in_field_47,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i24_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__13845\,
            in1 => \N__23526\,
            in2 => \N__13980\,
            in3 => \N__19124\,
            lcout => \c0.data_in_field_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29380\,
            in1 => \N__14865\,
            in2 => \_gnd_net_\,
            in3 => \N__13817\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_637_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19817\,
            in2 => \_gnd_net_\,
            in3 => \N__27854\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i154_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25346\,
            in1 => \N__15753\,
            in2 => \N__14055\,
            in3 => \N__31469\,
            lcout => \c0.data_in_frame_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35346\,
            ce => \N__28996\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_8004_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__15421\,
            in1 => \N__33116\,
            in2 => \N__14052\,
            in3 => \N__32033\,
            lcout => OPEN,
            ltout => \c0.n9704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9704_bdd_4_lut_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33120\,
            in1 => \N__20629\,
            in2 => \N__14040\,
            in3 => \N__17709\,
            lcout => OPEN,
            ltout => \c0.n9707_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31378\,
            in1 => \N__14037\,
            in2 => \N__14022\,
            in3 => \N__31245\,
            lcout => \c0.n22_adj_1682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_8014_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__32032\,
            in1 => \N__13972\,
            in2 => \N__33175\,
            in3 => \N__16500\,
            lcout => OPEN,
            ltout => \c0.n9722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9722_bdd_4_lut_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33121\,
            in1 => \N__13999\,
            in2 => \N__14007\,
            in3 => \N__16953\,
            lcout => \c0.n9240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_661_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13971\,
            lcout => \c0.n4514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_513_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14079\,
            in1 => \N__14085\,
            in2 => \N__14073\,
            in3 => \N__15458\,
            lcout => OPEN,
            ltout => \c0.n18_adj_1589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_514_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24606\,
            in1 => \N__14135\,
            in2 => \N__14118\,
            in3 => \N__26082\,
            lcout => OPEN,
            ltout => \c0.n20_adj_1590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i167_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22097\,
            in1 => \N__24351\,
            in2 => \N__14115\,
            in3 => \N__18471\,
            lcout => \c0.data_in_frame_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35354\,
            ce => \N__29025\,
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_592_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14108\,
            in1 => \N__14094\,
            in2 => \_gnd_net_\,
            in3 => \N__22685\,
            lcout => \c0.n8822\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_651_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26397\,
            in2 => \_gnd_net_\,
            in3 => \N__25481\,
            lcout => \c0.n4448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_742_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32118\,
            in1 => \N__26619\,
            in2 => \_gnd_net_\,
            in3 => \N__17942\,
            lcout => \c0.n4445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_739_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17943\,
            in1 => \N__17450\,
            in2 => \N__26627\,
            in3 => \N__32119\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9650_bdd_4_lut_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__15537\,
            in1 => \N__17756\,
            in2 => \N__32555\,
            in3 => \N__33176\,
            lcout => \c0.n9126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i64_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17595\,
            in1 => \N__21591\,
            in2 => \_gnd_net_\,
            in3 => \N__28990\,
            lcout => data_in_field_63,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_717_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22016\,
            in1 => \N__22524\,
            in2 => \N__24960\,
            in3 => \N__27853\,
            lcout => \c0.n8896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i45_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22463\,
            in1 => \N__14187\,
            in2 => \_gnd_net_\,
            in3 => \N__19150\,
            lcout => data_in_field_44,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_627_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14176\,
            in2 => \_gnd_net_\,
            in3 => \N__18057\,
            lcout => \c0.n9016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i106_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__14177\,
            in1 => \_gnd_net_\,
            in2 => \N__19611\,
            in3 => \N__28986\,
            lcout => data_in_field_105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i128_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21590\,
            in1 => \_gnd_net_\,
            in2 => \N__29062\,
            in3 => \N__15558\,
            lcout => data_in_field_127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i74_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19610\,
            in1 => \N__24489\,
            in2 => \_gnd_net_\,
            in3 => \N__28991\,
            lcout => data_in_field_73,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_601_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18061\,
            in1 => \N__19684\,
            in2 => \N__19737\,
            in3 => \N__21627\,
            lcout => \c0.n8890\,
            ltout => \c0.n8890_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_606_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24713\,
            in1 => \N__15740\,
            in2 => \N__14163\,
            in3 => \N__22261\,
            lcout => \c0.n14_adj_1638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_720_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15666\,
            in1 => \N__22017\,
            in2 => \N__15441\,
            in3 => \N__21549\,
            lcout => \c0.n8936\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_600_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21550\,
            in1 => \N__15440\,
            in2 => \_gnd_net_\,
            in3 => \N__15667\,
            lcout => \c0.n4285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i136_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18062\,
            in1 => \N__21090\,
            in2 => \_gnd_net_\,
            in3 => \N__28992\,
            lcout => data_in_field_135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i84_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14245\,
            in1 => \_gnd_net_\,
            in2 => \N__29063\,
            in3 => \N__19440\,
            lcout => data_in_field_83,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_710_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17446\,
            in1 => \N__15870\,
            in2 => \_gnd_net_\,
            in3 => \N__14244\,
            lcout => \c0.n8785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7885_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33137\,
            in1 => \N__25275\,
            in2 => \N__21793\,
            in3 => \N__32031\,
            lcout => \c0.n9572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9656_bdd_4_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__33182\,
            in1 => \N__15636\,
            in2 => \N__17451\,
            in3 => \N__14193\,
            lcout => OPEN,
            ltout => \c0.n9123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_8009_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__14223\,
            in1 => \N__31627\,
            in2 => \N__14214\,
            in3 => \N__31244\,
            lcout => OPEN,
            ltout => \c0.n9644_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9644_bdd_4_lut_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31628\,
            in1 => \N__14211\,
            in2 => \N__14199\,
            in3 => \N__14376\,
            lcout => OPEN,
            ltout => \c0.n9647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i7_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__18111\,
            in1 => \N__31629\,
            in2 => \N__14196\,
            in3 => \N__32384\,
            lcout => \c0.tx2.r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35376\,
            ce => \N__32228\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7955_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__27728\,
            in1 => \N__33177\,
            in2 => \N__21949\,
            in3 => \N__32056\,
            lcout => \c0.n9656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__17679\,
            in1 => \N__17604\,
            in2 => \N__33203\,
            in3 => \N__32034\,
            lcout => OPEN,
            ltout => \c0.n9752_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9752_bdd_4_lut_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__33181\,
            in1 => \N__15841\,
            in2 => \N__14421\,
            in3 => \N__14418\,
            lcout => \c0.n9120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_7999_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__14370\,
            in1 => \N__32292\,
            in2 => \N__16109\,
            in3 => \N__16172\,
            lcout => OPEN,
            ltout => \c0.tx2.n9692_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n9692_bdd_4_lut_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__30054\,
            in1 => \N__14358\,
            in2 => \N__14346\,
            in3 => \N__16102\,
            lcout => OPEN,
            ltout => \c0.tx2.n9695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i590722_i1_3_lut_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14333\,
            in2 => \N__14343\,
            in3 => \N__15891\,
            lcout => OPEN,
            ltout => \c0.tx2.o_Tx_Serial_N_1511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010101"
        )
    port map (
            in0 => \N__14300\,
            in1 => \_gnd_net_\,
            in2 => \N__14340\,
            in3 => \N__15939\,
            lcout => n3_adj_1749,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i657_2_lut_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16173\,
            lcout => OPEN,
            ltout => \n2207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i2_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101000000000"
        )
    port map (
            in0 => \N__14334\,
            in1 => \N__16144\,
            in2 => \N__14337\,
            in3 => \N__16121\,
            lcout => \r_Bit_Index_2_adj_1741\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i2_2_lut_3_lut_4_lut_adj_507_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__15937\,
            in1 => \N__14299\,
            in2 => \N__26934\,
            in3 => \N__20475\,
            lcout => \c0.tx2.n3760\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i7729_3_lut_4_lut_4_lut_LC_3_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001000000010"
        )
    port map (
            in0 => \N__20474\,
            in1 => \N__15938\,
            in2 => \N__14316\,
            in3 => \N__14268\,
            lcout => n8747,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i138_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29395\,
            in1 => \N__20133\,
            in2 => \_gnd_net_\,
            in3 => \N__16016\,
            lcout => data_in_17_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i112_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29954\,
            in1 => \N__15993\,
            in2 => \_gnd_net_\,
            in3 => \N__14492\,
            lcout => data_in_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i127_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29697\,
            in1 => \N__14481\,
            in2 => \_gnd_net_\,
            in3 => \N__14624\,
            lcout => data_in_15_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i157_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29699\,
            in1 => \N__14601\,
            in2 => \_gnd_net_\,
            in3 => \N__16286\,
            lcout => data_in_19_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i135_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29698\,
            in1 => \N__18159\,
            in2 => \_gnd_net_\,
            in3 => \N__14480\,
            lcout => data_in_16_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i79_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14460\,
            in1 => \N__29769\,
            in2 => \_gnd_net_\,
            in3 => \N__14471\,
            lcout => data_in_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i87_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__14451\,
            in1 => \_gnd_net_\,
            in2 => \N__29955\,
            in3 => \N__14459\,
            lcout => data_in_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i95_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14430\,
            in1 => \N__29770\,
            in2 => \_gnd_net_\,
            in3 => \N__14450\,
            lcout => data_in_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i103_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29766\,
            in1 => \N__14442\,
            in2 => \_gnd_net_\,
            in3 => \N__14429\,
            lcout => data_in_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i119_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29767\,
            in1 => \N__14625\,
            in2 => \_gnd_net_\,
            in3 => \N__14612\,
            lcout => data_in_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14583\,
            in1 => \N__14777\,
            in2 => \_gnd_net_\,
            in3 => \N__29774\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i165_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29768\,
            in1 => \N__20418\,
            in2 => \_gnd_net_\,
            in3 => \N__14600\,
            lcout => data_in_20_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_678_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15018\,
            in1 => \N__16542\,
            in2 => \N__14584\,
            in3 => \N__14551\,
            lcout => OPEN,
            ltout => \c0.n28_adj_1668_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_684_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__16518\,
            in2 => \N__14535\,
            in3 => \N__14526\,
            lcout => \c0.n30_adj_1674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_2_lut_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18573\,
            in2 => \_gnd_net_\,
            in3 => \N__14512\,
            lcout => \c0.n22_adj_1667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15022\,
            in1 => \N__16520\,
            in2 => \_gnd_net_\,
            in3 => \N__29393\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__16519\,
            in1 => \_gnd_net_\,
            in2 => \N__29623\,
            in3 => \N__16196\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14513\,
            in1 => \N__29389\,
            in2 => \_gnd_net_\,
            in3 => \N__15267\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i105_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29388\,
            in1 => \N__14792\,
            in2 => \_gnd_net_\,
            in3 => \N__18411\,
            lcout => data_in_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i33_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29840\,
            in1 => \N__14776\,
            in2 => \_gnd_net_\,
            in3 => \N__20526\,
            lcout => data_in_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_681_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18379\,
            in1 => \N__19185\,
            in2 => \N__16879\,
            in3 => \N__15263\,
            lcout => \c0.n13_adj_1671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_682_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15100\,
            in1 => \N__14652\,
            in2 => \N__16255\,
            in3 => \N__14679\,
            lcout => \c0.n13_adj_1672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18380\,
            in1 => \N__29956\,
            in2 => \_gnd_net_\,
            in3 => \N__14733\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i44_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__14709\,
            in1 => \_gnd_net_\,
            in2 => \N__30028\,
            in3 => \N__15211\,
            lcout => data_in_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__14680\,
            in1 => \N__29964\,
            in2 => \N__14660\,
            in3 => \_gnd_net_\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__15101\,
            in1 => \_gnd_net_\,
            in2 => \N__30029\,
            in3 => \N__14681\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14653\,
            in1 => \N__29957\,
            in2 => \_gnd_net_\,
            in3 => \N__14989\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_572_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21234\,
            in2 => \_gnd_net_\,
            in3 => \N__25166\,
            lcout => \c0.n4495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i22_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__23560\,
            in1 => \N__19066\,
            in2 => \N__16263\,
            in3 => \N__21357\,
            lcout => \c0.data_in_field_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_614_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16458\,
            in2 => \_gnd_net_\,
            in3 => \N__14934\,
            lcout => \c0.n8902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_708_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14897\,
            in1 => \N__15063\,
            in2 => \_gnd_net_\,
            in3 => \N__28041\,
            lcout => OPEN,
            ltout => \c0.n6_adj_1632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_596_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16697\,
            in1 => \N__16805\,
            in2 => \N__14874\,
            in3 => \N__14871\,
            lcout => \c0.n4107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_695_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16487\,
            lcout => \c0.n8804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i15_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__14861\,
            in1 => \N__23562\,
            in2 => \N__16413\,
            in3 => \N__19088\,
            lcout => \c0.data_in_field_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i32_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__23561\,
            in1 => \N__19067\,
            in2 => \N__14835\,
            in3 => \N__16488\,
            lcout => \c0.data_in_field_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i19_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__18384\,
            in1 => \N__23563\,
            in2 => \N__16818\,
            in3 => \N__19089\,
            lcout => \c0.data_in_field_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i39_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__16203\,
            in1 => \N__23470\,
            in2 => \N__22619\,
            in3 => \N__19087\,
            lcout => \c0.data_in_field_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_728_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18636\,
            in2 => \_gnd_net_\,
            in3 => \N__25603\,
            lcout => \c0.n4127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i4_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__19065\,
            in1 => \N__23471\,
            in2 => \N__15108\,
            in3 => \N__15084\,
            lcout => \c0.data_in_field_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_534_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15045\,
            in1 => \N__15036\,
            in2 => \N__16659\,
            in3 => \N__17019\,
            lcout => \c0.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i38_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__25604\,
            in1 => \N__23469\,
            in2 => \N__18300\,
            in3 => \N__19086\,
            lcout => data_in_field_37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7399_4_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__23668\,
            in1 => \N__20822\,
            in2 => \N__23545\,
            in3 => \N__20776\,
            lcout => n9069,
            ltout => \n9069_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i23_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__15026\,
            in1 => \N__23468\,
            in2 => \N__14997\,
            in3 => \N__16439\,
            lcout => \c0.data_in_field_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29394\,
            in1 => \N__15185\,
            in2 => \_gnd_net_\,
            in3 => \N__14985\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22778\,
            in1 => \_gnd_net_\,
            in2 => \N__25612\,
            in3 => \N__18640\,
            lcout => OPEN,
            ltout => \n4_adj_1750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__25640\,
            in1 => \N__14958\,
            in2 => \N__14949\,
            in3 => \N__18858\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i52_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15327\,
            in1 => \N__17501\,
            in2 => \_gnd_net_\,
            in3 => \N__19064\,
            lcout => data_in_field_51,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i53_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25262\,
            in1 => \N__19126\,
            in2 => \_gnd_net_\,
            in3 => \N__15315\,
            lcout => data_in_field_52,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_650_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22777\,
            in1 => \N__22604\,
            in2 => \N__25611\,
            in3 => \N__28009\,
            lcout => \c0.n8831\,
            ltout => \c0.n8831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_656_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15160\,
            in1 => \N__15292\,
            in2 => \N__15270\,
            in3 => \N__16434\,
            lcout => \c0.n4183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i9_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__15262\,
            in1 => \N__23451\,
            in2 => \N__28019\,
            in3 => \N__19063\,
            lcout => \c0.data_in_field_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i56_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19062\,
            in1 => \N__15231\,
            in2 => \_gnd_net_\,
            in3 => \N__17671\,
            lcout => data_in_field_55,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i36_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15178\,
            in1 => \N__29624\,
            in2 => \_gnd_net_\,
            in3 => \N__15216\,
            lcout => data_in_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_554_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24442\,
            in1 => \N__15414\,
            in2 => \_gnd_net_\,
            in3 => \N__22728\,
            lcout => \c0.n4556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_609_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18606\,
            in1 => \N__15161\,
            in2 => \N__15144\,
            in3 => \N__17153\,
            lcout => OPEN,
            ltout => \c0.n10_adj_1640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22675\,
            in1 => \N__16412\,
            in2 => \N__15477\,
            in3 => \N__15474\,
            lcout => \c0.n8933\,
            ltout => \c0.n8933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21410\,
            in2 => \N__15462\,
            in3 => \N__15491\,
            lcout => OPEN,
            ltout => \c0.n8314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_538_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111001"
        )
    port map (
            in0 => \N__24441\,
            in1 => \N__15459\,
            in2 => \N__15444\,
            in3 => \N__27233\,
            lcout => \c0.n23_adj_1608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i146_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15415\,
            in1 => \_gnd_net_\,
            in2 => \N__21044\,
            in3 => \N__28772\,
            lcout => data_in_field_145,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_555_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21233\,
            in1 => \N__15386\,
            in2 => \N__15568\,
            in3 => \N__17125\,
            lcout => \c0.n8974\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_645_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22468\,
            lcout => \c0.n8861\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_526_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22407\,
            in2 => \_gnd_net_\,
            in3 => \N__17124\,
            lcout => \c0.n4452\,
            ltout => \c0.n4452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23762\,
            in1 => \N__15360\,
            in2 => \N__15354\,
            in3 => \N__17393\,
            lcout => \c0.n8906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_702_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__21881\,
            in1 => \_gnd_net_\,
            in2 => \N__15569\,
            in3 => \N__24943\,
            lcout => \c0.n4253\,
            ltout => \c0.n4253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_531_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23845\,
            in1 => \N__15645\,
            in2 => \N__15639\,
            in3 => \N__15635\,
            lcout => \c0.n24_adj_1607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i148_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21155\,
            in2 => \N__29055\,
            in3 => \N__15594\,
            lcout => data_in_field_147,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i132_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__21154\,
            in1 => \_gnd_net_\,
            in2 => \N__23775\,
            in3 => \N__28968\,
            lcout => data_in_field_131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7950_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__32007\,
            in1 => \N__33189\,
            in2 => \N__15570\,
            in3 => \N__25741\,
            lcout => \c0.n9650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_4_lut_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26690\,
            in1 => \N__17541\,
            in2 => \N__21126\,
            in3 => \N__17593\,
            lcout => \c0.n16_adj_1598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_734_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17540\,
            in1 => \N__17594\,
            in2 => \_gnd_net_\,
            in3 => \N__26689\,
            lcout => \c0.n8980\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i60_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26728\,
            in1 => \N__17542\,
            in2 => \_gnd_net_\,
            in3 => \N__28972\,
            lcout => data_in_field_59,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_633_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25740\,
            lcout => OPEN,
            ltout => \c0.n6_adj_1645_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_634_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15518\,
            in1 => \N__21690\,
            in2 => \N__15498\,
            in3 => \N__15495\,
            lcout => \c0.n8788\,
            ltout => \c0.n8788_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_638_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27269\,
            in1 => \N__32508\,
            in2 => \N__15756\,
            in3 => \N__25553\,
            lcout => \c0.n14_adj_1648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_523_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26291\,
            in1 => \N__26031\,
            in2 => \N__15747\,
            in3 => \N__21821\,
            lcout => OPEN,
            ltout => \c0.n24_adj_1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15726\,
            in1 => \N__26556\,
            in2 => \N__15729\,
            in3 => \N__24860\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25718\,
            in1 => \N__21880\,
            in2 => \_gnd_net_\,
            in3 => \N__24948\,
            lcout => \c0.n18_adj_1603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_605_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22467\,
            in2 => \_gnd_net_\,
            in3 => \N__15719\,
            lcout => \c0.tx2_transmit_N_1334\,
            ltout => \c0.tx2_transmit_N_1334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_524_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28344\,
            in1 => \N__22749\,
            in2 => \N__15702\,
            in3 => \N__24903\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1601_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i165_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15699\,
            in1 => \N__18009\,
            in2 => \N__15690\,
            in3 => \N__15687\,
            lcout => \c0.data_in_frame_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35370\,
            ce => \N__28997\,
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15801\,
            in1 => \N__19927\,
            in2 => \N__21966\,
            in3 => \N__15879\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i116_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19439\,
            in1 => \N__15668\,
            in2 => \_gnd_net_\,
            in3 => \N__28985\,
            lcout => data_in_field_115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_648_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19473\,
            in2 => \_gnd_net_\,
            in3 => \N__25276\,
            lcout => OPEN,
            ltout => \c0.n4574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_558_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25808\,
            in1 => \N__21787\,
            in2 => \N__15882\,
            in3 => \N__26345\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17435\,
            in2 => \_gnd_net_\,
            in3 => \N__15878\,
            lcout => \c0.n24_adj_1615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i105_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19474\,
            in1 => \N__20675\,
            in2 => \_gnd_net_\,
            in3 => \N__28984\,
            lcout => data_in_field_104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_539_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26206\,
            in2 => \_gnd_net_\,
            in3 => \N__27879\,
            lcout => \c0.n8909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_613_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21432\,
            in2 => \_gnd_net_\,
            in3 => \N__15846\,
            lcout => \c0.n8945\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_570_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24183\,
            in2 => \_gnd_net_\,
            in3 => \N__24299\,
            lcout => \c0.n8825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_552_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__21891\,
            in1 => \_gnd_net_\,
            in2 => \N__20750\,
            in3 => \N__21730\,
            lcout => \c0.n4333\,
            ltout => \c0.n4333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_729_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__24300\,
            in1 => \_gnd_net_\,
            in2 => \N__15795\,
            in3 => \N__27328\,
            lcout => \c0.n8998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_45_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__26938\,
            in1 => \N__15769\,
            in2 => \_gnd_net_\,
            in3 => \N__15792\,
            lcout => tx2_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_559_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31685\,
            in1 => \N__15963\,
            in2 => \N__23916\,
            in3 => \N__15957\,
            lcout => \c0.n38_adj_1616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21554\,
            in1 => \N__27098\,
            in2 => \_gnd_net_\,
            in3 => \N__21731\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_47_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110000"
        )
    port map (
            in0 => \N__26943\,
            in1 => \N__15951\,
            in2 => \N__20495\,
            in3 => \N__15906\,
            lcout => tx2_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__15900\,
            in1 => \N__22872\,
            in2 => \N__16107\,
            in3 => \N__16171\,
            lcout => OPEN,
            ltout => \c0.tx2.n9716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.n9716_bdd_4_lut_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__25365\,
            in1 => \N__20010\,
            in2 => \N__15894\,
            in3 => \N__16095\,
            lcout => \c0.tx2.n9719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i0_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__16177\,
            in1 => \N__16145\,
            in2 => \_gnd_net_\,
            in3 => \N__16127\,
            lcout => \r_Bit_Index_0_adj_1743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_4_lut_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001010101"
        )
    port map (
            in0 => \N__30789\,
            in1 => \N__30647\,
            in2 => \N__30579\,
            in3 => \N__30723\,
            lcout => OPEN,
            ltout => \n4691_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__30648\,
            in1 => \N__29254\,
            in2 => \N__15885\,
            in3 => \N__30790\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7769_2_lut_3_lut_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__30788\,
            in1 => \N__30646\,
            in2 => \_gnd_net_\,
            in3 => \N__30722\,
            lcout => n8761,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_i1_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__16178\,
            in1 => \N__16146\,
            in2 => \N__16108\,
            in3 => \N__16128\,
            lcout => \r_Bit_Index_1_adj_1742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i122_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29883\,
            in1 => \N__16005\,
            in2 => \_gnd_net_\,
            in3 => \N__16061\,
            lcout => data_in_15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i132_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29953\,
            in1 => \N__18210\,
            in2 => \_gnd_net_\,
            in3 => \N__18230\,
            lcout => data_in_16_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i141_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29884\,
            in1 => \N__16275\,
            in2 => \_gnd_net_\,
            in3 => \N__16316\,
            lcout => data_in_17_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i37_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29885\,
            in1 => \N__16900\,
            in2 => \_gnd_net_\,
            in3 => \N__16049\,
            lcout => data_in_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i130_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16017\,
            in1 => \N__29886\,
            in2 => \_gnd_net_\,
            in3 => \N__16004\,
            lcout => data_in_16_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i120_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15981\,
            in1 => \N__29645\,
            in2 => \_gnd_net_\,
            in3 => \N__15992\,
            lcout => data_in_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i128_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15972\,
            in1 => \N__29649\,
            in2 => \_gnd_net_\,
            in3 => \N__15980\,
            lcout => data_in_15_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i136_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29647\,
            in1 => \N__16296\,
            in2 => \_gnd_net_\,
            in3 => \N__15971\,
            lcout => data_in_16_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i125_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__29646\,
            in2 => \_gnd_net_\,
            in3 => \N__16328\,
            lcout => data_in_15_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i133_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29643\,
            in1 => \N__16317\,
            in2 => \_gnd_net_\,
            in3 => \N__16304\,
            lcout => data_in_16_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i144_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29648\,
            in1 => \N__20226\,
            in2 => \_gnd_net_\,
            in3 => \N__16295\,
            lcout => data_in_17_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i149_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29644\,
            in1 => \N__16287\,
            in2 => \_gnd_net_\,
            in3 => \N__16274\,
            lcout => data_in_18_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16544\,
            in1 => \N__29795\,
            in2 => \_gnd_net_\,
            in3 => \N__16254\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i47_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16596\,
            in1 => \_gnd_net_\,
            in2 => \N__29965\,
            in3 => \N__16219\,
            lcout => data_in_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i39_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16220\,
            in1 => \N__29796\,
            in2 => \_gnd_net_\,
            in3 => \N__16195\,
            lcout => data_in_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29793\,
            in1 => \N__16907\,
            in2 => \_gnd_net_\,
            in3 => \N__18578\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i55_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16562\,
            in1 => \N__29800\,
            in2 => \_gnd_net_\,
            in3 => \N__16595\,
            lcout => data_in_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_54_i1_3_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16594\,
            in1 => \N__20879\,
            in2 => \_gnd_net_\,
            in3 => \N__23542\,
            lcout => n1889,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i63_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__16584\,
            in1 => \N__29801\,
            in2 => \N__16566\,
            in3 => \_gnd_net_\,
            lcout => data_in_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29794\,
            in1 => \N__18289\,
            in2 => \_gnd_net_\,
            in3 => \N__16543\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i31_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__16461\,
            in1 => \N__23553\,
            in2 => \N__16524\,
            in3 => \N__19119\,
            lcout => \c0.data_in_field_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_690_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22672\,
            in1 => \N__16616\,
            in2 => \N__16411\,
            in3 => \N__28042\,
            lcout => \c0.n8843\,
            ltout => \c0.n8843_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_621_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18743\,
            in1 => \N__18677\,
            in2 => \N__16503\,
            in3 => \N__16489\,
            lcout => \c0.n4151\,
            ltout => \c0.n4151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_623_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21430\,
            in1 => \N__27989\,
            in2 => \N__16464\,
            in3 => \N__16459\,
            lcout => \c0.n8852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7945_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__16460\,
            in1 => \N__32013\,
            in2 => \N__33032\,
            in3 => \N__16443\,
            lcout => OPEN,
            ltout => \c0.n9638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9638_bdd_4_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__16404\,
            in1 => \N__32955\,
            in2 => \N__16383\,
            in3 => \N__16380\,
            lcout => \c0.n9132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i17_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__28043\,
            in1 => \N__23554\,
            in2 => \N__16884\,
            in3 => \N__19118\,
            lcout => \c0.data_in_field_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i29_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__19117\,
            in1 => \N__18577\,
            in2 => \N__23565\,
            in3 => \N__18744\,
            lcout => \c0.data_in_field_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7910_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__32957\,
            in1 => \N__32012\,
            in2 => \N__21735\,
            in3 => \N__22147\,
            lcout => \c0.n9602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7840_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__32011\,
            in1 => \N__16848\,
            in2 => \N__16817\,
            in3 => \N__32956\,
            lcout => \c0.n9512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i18_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__16764\,
            in1 => \N__23501\,
            in2 => \N__19130\,
            in3 => \N__17304\,
            lcout => \c0.data_in_field_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_616_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16945\,
            in2 => \_gnd_net_\,
            in3 => \N__16614\,
            lcout => \c0.n4492\,
            ltout => \c0.n4492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_617_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16716\,
            in1 => \N__16698\,
            in2 => \N__16686\,
            in3 => \N__22991\,
            lcout => \c0.n8948\,
            ltout => \c0.n8948_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_525_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__22146\,
            in1 => \N__25019\,
            in2 => \N__16683\,
            in3 => \N__16676\,
            lcout => \c0.n19_adj_1602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i2_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__16615\,
            in1 => \N__23502\,
            in2 => \N__19131\,
            in3 => \N__16650\,
            lcout => \c0.data_in_field_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i16_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__16980\,
            in1 => \N__16946\,
            in2 => \N__23552\,
            in3 => \N__19074\,
            lcout => \c0.data_in_field_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i43_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19056\,
            in1 => \N__22923\,
            in2 => \_gnd_net_\,
            in3 => \N__18676\,
            lcout => data_in_field_42,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_48_i1_3_lut_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23506\,
            in1 => \_gnd_net_\,
            in2 => \N__20561\,
            in3 => \N__24128\,
            lcout => OPEN,
            ltout => \n1895_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i49_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19058\,
            in1 => \_gnd_net_\,
            in2 => \N__16932\,
            in3 => \N__19213\,
            lcout => data_in_field_48,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i55_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16929\,
            in1 => \N__24437\,
            in2 => \_gnd_net_\,
            in3 => \N__19061\,
            lcout => data_in_field_54,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i47_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19057\,
            in1 => \N__16920\,
            in2 => \_gnd_net_\,
            in3 => \N__22671\,
            lcout => data_in_field_46,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i37_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__23507\,
            in1 => \N__16908\,
            in2 => \N__22804\,
            in3 => \N__19059\,
            lcout => data_in_field_36,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i41_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19055\,
            in1 => \N__20643\,
            in2 => \_gnd_net_\,
            in3 => \N__18641\,
            lcout => data_in_field_40,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i51_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23202\,
            in1 => \N__26814\,
            in2 => \_gnd_net_\,
            in3 => \N__19060\,
            lcout => data_in_field_50,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7830_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__32883\,
            in1 => \N__26816\,
            in2 => \N__32035\,
            in3 => \N__24033\,
            lcout => OPEN,
            ltout => \c0.n9506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9506_bdd_4_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32890\,
            in1 => \N__18675\,
            in2 => \N__17073\,
            in3 => \N__17070\,
            lcout => \c0.n9195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_516_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17664\,
            lcout => OPEN,
            ltout => \c0.n4_adj_1592_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_522_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001101111"
        )
    port map (
            in0 => \N__26815\,
            in1 => \N__27119\,
            in2 => \N__17034\,
            in3 => \N__17031\,
            lcout => \c0.n21_adj_1599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i81_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24129\,
            in1 => \N__27930\,
            in2 => \_gnd_net_\,
            in3 => \N__28673\,
            lcout => data_in_field_80,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17136\,
            in1 => \N__17013\,
            in2 => \N__16995\,
            in3 => \N__16986\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i57_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20921\,
            in1 => \_gnd_net_\,
            in2 => \N__28749\,
            in3 => \N__24213\,
            lcout => data_in_field_56,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i140_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26739\,
            in1 => \N__17394\,
            in2 => \_gnd_net_\,
            in3 => \N__28578\,
            lcout => data_in_field_139,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i95_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__19365\,
            in1 => \_gnd_net_\,
            in2 => \N__28751\,
            in3 => \N__22523\,
            lcout => data_in_field_94,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_512_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23012\,
            in1 => \N__17235\,
            in2 => \N__17217\,
            in3 => \N__17205\,
            lcout => OPEN,
            ltout => \c0.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17190\,
            in2 => \N__17178\,
            in3 => \N__17175\,
            lcout => OPEN,
            ltout => \c0.n8421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_529_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111101"
        )
    port map (
            in0 => \N__25250\,
            in1 => \N__17163\,
            in2 => \N__17157\,
            in3 => \N__17154\,
            lcout => \c0.n24_adj_1605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i78_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22411\,
            in1 => \_gnd_net_\,
            in2 => \N__28750\,
            in3 => \N__21278\,
            lcout => data_in_field_77,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i93_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29108\,
            in1 => \N__24944\,
            in2 => \_gnd_net_\,
            in3 => \N__28585\,
            lcout => data_in_field_92,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i76_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19552\,
            in1 => \N__17126\,
            in2 => \_gnd_net_\,
            in3 => \N__28665\,
            lcout => data_in_field_75,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i79_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22304\,
            in2 => \N__28854\,
            in3 => \N__26381\,
            lcout => data_in_field_78,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i94_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21464\,
            in1 => \N__22000\,
            in2 => \_gnd_net_\,
            in3 => \N__28672\,
            lcout => data_in_field_93,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i68_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21156\,
            in1 => \_gnd_net_\,
            in2 => \N__28853\,
            in3 => \N__17097\,
            lcout => data_in_field_67,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i120_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19722\,
            in1 => \N__25745\,
            in2 => \_gnd_net_\,
            in3 => \N__28658\,
            lcout => data_in_field_119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i63_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19354\,
            in2 => \N__28852\,
            in3 => \N__22715\,
            lcout => data_in_field_62,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_647_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17340\,
            in1 => \N__17331\,
            in2 => \N__27621\,
            in3 => \N__19781\,
            lcout => \c0.n8939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i92_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26721\,
            in1 => \_gnd_net_\,
            in2 => \N__28855\,
            in3 => \N__21873\,
            lcout => data_in_field_91,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_727_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25220\,
            in1 => \N__21225\,
            in2 => \_gnd_net_\,
            in3 => \N__17703\,
            lcout => \c0.n8992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22562\,
            in1 => \N__21807\,
            in2 => \N__17325\,
            in3 => \N__17311\,
            lcout => \c0.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i86_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19676\,
            in1 => \N__19882\,
            in2 => \_gnd_net_\,
            in3 => \N__28885\,
            lcout => data_in_field_85,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i61_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29097\,
            in2 => \N__29011\,
            in3 => \N__21774\,
            lcout => data_in_field_60,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i142_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21459\,
            in1 => \N__19920\,
            in2 => \_gnd_net_\,
            in3 => \N__28881\,
            lcout => data_in_field_141,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_622_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23851\,
            in1 => \N__20739\,
            in2 => \N__21750\,
            in3 => \N__17261\,
            lcout => \c0.n19_adj_1643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i127_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19353\,
            in1 => \N__22563\,
            in2 => \_gnd_net_\,
            in3 => \N__28877\,
            lcout => data_in_field_126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i138_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__17704\,
            in1 => \_gnd_net_\,
            in2 => \N__29010\,
            in3 => \N__21661\,
            lcout => data_in_field_137,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_644_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17602\,
            in1 => \N__31419\,
            in2 => \N__17550\,
            in3 => \N__21623\,
            lcout => \c0.n22_adj_1617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i73_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20671\,
            in2 => \N__29014\,
            in3 => \N__27886\,
            lcout => data_in_field_72,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i137_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20916\,
            in1 => \N__26212\,
            in2 => \_gnd_net_\,
            in3 => \N__28892\,
            lcout => data_in_field_136,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_604_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17643\,
            in1 => \N__17885\,
            in2 => \N__20749\,
            in3 => \N__17510\,
            lcout => \c0.n4302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i80_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19501\,
            in1 => \N__17436\,
            in2 => \_gnd_net_\,
            in3 => \N__28896\,
            lcout => data_in_field_79,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_726_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23849\,
            in1 => \N__27784\,
            in2 => \N__17402\,
            in3 => \N__17357\,
            lcout => \c0.n8782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_709_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27785\,
            in1 => \N__23850\,
            in2 => \_gnd_net_\,
            in3 => \N__22516\,
            lcout => \c0.n8977\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i112_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19500\,
            in2 => \N__29013\,
            in3 => \N__17755\,
            lcout => data_in_field_111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_718_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25334\,
            in1 => \N__25219\,
            in2 => \N__19782\,
            in3 => \N__22327\,
            lcout => \c0.n4525\,
            ltout => \c0.n4525_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_557_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19677\,
            in1 => \N__17913\,
            in2 => \N__17736\,
            in3 => \N__22570\,
            lcout => \c0.n8924\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_589_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17733\,
            in2 => \_gnd_net_\,
            in3 => \N__17705\,
            lcout => \c0.n8874\,
            ltout => \c0.n8874_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_560_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22245\,
            in1 => \N__27137\,
            in2 => \N__17682\,
            in3 => \N__25722\,
            lcout => \c0.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_602_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24390\,
            in2 => \_gnd_net_\,
            in3 => \N__17678\,
            lcout => \c0.n6_adj_1636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i134_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19304\,
            in1 => \N__32586\,
            in2 => \_gnd_net_\,
            in3 => \N__29057\,
            lcout => data_in_field_133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_701_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19475\,
            in1 => \N__25277\,
            in2 => \_gnd_net_\,
            in3 => \N__27045\,
            lcout => \c0.n8989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i70_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24391\,
            in1 => \N__19299\,
            in2 => \_gnd_net_\,
            in3 => \N__29058\,
            lcout => data_in_field_69,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_528_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17912\,
            in2 => \_gnd_net_\,
            in3 => \N__21928\,
            lcout => OPEN,
            ltout => \c0.n6_adj_1604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_530_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24047\,
            in1 => \N__22729\,
            in2 => \N__18012\,
            in3 => \N__27429\,
            lcout => \c0.n8983\,
            ltout => \c0.n8983_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17997\,
            in1 => \N__17985\,
            in2 => \N__17976\,
            in3 => \N__17973\,
            lcout => \c0.n26_adj_1606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_556_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17954\,
            in1 => \N__25139\,
            in2 => \N__26462\,
            in3 => \N__32121\,
            lcout => \c0.n4203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_532_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17898\,
            in1 => \N__26115\,
            in2 => \N__20583\,
            in3 => \N__17886\,
            lcout => OPEN,
            ltout => \c0.n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i164_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17874\,
            in1 => \N__17862\,
            in2 => \N__17856\,
            in3 => \N__17853\,
            lcout => \c0.data_in_frame_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35392\,
            ce => \N__29021\,
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_561_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24365\,
            in1 => \N__17828\,
            in2 => \N__17805\,
            in3 => \N__17790\,
            lcout => \c0.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1509_2_lut_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32045\,
            in2 => \_gnd_net_\,
            in3 => \N__33138\,
            lcout => \c0.n3056\,
            ltout => \c0.n3056_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__17778\,
            in1 => \N__18036\,
            in2 => \N__18114\,
            in3 => \N__31263\,
            lcout => \c0.n22_adj_1676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i160_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24999\,
            in1 => \N__18099\,
            in2 => \N__18093\,
            in3 => \N__18081\,
            lcout => \c0.data_in_frame_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35398\,
            ce => \N__29072\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7960_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25213\,
            in1 => \N__33148\,
            in2 => \N__18075\,
            in3 => \N__32046\,
            lcout => OPEN,
            ltout => \c0.n9662_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9662_bdd_4_lut_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33149\,
            in1 => \N__18066\,
            in2 => \N__18039\,
            in3 => \N__21555\,
            lcout => \c0.n9665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i84_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29975\,
            in1 => \N__20070\,
            in2 => \_gnd_net_\,
            in3 => \N__18140\,
            lcout => data_in_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i110_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29966\,
            in1 => \N__19973\,
            in2 => \_gnd_net_\,
            in3 => \N__19953\,
            lcout => data_in_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i100_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18030\,
            in1 => \N__29969\,
            in2 => \_gnd_net_\,
            in3 => \N__20081\,
            lcout => data_in_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i108_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18021\,
            in1 => \N__29976\,
            in2 => \_gnd_net_\,
            in3 => \N__18029\,
            lcout => data_in_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i116_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18219\,
            in1 => \N__29970\,
            in2 => \_gnd_net_\,
            in3 => \N__18020\,
            lcout => data_in_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i124_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29967\,
            in1 => \N__18231\,
            in2 => \_gnd_net_\,
            in3 => \N__18218\,
            lcout => data_in_15_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i140_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29968\,
            in1 => \N__18198\,
            in2 => \_gnd_net_\,
            in3 => \N__18209\,
            lcout => data_in_17_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i148_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18186\,
            in1 => \N__29652\,
            in2 => \_gnd_net_\,
            in3 => \N__18197\,
            lcout => data_in_18_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i156_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18177\,
            in1 => \N__29654\,
            in2 => \_gnd_net_\,
            in3 => \N__18185\,
            lcout => data_in_19_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i164_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29656\,
            in1 => \N__20271\,
            in2 => \_gnd_net_\,
            in3 => \N__18176\,
            lcout => data_in_20_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i150_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18168\,
            in1 => \N__29653\,
            in2 => \_gnd_net_\,
            in3 => \N__20165\,
            lcout => data_in_18_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i158_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29655\,
            in1 => \N__18324\,
            in2 => \_gnd_net_\,
            in3 => \N__18167\,
            lcout => data_in_19_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i143_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29651\,
            in1 => \N__20145\,
            in2 => \_gnd_net_\,
            in3 => \N__18155\,
            lcout => data_in_17_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35314\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_31_i4_2_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27552\,
            in2 => \_gnd_net_\,
            in3 => \N__25874\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i76_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29924\,
            in1 => \N__18125\,
            in2 => \_gnd_net_\,
            in3 => \N__18144\,
            lcout => data_in_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i166_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29923\,
            in1 => \N__20351\,
            in2 => \_gnd_net_\,
            in3 => \N__18323\,
            lcout => data_in_20_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_45_i1_3_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21274\,
            in1 => \N__18310\,
            in2 => \_gnd_net_\,
            in3 => \N__23543\,
            lcout => n1898,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i46_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18311\,
            in1 => \N__29803\,
            in2 => \_gnd_net_\,
            in3 => \N__18270\,
            lcout => data_in_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i38_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29802\,
            in1 => \N__18312\,
            in2 => \_gnd_net_\,
            in3 => \N__18290\,
            lcout => data_in_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i54_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29838\,
            in1 => \N__18258\,
            in2 => \_gnd_net_\,
            in3 => \N__18269\,
            lcout => data_in_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_53_i1_3_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18268\,
            in1 => \N__19887\,
            in2 => \_gnd_net_\,
            in3 => \N__23544\,
            lcout => n1890,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i62_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18249\,
            in1 => \N__29804\,
            in2 => \_gnd_net_\,
            in3 => \N__18257\,
            lcout => data_in_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i70_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18240\,
            in1 => \N__29837\,
            in2 => \_gnd_net_\,
            in3 => \N__18248\,
            lcout => data_in_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i78_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29839\,
            in1 => \N__18239\,
            in2 => \_gnd_net_\,
            in3 => \N__20001\,
            lcout => data_in_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35328\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i113_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18393\,
            in1 => \N__29983\,
            in2 => \_gnd_net_\,
            in3 => \N__18404\,
            lcout => data_in_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i121_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29980\,
            in1 => \N__18354\,
            in2 => \_gnd_net_\,
            in3 => \N__18392\,
            lcout => data_in_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i135_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24657\,
            in1 => \N__25784\,
            in2 => \_gnd_net_\,
            in3 => \N__29012\,
            lcout => data_in_field_134,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29982\,
            in1 => \N__18544\,
            in2 => \_gnd_net_\,
            in3 => \N__18375\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i153_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18341\,
            in1 => \N__29984\,
            in2 => \_gnd_net_\,
            in3 => \N__29147\,
            lcout => data_in_19_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i129_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29981\,
            in1 => \N__18483\,
            in2 => \_gnd_net_\,
            in3 => \N__18353\,
            lcout => data_in_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i161_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__20247\,
            in1 => \N__29985\,
            in2 => \N__18345\,
            in3 => \_gnd_net_\,
            lcout => data_in_20_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i46_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18333\,
            in1 => \N__18850\,
            in2 => \_gnd_net_\,
            in3 => \N__19148\,
            lcout => data_in_field_45,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_8029_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__31910\,
            in1 => \N__32871\,
            in2 => \N__19215\,
            in3 => \N__24223\,
            lcout => OPEN,
            ltout => \c0.n9746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9746_bdd_4_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__18635\,
            in1 => \N__32872\,
            in2 => \N__18720\,
            in3 => \N__18717\,
            lcout => \c0.n9228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_686_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18801\,
            in1 => \N__18668\,
            in2 => \_gnd_net_\,
            in3 => \N__18634\,
            lcout => \c0.n4208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18582\,
            in1 => \N__18507\,
            in2 => \_gnd_net_\,
            in3 => \N__29873\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29871\,
            in1 => \N__26978\,
            in2 => \_gnd_net_\,
            in3 => \N__18543\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19181\,
            in1 => \N__18508\,
            in2 => \_gnd_net_\,
            in3 => \N__29872\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i137_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29870\,
            in1 => \N__29136\,
            in2 => \_gnd_net_\,
            in3 => \N__18482\,
            lcout => data_in_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_689_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33303\,
            in1 => \N__25034\,
            in2 => \N__26541\,
            in3 => \N__27926\,
            lcout => \c0.n8960\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30032\,
            in1 => \N__18439\,
            in2 => \_gnd_net_\,
            in3 => \N__19180\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i54_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22151\,
            in1 => \N__18420\,
            in2 => \_gnd_net_\,
            in3 => \N__19113\,
            lcout => data_in_field_53,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i131_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23714\,
            in1 => \N__26532\,
            in2 => \_gnd_net_\,
            in3 => \N__28752\,
            lcout => data_in_field_130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i13_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__19179\,
            in1 => \N__23508\,
            in2 => \N__18812\,
            in3 => \N__19112\,
            lcout => \c0.data_in_field_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9602_bdd_4_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32789\,
            in1 => \N__18849\,
            in2 => \N__18822\,
            in3 => \N__25613\,
            lcout => \c0.n9150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_586_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19206\,
            in2 => \_gnd_net_\,
            in3 => \N__18802\,
            lcout => \c0.n9019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_665_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18757\,
            in2 => \_gnd_net_\,
            in3 => \N__22208\,
            lcout => \c0.n8813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i59_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23944\,
            in2 => \N__28748\,
            in3 => \N__24040\,
            lcout => data_in_field_58,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_551_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26484\,
            in2 => \_gnd_net_\,
            in3 => \N__26813\,
            lcout => \c0.n8828\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i150_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19305\,
            in2 => \N__28747\,
            in3 => \N__19769\,
            lcout => data_in_field_149,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i139_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23943\,
            in1 => \N__26485\,
            in2 => \_gnd_net_\,
            in3 => \N__28567\,
            lcout => data_in_field_138,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i125_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29107\,
            in2 => \N__28745\,
            in3 => \N__24281\,
            lcout => data_in_field_124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i109_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21506\,
            in1 => \N__24887\,
            in2 => \_gnd_net_\,
            in3 => \N__28563\,
            lcout => data_in_field_108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i143_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19361\,
            in2 => \N__28746\,
            in3 => \N__26441\,
            lcout => data_in_field_142,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i65_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27843\,
            in1 => \N__25987\,
            in2 => \_gnd_net_\,
            in3 => \N__28577\,
            lcout => data_in_field_64,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7420_4_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001010000"
        )
    port map (
            in0 => \N__30269\,
            in1 => \N__30296\,
            in2 => \N__30360\,
            in3 => \N__30323\,
            lcout => n9091,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7421_4_lut_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010001010"
        )
    port map (
            in0 => \N__30297\,
            in1 => \N__30270\,
            in2 => \N__30327\,
            in3 => \N__30359\,
            lcout => OPEN,
            ltout => \n9092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7422_3_lut_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__19251\,
            in1 => \_gnd_net_\,
            in2 => \N__19245\,
            in3 => \N__30243\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__31086\,
            in1 => \N__27447\,
            in2 => \N__31032\,
            in3 => \N__30972\,
            lcout => \r_SM_Main_2_adj_1734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35364\,
            ce => 'H',
            sr => \N__19227\
        );

    \c0.i1_2_lut_3_lut_adj_699_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26380\,
            in1 => \N__25480\,
            in2 => \_gnd_net_\,
            in3 => \N__19214\,
            lcout => \c0.n8883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__23662\,
            in1 => \N__23401\,
            in2 => \_gnd_net_\,
            in3 => \N__20774\,
            lcout => \c0.n4897\,
            ltout => \c0.n4897_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3607_2_lut_3_lut_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__23402\,
            in1 => \_gnd_net_\,
            in2 => \N__19323\,
            in3 => \N__23663\,
            lcout => \c0.n5154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7744_3_lut_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__23661\,
            in1 => \N__23400\,
            in2 => \_gnd_net_\,
            in3 => \N__20775\,
            lcout => n4806,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i0_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25976\,
            in2 => \_gnd_net_\,
            in3 => \N__19320\,
            lcout => rand_data_0,
            ltout => OPEN,
            carryin => \bfn_6_27_0_\,
            carryout => n8155,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i1_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21018\,
            in2 => \_gnd_net_\,
            in3 => \N__19317\,
            lcout => rand_data_1,
            ltout => OPEN,
            carryin => n8155,
            carryout => n8156,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i2_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23706\,
            in2 => \_gnd_net_\,
            in3 => \N__19314\,
            lcout => rand_data_2,
            ltout => OPEN,
            carryin => n8156,
            carryout => n8157,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i3_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21144\,
            in2 => \_gnd_net_\,
            in3 => \N__19311\,
            lcout => rand_data_3,
            ltout => OPEN,
            carryin => n8157,
            carryout => n8158,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i4_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21179\,
            in2 => \_gnd_net_\,
            in3 => \N__19308\,
            lcout => rand_data_4,
            ltout => OPEN,
            carryin => n8158,
            carryout => n8159,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i5_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19272\,
            in2 => \_gnd_net_\,
            in3 => \N__19257\,
            lcout => rand_data_5,
            ltout => OPEN,
            carryin => n8159,
            carryout => n8160,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i6_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24629\,
            in2 => \_gnd_net_\,
            in3 => \N__19254\,
            lcout => rand_data_6,
            ltout => OPEN,
            carryin => n8160,
            carryout => n8161,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i7_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21063\,
            in2 => \_gnd_net_\,
            in3 => \N__19386\,
            lcout => rand_data_7,
            ltout => OPEN,
            carryin => n8161,
            carryout => n8162,
            clk => \N__35372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i8_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20903\,
            in2 => \_gnd_net_\,
            in3 => \N__19383\,
            lcout => rand_data_8,
            ltout => OPEN,
            carryin => \bfn_6_28_0_\,
            carryout => n8163,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i9_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21650\,
            in2 => \_gnd_net_\,
            in3 => \N__19380\,
            lcout => rand_data_9,
            ltout => OPEN,
            carryin => n8163,
            carryout => n8164,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i10_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23932\,
            in2 => \_gnd_net_\,
            in3 => \N__19377\,
            lcout => rand_data_10,
            ltout => OPEN,
            carryin => n8164,
            carryout => n8165,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i11_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26717\,
            in2 => \_gnd_net_\,
            in3 => \N__19374\,
            lcout => rand_data_11,
            ltout => OPEN,
            carryin => n8165,
            carryout => n8166,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i12_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29096\,
            in2 => \_gnd_net_\,
            in3 => \N__19371\,
            lcout => rand_data_12,
            ltout => OPEN,
            carryin => n8166,
            carryout => n8167,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i13_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21458\,
            in2 => \_gnd_net_\,
            in3 => \N__19368\,
            lcout => rand_data_13,
            ltout => OPEN,
            carryin => n8167,
            carryout => n8168,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i14_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19352\,
            in2 => \_gnd_net_\,
            in3 => \N__19329\,
            lcout => rand_data_14,
            ltout => OPEN,
            carryin => n8168,
            carryout => n8169,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i15_LC_6_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21576\,
            in2 => \_gnd_net_\,
            in3 => \N__19326\,
            lcout => rand_data_15,
            ltout => OPEN,
            carryin => n8169,
            carryout => n8170,
            clk => \N__35379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i16_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24106\,
            in2 => \_gnd_net_\,
            in3 => \N__19449\,
            lcout => rand_data_16,
            ltout => OPEN,
            carryin => \bfn_6_29_0_\,
            carryout => n8171,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i17_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19839\,
            in2 => \_gnd_net_\,
            in3 => \N__19446\,
            lcout => rand_data_17,
            ltout => OPEN,
            carryin => n8171,
            carryout => n8172,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i18_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26126\,
            in2 => \_gnd_net_\,
            in3 => \N__19443\,
            lcout => rand_data_18,
            ltout => OPEN,
            carryin => n8172,
            carryout => n8173,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i19_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19420\,
            in2 => \_gnd_net_\,
            in3 => \N__19404\,
            lcout => rand_data_19,
            ltout => OPEN,
            carryin => n8173,
            carryout => n8174,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i20_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24313\,
            in2 => \_gnd_net_\,
            in3 => \N__19401\,
            lcout => rand_data_20,
            ltout => OPEN,
            carryin => n8174,
            carryout => n8175,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i21_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19875\,
            in2 => \_gnd_net_\,
            in3 => \N__19398\,
            lcout => rand_data_21,
            ltout => OPEN,
            carryin => n8175,
            carryout => n8176,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i22_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20848\,
            in2 => \_gnd_net_\,
            in3 => \N__19395\,
            lcout => rand_data_22,
            ltout => OPEN,
            carryin => n8176,
            carryout => n8177,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i23_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19704\,
            in2 => \_gnd_net_\,
            in3 => \N__19392\,
            lcout => rand_data_23,
            ltout => OPEN,
            carryin => n8177,
            carryout => n8178,
            clk => \N__35386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i24_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20664\,
            in2 => \_gnd_net_\,
            in3 => \N__19389\,
            lcout => rand_data_24,
            ltout => OPEN,
            carryin => \bfn_6_30_0_\,
            carryout => n8179,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i25_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19588\,
            in2 => \_gnd_net_\,
            in3 => \N__19572\,
            lcout => rand_data_25,
            ltout => OPEN,
            carryin => n8179,
            carryout => n8180,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i26_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24070\,
            in2 => \_gnd_net_\,
            in3 => \N__19569\,
            lcout => rand_data_26,
            ltout => OPEN,
            carryin => n8180,
            carryout => n8181,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i27_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19539\,
            in2 => \_gnd_net_\,
            in3 => \N__19521\,
            lcout => rand_data_27,
            ltout => OPEN,
            carryin => n8181,
            carryout => n8182,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i28_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21486\,
            in2 => \_gnd_net_\,
            in3 => \N__19518\,
            lcout => rand_data_28,
            ltout => OPEN,
            carryin => n8182,
            carryout => n8183,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i29_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21258\,
            in2 => \_gnd_net_\,
            in3 => \N__19515\,
            lcout => rand_data_29,
            ltout => OPEN,
            carryin => n8183,
            carryout => n8184,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i30_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22284\,
            in2 => \_gnd_net_\,
            in3 => \N__19512\,
            lcout => rand_data_30,
            ltout => OPEN,
            carryin => n8184,
            carryout => n8185,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rand_data_422__i31_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19502\,
            in2 => \_gnd_net_\,
            in3 => \N__19509\,
            lcout => rand_data_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_8019_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__22326\,
            in1 => \N__27041\,
            in2 => \N__33014\,
            in3 => \N__32015\,
            lcout => OPEN,
            ltout => \c0.n9734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9734_bdd_4_lut_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__19479\,
            in1 => \N__32918\,
            in2 => \N__19452\,
            in3 => \N__27672\,
            lcout => \c0.n9234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_533_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19928\,
            in1 => \N__22058\,
            in2 => \_gnd_net_\,
            in3 => \N__19800\,
            lcout => \c0.n9013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i121_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22329\,
            in1 => \N__20920\,
            in2 => \_gnd_net_\,
            in3 => \N__29019\,
            lcout => data_in_field_120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i118_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19886\,
            in2 => \N__29065\,
            in3 => \N__19631\,
            lcout => data_in_field_117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i114_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19801\,
            in1 => \N__19852\,
            in2 => \_gnd_net_\,
            in3 => \N__29015\,
            lcout => data_in_field_113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1290_2_lut_3_lut_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19771\,
            in1 => \N__25214\,
            in2 => \_gnd_net_\,
            in3 => \N__25338\,
            lcout => \c0.n1893_adj_1635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i88_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19715\,
            in1 => \N__21929\,
            in2 => \_gnd_net_\,
            in3 => \N__29020\,
            lcout => data_in_field_87,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7905_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__19685\,
            in1 => \N__32052\,
            in2 => \N__33098\,
            in3 => \N__22022\,
            lcout => OPEN,
            ltout => \c0.n9596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9596_bdd_4_lut_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__22418\,
            in1 => \N__24398\,
            in2 => \N__19638\,
            in3 => \N__33028\,
            lcout => \c0.n9153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7900_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33029\,
            in1 => \N__19627\,
            in2 => \N__24559\,
            in3 => \N__32053\,
            lcout => OPEN,
            ltout => \c0.n9590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9590_bdd_4_lut_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__24188\,
            in1 => \N__21232\,
            in2 => \N__20055\,
            in3 => \N__33030\,
            lcout => OPEN,
            ltout => \c0.n9156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_7915_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__20052\,
            in1 => \N__31604\,
            in2 => \N__20046\,
            in3 => \N__31243\,
            lcout => OPEN,
            ltout => \c0.n9584_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9584_bdd_4_lut_LC_6_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__31605\,
            in1 => \N__21291\,
            in2 => \N__20043\,
            in3 => \N__20040\,
            lcout => OPEN,
            ltout => \c0.n9587_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i5_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32383\,
            in1 => \N__20028\,
            in2 => \N__20013\,
            in3 => \N__31606\,
            lcout => \c0.tx2.r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35406\,
            ce => \N__32229\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i86_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19983\,
            in1 => \N__29974\,
            in2 => \_gnd_net_\,
            in3 => \N__19994\,
            lcout => data_in_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i94_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19962\,
            in1 => \N__29979\,
            in2 => \_gnd_net_\,
            in3 => \N__19982\,
            lcout => data_in_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i102_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29977\,
            in1 => \N__19974\,
            in2 => \_gnd_net_\,
            in3 => \N__19961\,
            lcout => data_in_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i118_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19941\,
            in1 => \N__29972\,
            in2 => \_gnd_net_\,
            in3 => \N__19952\,
            lcout => data_in_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i126_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__29978\,
            in2 => \_gnd_net_\,
            in3 => \N__19940\,
            lcout => data_in_15_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i134_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20154\,
            in1 => \N__29973\,
            in2 => \_gnd_net_\,
            in3 => \N__20174\,
            lcout => data_in_16_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i142_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29971\,
            in1 => \N__20166\,
            in2 => \_gnd_net_\,
            in3 => \N__20153\,
            lcout => data_in_17_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i151_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20259\,
            in1 => \_gnd_net_\,
            in2 => \N__29988\,
            in3 => \N__20144\,
            lcout => data_in_18_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i146_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20115\,
            in1 => \N__29874\,
            in2 => \_gnd_net_\,
            in3 => \N__20126\,
            lcout => data_in_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i154_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20106\,
            in1 => \_gnd_net_\,
            in2 => \N__29989\,
            in3 => \N__20114\,
            lcout => data_in_19_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i162_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20190\,
            in1 => \N__29875\,
            in2 => \_gnd_net_\,
            in3 => \N__20105\,
            lcout => data_in_20_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__20282\,
            in1 => \N__28167\,
            in2 => \N__20097\,
            in3 => \N__20337\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i163_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29882\,
            in1 => \N__20093\,
            in2 => \_gnd_net_\,
            in3 => \N__23078\,
            lcout => data_in_20_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35322\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i92_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29926\,
            in1 => \N__20085\,
            in2 => \_gnd_net_\,
            in3 => \N__20066\,
            lcout => data_in_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__20270\,
            in1 => \N__28159\,
            in2 => \N__20289\,
            in3 => \N__20366\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i159_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20208\,
            in1 => \N__29927\,
            in2 => \_gnd_net_\,
            in3 => \N__20258\,
            lcout => data_in_19_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__20199\,
            in1 => \N__28157\,
            in2 => \N__20246\,
            in3 => \N__20336\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i152_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29925\,
            in1 => \N__20379\,
            in2 => \_gnd_net_\,
            in3 => \N__20219\,
            lcout => data_in_18_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i167_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29928\,
            in1 => \N__20430\,
            in2 => \_gnd_net_\,
            in3 => \N__20207\,
            lcout => data_in_20_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_32_i4_2_lut_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27551\,
            in2 => \_gnd_net_\,
            in3 => \N__25873\,
            lcout => n4_adj_1725,
            ltout => \n4_adj_1725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__20189\,
            in1 => \N__28158\,
            in2 => \N__20193\,
            in3 => \N__20365\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_506_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25926\,
            in2 => \_gnd_net_\,
            in3 => \N__27473\,
            lcout => n4044,
            ltout => \n4044_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__23058\,
            in1 => \N__20397\,
            in2 => \N__20178\,
            in3 => \N__28156\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__20335\,
            in1 => \N__20429\,
            in2 => \N__28166\,
            in3 => \N__23057\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__25823\,
            in1 => \N__28151\,
            in2 => \N__20414\,
            in3 => \N__20334\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i168_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20396\,
            in1 => \_gnd_net_\,
            in2 => \N__29987\,
            in3 => \N__20387\,
            lcout => data_in_20_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i160_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20388\,
            in1 => \N__29866\,
            in2 => \_gnd_net_\,
            in3 => \N__20378\,
            lcout => data_in_19_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__28152\,
            in1 => \N__25824\,
            in2 => \N__20352\,
            in3 => \N__20367\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25925\,
            in2 => \_gnd_net_\,
            in3 => \N__27474\,
            lcout => n4049,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_566_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26623\,
            in1 => \N__25128\,
            in2 => \N__27330\,
            in3 => \N__26500\,
            lcout => \c0.n28_adj_1619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7805_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__32870\,
            in1 => \N__31952\,
            in2 => \N__22057\,
            in3 => \N__22382\,
            lcout => \c0.n9476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_2056_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__23667\,
            in1 => \N__23524\,
            in2 => \N__20700\,
            in3 => \N__20789\,
            lcout => \c0.r_SM_Main_2_N_1483_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7965_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25303\,
            in1 => \N__32806\,
            in2 => \N__22935\,
            in3 => \N__31897\,
            lcout => \c0.n9668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_40_i1_3_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__20518\,
            in1 => \N__20676\,
            in2 => \N__23559\,
            in3 => \_gnd_net_\,
            lcout => n1903,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i130_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__20605\,
            in1 => \_gnd_net_\,
            in2 => \N__21045\,
            in3 => \N__28998\,
            lcout => data_in_field_129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_610_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20604\,
            in2 => \_gnd_net_\,
            in3 => \N__26060\,
            lcout => \c0.n8791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i145_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26061\,
            in1 => \N__25998\,
            in2 => \_gnd_net_\,
            in3 => \N__28999\,
            lcout => data_in_field_144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i41_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20519\,
            in1 => \N__29387\,
            in2 => \_gnd_net_\,
            in3 => \N__20562\,
            lcout => data_in_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_676_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20978\,
            in1 => \N__20993\,
            in2 => \N__20961\,
            in3 => \N__22818\,
            lcout => \c0.n19_adj_1665\,
            ltout => \c0.n19_adj_1665_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7763_2_lut_3_lut_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \N__20505\,
            in3 => \N__20501\,
            lcout => \c0.tx2_transmit_N_1444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5656_2_lut_3_lut_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__20502\,
            in1 => \_gnd_net_\,
            in2 => \N__20456\,
            in3 => \N__20436\,
            lcout => \c0.n7194\,
            ltout => \c0.n7194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_4_lut_adj_733_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001001110011"
        )
    port map (
            in0 => \N__23520\,
            in1 => \N__23659\,
            in2 => \N__20832\,
            in3 => \N__20829\,
            lcout => n4839,
            ltout => \n4839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state__i2_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__23660\,
            in1 => \N__23589\,
            in2 => \N__20793\,
            in3 => \N__20790\,
            lcout => \FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i66_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21040\,
            in1 => \N__20718\,
            in2 => \_gnd_net_\,
            in3 => \N__28873\,
            lcout => data_in_field_65,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i151_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24655\,
            in1 => \_gnd_net_\,
            in2 => \N__29008\,
            in3 => \N__25318\,
            lcout => data_in_field_150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i119_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__20880\,
            in1 => \_gnd_net_\,
            in2 => \N__24010\,
            in3 => \N__28869\,
            lcout => data_in_field_118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_425__i0_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20696\,
            in2 => \N__31971\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter2_0\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \c0.n8113\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i1_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32790\,
            in2 => \_gnd_net_\,
            in3 => \N__20685\,
            lcout => \c0.byte_transmit_counter2_1\,
            ltout => OPEN,
            carryin => \c0.n8113\,
            carryout => \c0.n8114\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i2_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31178\,
            in2 => \_gnd_net_\,
            in3 => \N__20682\,
            lcout => \c0.byte_transmit_counter2_2\,
            ltout => OPEN,
            carryin => \c0.n8114\,
            carryout => \c0.n8115\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i3_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31532\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => \c0.byte_transmit_counter2_3\,
            ltout => OPEN,
            carryin => \c0.n8115\,
            carryout => \c0.n8116\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i4_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32319\,
            in2 => \_gnd_net_\,
            in3 => \N__20997\,
            lcout => \c0.byte_transmit_counter2_4\,
            ltout => OPEN,
            carryin => \c0.n8116\,
            carryout => \c0.n8117\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i5_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20994\,
            in2 => \_gnd_net_\,
            in3 => \N__20982\,
            lcout => \c0.byte_transmit_counter2_5\,
            ltout => OPEN,
            carryin => \c0.n8117\,
            carryout => \c0.n8118\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i6_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20979\,
            in2 => \_gnd_net_\,
            in3 => \N__20967\,
            lcout => \c0.byte_transmit_counter2_6\,
            ltout => OPEN,
            carryin => \c0.n8118\,
            carryout => \c0.n8119\,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.byte_transmit_counter2_425__i7_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20960\,
            in2 => \_gnd_net_\,
            in3 => \N__20964\,
            lcout => \c0.byte_transmit_counter2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35365\,
            ce => \N__20946\,
            sr => \N__20934\
        );

    \c0.data_in_frame_0___i83_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26146\,
            in2 => \N__28743\,
            in3 => \N__32158\,
            lcout => data_in_field_82,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i89_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20922\,
            in1 => \N__28381\,
            in2 => \_gnd_net_\,
            in3 => \N__28558\,
            lcout => data_in_field_88,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i133_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21182\,
            in2 => \N__28742\,
            in3 => \N__33302\,
            lcout => data_in_field_132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i87_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20875\,
            in1 => \N__25118\,
            in2 => \_gnd_net_\,
            in3 => \N__28557\,
            lcout => data_in_field_86,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i96_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21584\,
            in1 => \_gnd_net_\,
            in2 => \N__28744\,
            in3 => \N__27703\,
            lcout => data_in_field_95,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i100_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21153\,
            in1 => \N__23824\,
            in2 => \_gnd_net_\,
            in3 => \N__28550\,
            lcout => data_in_field_99,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_577_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21125\,
            in1 => \N__23898\,
            in2 => \N__22128\,
            in3 => \N__23145\,
            lcout => \c0.n21_adj_1624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i91_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23951\,
            in1 => \N__32104\,
            in2 => \_gnd_net_\,
            in3 => \N__28559\,
            lcout => data_in_field_90,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i104_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21075\,
            in1 => \N__32538\,
            in2 => \_gnd_net_\,
            in3 => \N__28643\,
            lcout => data_in_field_103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i99_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23707\,
            in1 => \_gnd_net_\,
            in2 => \N__28851\,
            in3 => \N__31462\,
            lcout => data_in_field_98,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i101_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21180\,
            in1 => \N__24845\,
            in2 => \_gnd_net_\,
            in3 => \N__28642\,
            lcout => data_in_field_100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i69_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21181\,
            in2 => \N__28850\,
            in3 => \N__25511\,
            lcout => data_in_field_68,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i129_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25977\,
            in1 => \N__26179\,
            in2 => \_gnd_net_\,
            in3 => \N__28647\,
            lcout => data_in_field_128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i126_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21463\,
            in2 => \N__28848\,
            in3 => \N__24539\,
            lcout => data_in_field_125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i98_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21019\,
            in1 => \N__27763\,
            in2 => \_gnd_net_\,
            in3 => \N__28654\,
            lcout => data_in_field_97,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i144_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21577\,
            in2 => \N__28849\,
            in3 => \N__21537\,
            lcout => data_in_field_143,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35380\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_626_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26172\,
            lcout => \c0.n4288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i77_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21505\,
            in2 => \N__29007\,
            in3 => \N__25476\,
            lcout => data_in_field_76,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i62_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21465\,
            in1 => \N__21717\,
            in2 => \_gnd_net_\,
            in3 => \N__28863\,
            lcout => data_in_field_61,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7920_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__21431\,
            in1 => \N__32016\,
            in2 => \N__33024\,
            in3 => \N__21374\,
            lcout => OPEN,
            ltout => \c0.n9608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9608_bdd_4_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32946\,
            in1 => \N__22223\,
            in2 => \N__21330\,
            in3 => \N__21327\,
            lcout => \c0.n9147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i110_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21279\,
            in1 => \_gnd_net_\,
            in2 => \N__29005\,
            in3 => \N__21218\,
            lcout => data_in_field_109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i107_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24082\,
            in1 => \N__31414\,
            in2 => \_gnd_net_\,
            in3 => \N__28856\,
            lcout => data_in_field_106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i149_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21183\,
            in1 => \_gnd_net_\,
            in2 => \N__29006\,
            in3 => \N__32497\,
            lcout => data_in_field_148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_515_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24249\,
            lcout => \c0.n8942\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i58_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22056\,
            in1 => \_gnd_net_\,
            in2 => \N__21662\,
            in3 => \N__28868\,
            lcout => data_in_field_57,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_698_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24959\,
            in1 => \N__22023\,
            in2 => \_gnd_net_\,
            in3 => \N__22531\,
            lcout => \c0.n4390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_730_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21942\,
            in1 => \N__21892\,
            in2 => \N__21828\,
            in3 => \N__21675\,
            lcout => \c0.n4197\,
            ltout => \c0.n4197_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_545_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__21795\,
            in1 => \_gnd_net_\,
            in2 => \N__21753\,
            in3 => \_gnd_net_\,
            lcout => \c0.n8834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_619_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31407\,
            in2 => \_gnd_net_\,
            in3 => \N__21611\,
            lcout => \c0.n4399\,
            ltout => \c0.n4399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_541_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21718\,
            in1 => \N__25454\,
            in2 => \N__21693\,
            in3 => \N__21686\,
            lcout => \c0.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i122_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21654\,
            in1 => \N__21612\,
            in2 => \_gnd_net_\,
            in3 => \N__28867\,
            lcout => data_in_field_121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9572_bdd_4_lut_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__32945\,
            in1 => \N__22475\,
            in2 => \N__22809\,
            in3 => \N__22431\,
            lcout => \c0.n9165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_707_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22157\,
            in1 => \N__25512\,
            in2 => \N__22422\,
            in3 => \N__22383\,
            lcout => \c0.n8887\,
            ltout => \c0.n8887_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_705_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__32598\,
            in2 => \N__22332\,
            in3 => \N__22328\,
            lcout => \c0.n8893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i111_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27308\,
            in1 => \N__22294\,
            in2 => \_gnd_net_\,
            in3 => \N__29056\,
            lcout => data_in_field_110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_632_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22263\,
            in1 => \N__22238\,
            in2 => \_gnd_net_\,
            in3 => \N__32599\,
            lcout => OPEN,
            ltout => \c0.n4240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22164\,
            in1 => \N__26628\,
            in2 => \N__22227\,
            in3 => \N__22224\,
            lcout => \c0.n44_adj_1609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_553_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27307\,
            in2 => \_gnd_net_\,
            in3 => \N__24298\,
            lcout => \c0.n4553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_630_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22158\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25513\,
            lcout => \c0.n8964\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_50_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22116\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__31569\,
            in1 => \N__32348\,
            in2 => \_gnd_net_\,
            in3 => \N__31179\,
            lcout => \c0.n18_adj_1666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_652_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24003\,
            in1 => \N__22574\,
            in2 => \N__22737\,
            in3 => \N__22805\,
            lcout => \c0.n8810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1042_2_lut_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25218\,
            in2 => \_gnd_net_\,
            in3 => \N__25339\,
            lcout => \c0.n1645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7935_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__24450\,
            in1 => \N__32947\,
            in2 => \N__22736\,
            in3 => \N__32030\,
            lcout => OPEN,
            ltout => \c0.n9632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9632_bdd_4_lut_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32948\,
            in1 => \N__22686\,
            in2 => \N__22626\,
            in3 => \N__22623\,
            lcout => \c0.n9135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7925_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__32054\,
            in1 => \N__24011\,
            in2 => \N__22575\,
            in3 => \N__32848\,
            lcout => OPEN,
            ltout => \c0.n9620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9620_bdd_4_lut_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__32849\,
            in1 => \N__24604\,
            in2 => \N__22536\,
            in3 => \N__27327\,
            lcout => \c0.n9141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7930_LC_7_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__32055\,
            in1 => \N__32850\,
            in2 => \N__25138\,
            in3 => \N__22533\,
            lcout => OPEN,
            ltout => \c0.n9626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9626_bdd_4_lut_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32851\,
            in1 => \N__26404\,
            in2 => \N__22479\,
            in3 => \N__27081\,
            lcout => OPEN,
            ltout => \c0.n9138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_7940_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__31570\,
            in1 => \N__22911\,
            in2 => \N__22905\,
            in3 => \N__31192\,
            lcout => OPEN,
            ltout => \c0.n9614_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9614_bdd_4_lut_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__22902\,
            in1 => \N__22884\,
            in2 => \N__22878\,
            in3 => \N__31571\,
            lcout => OPEN,
            ltout => \c0.n9617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i6_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31572\,
            in1 => \N__31107\,
            in2 => \N__22875\,
            in3 => \N__32349\,
            lcout => \c0.tx2.r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35411\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i83_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22863\,
            in1 => \_gnd_net_\,
            in2 => \N__30034\,
            in3 => \N__23165\,
            lcout => data_in_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i91_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22854\,
            in1 => \N__30008\,
            in2 => \_gnd_net_\,
            in3 => \N__22862\,
            lcout => data_in_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i99_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22845\,
            in1 => \_gnd_net_\,
            in2 => \N__30035\,
            in3 => \N__22853\,
            lcout => data_in_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i107_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22836\,
            in1 => \N__30006\,
            in2 => \_gnd_net_\,
            in3 => \N__22844\,
            lcout => data_in_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i115_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22827\,
            in1 => \_gnd_net_\,
            in2 => \N__30033\,
            in3 => \N__22835\,
            lcout => data_in_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i123_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23115\,
            in1 => \N__30007\,
            in2 => \_gnd_net_\,
            in3 => \N__22826\,
            lcout => data_in_15_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i131_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30005\,
            in1 => \N__23097\,
            in2 => \_gnd_net_\,
            in3 => \N__23114\,
            lcout => data_in_16_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i147_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29990\,
            in1 => \N__23105\,
            in2 => \_gnd_net_\,
            in3 => \N__23067\,
            lcout => data_in_18_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i139_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23106\,
            in1 => \N__29992\,
            in2 => \_gnd_net_\,
            in3 => \N__23096\,
            lcout => data_in_17_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i155_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29991\,
            in1 => \N__23085\,
            in2 => \_gnd_net_\,
            in3 => \N__23066\,
            lcout => data_in_19_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5633_2_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27529\,
            in2 => \_gnd_net_\,
            in3 => \N__25863\,
            lcout => n7171,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9668_bdd_4_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__23043\,
            in1 => \N__26457\,
            in2 => \N__25809\,
            in3 => \N__32978\,
            lcout => \c0.n9671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_567_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23034\,
            in1 => \N__23016\,
            in2 => \N__26313\,
            in3 => \N__22995\,
            lcout => OPEN,
            ltout => \c0.n29_adj_1620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i159_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22950\,
            in1 => \N__23964\,
            in2 => \N__22938\,
            in3 => \N__23685\,
            lcout => \c0.data_in_frame_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35366\,
            ce => \N__29009\,
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_42_i1_3_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24089\,
            in1 => \N__26995\,
            in2 => \_gnd_net_\,
            in3 => \N__23551\,
            lcout => n1901,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i43_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26996\,
            in1 => \_gnd_net_\,
            in2 => \N__30030\,
            in3 => \N__23577\,
            lcout => data_in_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7655_2_lut_1_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \N__23669\,
            in1 => \N__23550\,
            in2 => \_gnd_net_\,
            in3 => \N__23609\,
            lcout => n9262,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i51_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29993\,
            in1 => \N__23190\,
            in2 => \_gnd_net_\,
            in3 => \N__23576\,
            lcout => data_in_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.mux_358_Mux_50_i1_3_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23575\,
            in1 => \N__26147\,
            in2 => \_gnd_net_\,
            in3 => \N__23549\,
            lcout => n1893,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i59_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23181\,
            in1 => \_gnd_net_\,
            in2 => \N__30031\,
            in3 => \N__23189\,
            lcout => data_in_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i67_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23154\,
            in1 => \N__29995\,
            in2 => \_gnd_net_\,
            in3 => \N__23180\,
            lcout => data_in_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i75_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29994\,
            in1 => \N__23153\,
            in2 => \_gnd_net_\,
            in3 => \N__23172\,
            lcout => data_in_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_724_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24888\,
            in1 => \N__26654\,
            in2 => \N__23787\,
            in3 => \N__23144\,
            lcout => \c0.n4562\,
            ltout => \c0.n4562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_582_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26004\,
            in1 => \N__26267\,
            in2 => \N__23118\,
            in3 => \N__26750\,
            lcout => \c0.n8837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_654_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32116\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26605\,
            lcout => OPEN,
            ltout => \c0.n4235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_549_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23877\,
            in1 => \N__27390\,
            in2 => \N__23862\,
            in3 => \N__23859\,
            lcout => \c0.n25_adj_1614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_618_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27932\,
            in2 => \_gnd_net_\,
            in3 => \N__26219\,
            lcout => \c0.n4365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_649_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27787\,
            in1 => \N__24184\,
            in2 => \N__23853\,
            in3 => \N__24291\,
            lcout => \c0.n4534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_725_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26655\,
            in1 => \N__23786\,
            in2 => \_gnd_net_\,
            in3 => \N__24889\,
            lcout => \c0.n8846\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i71_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27067\,
            in1 => \_gnd_net_\,
            in2 => \N__29053\,
            in3 => \N__24656\,
            lcout => data_in_field_70,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i67_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23721\,
            in1 => \N__31722\,
            in2 => \_gnd_net_\,
            in3 => \N__28957\,
            lcout => data_in_field_66,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i147_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23720\,
            in2 => \N__29052\,
            in3 => \N__26606\,
            lcout => data_in_field_146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_565_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28320\,
            in1 => \N__32447\,
            in2 => \N__24459\,
            in3 => \N__23894\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_721_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27066\,
            in1 => \N__27704\,
            in2 => \_gnd_net_\,
            in3 => \N__27411\,
            lcout => \c0.n8918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i75_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24090\,
            in1 => \N__31673\,
            in2 => \_gnd_net_\,
            in3 => \N__28961\,
            lcout => data_in_field_74,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_568_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24048\,
            in1 => \N__24012\,
            in2 => \N__23973\,
            in3 => \N__28388\,
            lcout => \c0.n27_adj_1621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i123_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27412\,
            in1 => \N__23952\,
            in2 => \_gnd_net_\,
            in3 => \N__28953\,
            lcout => data_in_field_122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_571_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33314\,
            in1 => \N__24579\,
            in2 => \_gnd_net_\,
            in3 => \N__27896\,
            lcout => \c0.n4473\,
            ltout => \c0.n4473_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_573_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27659\,
            in2 => \N__23901\,
            in3 => \N__26769\,
            lcout => \c0.n9010\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_597_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31460\,
            in2 => \_gnd_net_\,
            in3 => \N__24846\,
            lcout => \c0.n4511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_719_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31461\,
            in1 => \N__25804\,
            in2 => \N__24987\,
            in3 => \N__32513\,
            lcout => \c0.n4244\,
            ltout => \c0.n4244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_738_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28343\,
            in1 => \N__33247\,
            in2 => \N__23880\,
            in3 => \N__24224\,
            lcout => \c0.n8995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i103_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24580\,
            in1 => \N__24654\,
            in2 => \_gnd_net_\,
            in3 => \N__28924\,
            lcout => data_in_field_102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_716_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24549\,
            in1 => \N__24504\,
            in2 => \_gnd_net_\,
            in3 => \N__24984\,
            lcout => \c0.n18_adj_1618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_615_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25523\,
            in1 => \N__24449\,
            in2 => \_gnd_net_\,
            in3 => \N__24402\,
            lcout => \c0.n8912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_4_lut_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24372\,
            in1 => \N__31678\,
            in2 => \N__33257\,
            in3 => \N__28398\,
            lcout => \c0.n16_adj_1591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i117_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24331\,
            in2 => \N__29071\,
            in3 => \N__24242\,
            lcout => data_in_field_116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i85_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24332\,
            in1 => \N__24986\,
            in2 => \_gnd_net_\,
            in3 => \N__29046\,
            lcout => data_in_field_84,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7875_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__24292\,
            in1 => \N__24240\,
            in2 => \N__33204\,
            in3 => \N__31975\,
            lcout => \c0.n9560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_585_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24241\,
            in1 => \N__24225\,
            in2 => \N__24189\,
            in3 => \N__24985\,
            lcout => \c0.n16_adj_1629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i113_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24127\,
            in1 => \N__27033\,
            in2 => \_gnd_net_\,
            in3 => \N__29042\,
            lcout => data_in_field_112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_562_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24800\,
            in1 => \N__25059\,
            in2 => \N__25044\,
            in3 => \N__25023\,
            lcout => \c0.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7880_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__24980\,
            in1 => \N__31976\,
            in2 => \N__33135\,
            in3 => \N__24958\,
            lcout => \c0.n9566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_612_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26108\,
            in2 => \_gnd_net_\,
            in3 => \N__26186\,
            lcout => \c0.n8954\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9560_bdd_4_lut_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__24909\,
            in1 => \N__24902\,
            in2 => \N__33136\,
            in3 => \N__24856\,
            lcout => \c0.n9171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_587_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24813\,
            in1 => \N__24801\,
            in2 => \N__25079\,
            in3 => \N__24789\,
            lcout => \c0.n17_adj_1630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7975_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__32988\,
            in1 => \N__32509\,
            in2 => \N__24684\,
            in3 => \N__32037\,
            lcout => \c0.n9680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i157_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26030\,
            in1 => \N__24729\,
            in2 => \N__24720\,
            in3 => \N__24690\,
            lcout => \c0.data_in_frame_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35412\,
            ce => \N__29073\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__31343\,
            in1 => \N__32631\,
            in2 => \N__24675\,
            in3 => \N__31255\,
            lcout => \c0.n22_adj_1679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9566_bdd_4_lut_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__33023\,
            in1 => \N__25527\,
            in2 => \N__25482\,
            in3 => \N__25437\,
            lcout => OPEN,
            ltout => \c0.n9168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_7890_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__25428\,
            in1 => \N__31614\,
            in2 => \N__25419\,
            in3 => \N__31242\,
            lcout => \c0.n9554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9554_bdd_4_lut_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__31615\,
            in1 => \N__25416\,
            in2 => \N__25404\,
            in3 => \N__25383\,
            lcout => OPEN,
            ltout => \c0.n9557_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i4_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__25377\,
            in1 => \N__31616\,
            in2 => \N__25368\,
            in3 => \N__32382\,
            lcout => \c0.tx2.r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35417\,
            ce => \N__32277\,
            sr => \_gnd_net_\
        );

    \c0.rx.i7410_3_lut_4_lut_LC_9_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__27518\,
            in1 => \N__30792\,
            in2 => \N__27570\,
            in3 => \N__25947\,
            lcout => n5185,
            ltout => \n5185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_9_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000011000000"
        )
    port map (
            in0 => \N__25950\,
            in1 => \N__27519\,
            in2 => \N__25350\,
            in3 => \N__27568\,
            lcout => \r_Bit_Index_2_adj_1731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i7406_4_lut_LC_9_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30567\,
            in1 => \N__30724\,
            in2 => \N__30657\,
            in3 => \N__30791\,
            lcout => n9077,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_722_LC_9_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25347\,
            in1 => \N__25278\,
            in2 => \N__25224\,
            in3 => \N__25140\,
            lcout => \c0.n8915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_9_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000101000"
        )
    port map (
            in0 => \N__25935\,
            in1 => \N__25843\,
            in2 => \N__25906\,
            in3 => \N__25949\,
            lcout => \r_Bit_Index_1_adj_1732\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i635_2_lut_LC_9_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25842\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25895\,
            lcout => n2185,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_9_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__25948\,
            in1 => \N__25896\,
            in2 => \_gnd_net_\,
            in3 => \N__25934\,
            lcout => \r_Bit_Index_0_adj_1733\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.equal_29_i4_2_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27544\,
            in2 => \_gnd_net_\,
            in3 => \N__25875\,
            lcout => n4_adj_1724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_653_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25791\,
            in2 => \_gnd_net_\,
            in3 => \N__32514\,
            lcout => \c0.n8770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_3_lut_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32117\,
            in1 => \N__26612\,
            in2 => \_gnd_net_\,
            in3 => \N__25752\,
            lcout => \c0.n16_adj_1657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_657_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25711\,
            in1 => \N__25686\,
            in2 => \N__25673\,
            in3 => \N__25647\,
            lcout => OPEN,
            ltout => \c0.n22_adj_1655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_659_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25623\,
            in1 => \N__31731\,
            in2 => \N__25617\,
            in3 => \N__25614\,
            lcout => \c0.n24_adj_1658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i153_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28319\,
            in1 => \N__25572\,
            in2 => \N__25566\,
            in3 => \N__25542\,
            lcout => \c0.data_in_frame_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35381\,
            ce => \N__29047\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7855_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__26080\,
            in1 => \N__32884\,
            in2 => \N__32036\,
            in3 => \N__26229\,
            lcout => OPEN,
            ltout => \c0.n9536_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9536_bdd_4_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__32885\,
            in1 => \N__26223\,
            in2 => \N__26190\,
            in3 => \N__26187\,
            lcout => OPEN,
            ltout => \c0.n9539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__27195\,
            in1 => \N__31383\,
            in2 => \N__26154\,
            in3 => \N__31203\,
            lcout => \c0.n22_adj_1661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i115_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26096\,
            in1 => \N__26151\,
            in2 => \_gnd_net_\,
            in3 => \N__28962\,
            lcout => data_in_field_114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7820_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__27410\,
            in1 => \N__26095\,
            in2 => \N__33090\,
            in3 => \N__31993\,
            lcout => \c0.n9494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_584_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26079\,
            in2 => \_gnd_net_\,
            in3 => \N__26501\,
            lcout => \c0.n8971\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_581_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26592\,
            in2 => \_gnd_net_\,
            in3 => \N__32160\,
            lcout => \c0.n6_adj_1628\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i97_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27647\,
            in1 => \N__25997\,
            in2 => \_gnd_net_\,
            in3 => \N__28966\,
            lcout => data_in_field_96,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_595_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31712\,
            in2 => \_gnd_net_\,
            in3 => \N__27646\,
            lcout => OPEN,
            ltout => \c0.n8840_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_599_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26554\,
            in1 => \N__26783\,
            in2 => \N__26772\,
            in3 => \N__26768\,
            lcout => \c0.n4309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i124_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26738\,
            in2 => \N__29054\,
            in3 => \N__26659\,
            lcout => data_in_field_123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7989_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__26591\,
            in1 => \N__33018\,
            in2 => \N__26238\,
            in3 => \N__31977\,
            lcout => OPEN,
            ltout => \c0.n9698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9698_bdd_4_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33019\,
            in1 => \N__26555\,
            in2 => \N__26508\,
            in3 => \N__26505\,
            lcout => OPEN,
            ltout => \c0.n9701_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31379\,
            in1 => \N__27009\,
            in2 => \N__26466\,
            in3 => \N__31233\,
            lcout => \c0.n22_adj_1681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_713_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26463\,
            in1 => \N__32171\,
            in2 => \N__26408\,
            in3 => \N__26346\,
            lcout => \c0.n8819\,
            ltout => \c0.n8819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_624_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26303\,
            in1 => \N__26292\,
            in2 => \N__26274\,
            in3 => \N__26271\,
            lcout => OPEN,
            ltout => \c0.n21_adj_1644_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i155_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__27489\,
            in1 => \_gnd_net_\,
            in2 => \N__26256\,
            in3 => \N__26253\,
            lcout => \c0.data_in_frame_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35396\,
            ce => \N__29048\,
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_547_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27372\,
            in1 => \N__32554\,
            in2 => \N__27345\,
            in3 => \N__27329\,
            lcout => \c0.n26_adj_1613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_548_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27276\,
            in1 => \N__27162\,
            in2 => \N__27270\,
            in3 => \N__27240\,
            lcout => OPEN,
            ltout => \c0.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i161_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27222\,
            in1 => \N__27213\,
            in2 => \N__27207\,
            in3 => \N__27204\,
            lcout => \c0.data_in_frame_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => \N__29030\,
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_535_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27176\,
            in1 => \N__27161\,
            in2 => \N__27147\,
            in3 => \N__27123\,
            lcout => OPEN,
            ltout => \c0.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i163_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__27102\,
            in1 => \N__27077\,
            in2 => \N__27048\,
            in3 => \N__27034\,
            lcout => \c0.data_in_frame_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35402\,
            ce => \N__29030\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i35_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29842\,
            in1 => \N__26959\,
            in2 => \_gnd_net_\,
            in3 => \N__27003\,
            lcout => data_in_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.i6_1_lut_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26942\,
            lcout => \c0.tx2.n4880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_620_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27614\,
            in1 => \N__26853\,
            in2 => \N__26838\,
            in3 => \N__26823\,
            lcout => \c0.n20_adj_1642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__30450\,
            in1 => \N__31016\,
            in2 => \N__30530\,
            in3 => \N__30489\,
            lcout => OPEN,
            ltout => \n12_adj_1753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7695_4_lut_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30965\,
            in1 => \N__31074\,
            in2 => \N__27480\,
            in3 => \N__30411\,
            lcout => n9246,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__31073\,
            in1 => \N__27440\,
            in2 => \N__31021\,
            in3 => \N__30964\,
            lcout => \r_SM_Main_2_N_1537_2\,
            ltout => \r_SM_Main_2_N_1537_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__30641\,
            in1 => \N__30721\,
            in2 => \N__27477\,
            in3 => \N__30786\,
            lcout => \c0.rx.n4090\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5849_3_lut_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__30488\,
            in1 => \N__30410\,
            in2 => \_gnd_net_\,
            in3 => \N__30449\,
            lcout => \c0.rx.n7393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i7_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__31012\,
            in1 => \N__30909\,
            in2 => \N__30876\,
            in3 => \N__30978\,
            lcout => \r_Clock_Count_7_adj_1727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_590_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27720\,
            in2 => \_gnd_net_\,
            in3 => \N__27425\,
            lcout => \c0.n4537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i6_4_lut_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__30491\,
            in1 => \N__30451\,
            in2 => \N__27594\,
            in3 => \N__30963\,
            lcout => \c0.rx.r_SM_Main_2_N_1543_0\,
            ltout => \c0.rx.r_SM_Main_2_N_1543_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_2_lut_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__28163\,
            in1 => \_gnd_net_\,
            in2 => \N__27375\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n6_adj_1751_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__30714\,
            in1 => \N__30658\,
            in2 => \N__27798\,
            in3 => \N__30783\,
            lcout => n30,
            ltout => \n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_10_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__30504\,
            in1 => \N__30523\,
            in2 => \N__27795\,
            in3 => \N__30873\,
            lcout => \r_Clock_Count_0_adj_1730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_643_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27786\,
            in1 => \N__27727\,
            in2 => \_gnd_net_\,
            in3 => \N__27671\,
            lcout => \c0.n4296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i5_4_lut_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__31072\,
            in1 => \N__30522\,
            in2 => \N__31022\,
            in3 => \N__30412\,
            lcout => \c0.rx.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_I_0_1_lut_LC_10_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34112\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_10_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101010101"
        )
    port map (
            in0 => \N__30720\,
            in1 => \N__27569\,
            in2 => \N__27535\,
            in3 => \N__30569\,
            lcout => OPEN,
            ltout => \n7415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_10_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__30659\,
            in1 => \N__30784\,
            in2 => \N__27495\,
            in3 => \N__28173\,
            lcout => \r_SM_Main_0_adj_1736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i7714_2_lut_LC_10_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30719\,
            in2 => \_gnd_net_\,
            in3 => \N__30568\,
            lcout => OPEN,
            ltout => \n9301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_10_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000010101"
        )
    port map (
            in0 => \N__30660\,
            in1 => \N__30785\,
            in2 => \N__27492\,
            in3 => \N__28089\,
            lcout => \r_SM_Main_1_adj_1735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_10_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__28098\,
            in1 => \_gnd_net_\,
            in2 => \N__30728\,
            in3 => \N__28164\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i7683_3_lut_LC_10_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__28165\,
            in1 => \N__28097\,
            in2 => \_gnd_net_\,
            in3 => \N__30715\,
            lcout => n9300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7790_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__32044\,
            in1 => \N__28083\,
            in2 => \N__33150\,
            in3 => \N__28053\,
            lcout => OPEN,
            ltout => \c0.n9446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9446_bdd_4_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__28023\,
            in1 => \N__27993\,
            in2 => \N__27957\,
            in3 => \N__33095\,
            lcout => OPEN,
            ltout => \c0.n9449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9728_bdd_4_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__27954\,
            in1 => \N__27804\,
            in2 => \N__27939\,
            in3 => \N__31583\,
            lcout => \c0.n9731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_8024_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__27931\,
            in1 => \N__28395\,
            in2 => \N__32987\,
            in3 => \N__31967\,
            lcout => OPEN,
            ltout => \c0.n9740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9740_bdd_4_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__27897\,
            in1 => \N__32889\,
            in2 => \N__27858\,
            in3 => \N__27855\,
            lcout => OPEN,
            ltout => \c0.n9231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__27822\,
            in1 => \N__31551\,
            in2 => \N__27807\,
            in3 => \N__31193\,
            lcout => \c0.n9728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i0_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__31552\,
            in1 => \N__32344\,
            in2 => \N__30072\,
            in3 => \N__30060\,
            lcout => \c0.tx2.r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35390\,
            ce => \N__32271\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i145_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29841\,
            in1 => \N__29126\,
            in2 => \_gnd_net_\,
            in3 => \N__29157\,
            lcout => data_in_18_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0___i141_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29115\,
            in1 => \N__33234\,
            in2 => \_gnd_net_\,
            in3 => \N__28967\,
            lcout => data_in_field_140,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_537_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31674\,
            in2 => \_gnd_net_\,
            in3 => \N__28396\,
            lcout => \c0.n4292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_646_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32164\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33233\,
            lcout => \c0.n8957\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_688_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28301\,
            in2 => \_gnd_net_\,
            in3 => \N__28248\,
            lcout => \c0.n8871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i0_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28191\,
            in2 => \_gnd_net_\,
            in3 => \N__28185\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_11_27_0_\,
            carryout => n8130,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i1_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28182\,
            in2 => \_gnd_net_\,
            in3 => \N__28176\,
            lcout => n25_adj_1722,
            ltout => OPEN,
            carryin => n8130,
            carryout => n8131,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i2_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30153\,
            in2 => \_gnd_net_\,
            in3 => \N__30147\,
            lcout => n24,
            ltout => OPEN,
            carryin => n8131,
            carryout => n8132,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i3_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30144\,
            in2 => \_gnd_net_\,
            in3 => \N__30138\,
            lcout => n23,
            ltout => OPEN,
            carryin => n8132,
            carryout => n8133,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i4_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30135\,
            in2 => \_gnd_net_\,
            in3 => \N__30129\,
            lcout => n22,
            ltout => OPEN,
            carryin => n8133,
            carryout => n8134,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i5_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30126\,
            in2 => \_gnd_net_\,
            in3 => \N__30120\,
            lcout => n21,
            ltout => OPEN,
            carryin => n8134,
            carryout => n8135,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i6_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30117\,
            in2 => \_gnd_net_\,
            in3 => \N__30111\,
            lcout => n20,
            ltout => OPEN,
            carryin => n8135,
            carryout => n8136,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i7_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30108\,
            in2 => \_gnd_net_\,
            in3 => \N__30102\,
            lcout => n19,
            ltout => OPEN,
            carryin => n8136,
            carryout => n8137,
            clk => \N__35403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i8_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30099\,
            in2 => \_gnd_net_\,
            in3 => \N__30093\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_11_28_0_\,
            carryout => n8138,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i9_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30090\,
            in2 => \_gnd_net_\,
            in3 => \N__30084\,
            lcout => n17,
            ltout => OPEN,
            carryin => n8138,
            carryout => n8139,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i10_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30081\,
            in2 => \_gnd_net_\,
            in3 => \N__30075\,
            lcout => n16,
            ltout => OPEN,
            carryin => n8139,
            carryout => n8140,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i11_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30225\,
            in2 => \_gnd_net_\,
            in3 => \N__30219\,
            lcout => n15,
            ltout => OPEN,
            carryin => n8140,
            carryout => n8141,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i12_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30216\,
            in2 => \_gnd_net_\,
            in3 => \N__30210\,
            lcout => n14,
            ltout => OPEN,
            carryin => n8141,
            carryout => n8142,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i13_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30207\,
            in2 => \_gnd_net_\,
            in3 => \N__30201\,
            lcout => n13,
            ltout => OPEN,
            carryin => n8142,
            carryout => n8143,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i14_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30198\,
            in2 => \_gnd_net_\,
            in3 => \N__30192\,
            lcout => n12,
            ltout => OPEN,
            carryin => n8143,
            carryout => n8144,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i15_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30189\,
            in2 => \_gnd_net_\,
            in3 => \N__30183\,
            lcout => n11,
            ltout => OPEN,
            carryin => n8144,
            carryout => n8145,
            clk => \N__35409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i16_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30180\,
            in2 => \_gnd_net_\,
            in3 => \N__30174\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_11_29_0_\,
            carryout => n8146,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i17_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30171\,
            in2 => \_gnd_net_\,
            in3 => \N__30165\,
            lcout => n9,
            ltout => OPEN,
            carryin => n8146,
            carryout => n8147,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i18_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30162\,
            in2 => \_gnd_net_\,
            in3 => \N__30156\,
            lcout => n8,
            ltout => OPEN,
            carryin => n8147,
            carryout => n8148,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i19_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30378\,
            in2 => \_gnd_net_\,
            in3 => \N__30372\,
            lcout => n7,
            ltout => OPEN,
            carryin => n8148,
            carryout => n8149,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i20_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30369\,
            in2 => \_gnd_net_\,
            in3 => \N__30363\,
            lcout => n6,
            ltout => OPEN,
            carryin => n8149,
            carryout => n8150,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i21_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30341\,
            in2 => \_gnd_net_\,
            in3 => \N__30330\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n8150,
            carryout => n8151,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i22_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30311\,
            in2 => \_gnd_net_\,
            in3 => \N__30300\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n8151,
            carryout => n8152,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i23_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30284\,
            in2 => \_gnd_net_\,
            in3 => \N__30273\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n8152,
            carryout => n8153,
            clk => \N__35414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i24_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30260\,
            in2 => \_gnd_net_\,
            in3 => \N__30249\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_11_30_0_\,
            carryout => n8154,
            clk => \N__35419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_423__i25_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30236\,
            in2 => \_gnd_net_\,
            in3 => \N__30246\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i6_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__30913\,
            in1 => \N__31076\,
            in2 => \N__31044\,
            in3 => \N__30869\,
            lcout => \r_Clock_Count_6_adj_1728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i2_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__30867\,
            in1 => \N__30911\,
            in2 => \N__30426\,
            in3 => \N__30453\,
            lcout => \r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i1_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__30910\,
            in1 => \N__30868\,
            in2 => \N__30495\,
            in3 => \N__30465\,
            lcout => \r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i48_4_lut_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000101"
        )
    port map (
            in0 => \N__30787\,
            in1 => \N__30738\,
            in2 => \N__30732\,
            in3 => \N__30537\,
            lcout => n44,
            ltout => \n44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i3_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__30912\,
            in1 => \N__30387\,
            in2 => \N__30663\,
            in3 => \N__30414\,
            lcout => \r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7646_2_lut_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30563\,
            lcout => n9245,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_2_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30531\,
            in3 => \N__30498\,
            lcout => n226,
            ltout => OPEN,
            carryin => \bfn_11_31_0_\,
            carryout => \c0.rx.n8098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_3_lut_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30490\,
            in2 => \_gnd_net_\,
            in3 => \N__30456\,
            lcout => n225,
            ltout => OPEN,
            carryin => \c0.rx.n8098\,
            carryout => \c0.rx.n8099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_4_lut_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30452\,
            in2 => \_gnd_net_\,
            in3 => \N__30417\,
            lcout => n224,
            ltout => OPEN,
            carryin => \c0.rx.n8099\,
            carryout => \c0.rx.n8100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_5_lut_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30413\,
            in2 => \_gnd_net_\,
            in3 => \N__30381\,
            lcout => n223,
            ltout => OPEN,
            carryin => \c0.rx.n8100\,
            carryout => \c0.rx.n8101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_6_lut_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30837\,
            in2 => \_gnd_net_\,
            in3 => \N__31092\,
            lcout => n222,
            ltout => OPEN,
            carryin => \c0.rx.n8101\,
            carryout => \c0.rx.n8102\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_7_lut_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30930\,
            in2 => \_gnd_net_\,
            in3 => \N__31089\,
            lcout => n221,
            ltout => OPEN,
            carryin => \c0.rx.n8102\,
            carryout => \c0.rx.n8103\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_8_lut_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31075\,
            in2 => \_gnd_net_\,
            in3 => \N__31035\,
            lcout => n220,
            ltout => OPEN,
            carryin => \c0.rx.n8103\,
            carryout => \c0.rx.n8104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.add_62_9_lut_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31020\,
            in2 => \_gnd_net_\,
            in3 => \N__30981\,
            lcout => n219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_505_LC_11_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30928\,
            in2 => \_gnd_net_\,
            in3 => \N__30835\,
            lcout => n4084,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i5_LC_11_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__30929\,
            in1 => \N__30915\,
            in2 => \N__30942\,
            in3 => \N__30875\,
            lcout => \r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i4_LC_11_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__30836\,
            in1 => \N__30914\,
            in2 => \N__30885\,
            in3 => \N__30874\,
            lcout => \r_Clock_Count_4_adj_1729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9488_bdd_4_lut_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__30822\,
            in1 => \N__31476\,
            in2 => \N__30807\,
            in3 => \N__31585\,
            lcout => OPEN,
            ltout => \c0.n9491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_i2_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31586\,
            in1 => \N__32403\,
            in2 => \N__32391\,
            in3 => \N__32381\,
            lcout => \c0.tx2.r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35404\,
            ce => \N__32272\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0__bdd_4_lut_7825_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__32159\,
            in1 => \N__33091\,
            in2 => \N__32120\,
            in3 => \N__32043\,
            lcout => \c0.n9500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9500_bdd_4_lut_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__33097\,
            in1 => \N__31732\,
            in2 => \N__31686\,
            in3 => \N__31638\,
            lcout => OPEN,
            ltout => \c0.n9198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_2__bdd_4_lut_7835_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__31389\,
            in1 => \N__31584\,
            in2 => \N__31479\,
            in3 => \N__31232\,
            lcout => \c0.n9488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9494_bdd_4_lut_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000010"
        )
    port map (
            in0 => \N__31470\,
            in1 => \N__31431\,
            in2 => \N__33210\,
            in3 => \N__31415\,
            lcout => \c0.n9201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__31360\,
            in1 => \N__31296\,
            in2 => \N__31281\,
            in3 => \N__31259\,
            lcout => \c0.n22_adj_1677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34031\,
            in2 => \_gnd_net_\,
            in3 => \N__33985\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_3_lut_4_lut_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__33986\,
            in1 => \N__35638\,
            in2 => \N__34440\,
            in3 => \N__34032\,
            lcout => n5062,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i3_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__34351\,
            in1 => \N__33673\,
            in2 => \N__35814\,
            in3 => \N__33420\,
            lcout => \c0.byte_transmit_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35405\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_2_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33849\,
            in2 => \N__33836\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_out_6_7_N_965_0\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \c0.n8083\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_3_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33896\,
            in2 => \_gnd_net_\,
            in3 => \N__32424\,
            lcout => \c0.data_out_6_7_N_965_1\,
            ltout => OPEN,
            carryin => \c0.n8083\,
            carryout => \c0.n8084\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_4_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33700\,
            in2 => \_gnd_net_\,
            in3 => \N__32421\,
            lcout => \c0.data_out_6_7_N_965_2\,
            ltout => OPEN,
            carryin => \c0.n8084\,
            carryout => \c0.n8085\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_5_lut_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33660\,
            in2 => \_gnd_net_\,
            in3 => \N__32418\,
            lcout => \c0.data_out_6_7_N_965_3\,
            ltout => OPEN,
            carryin => \c0.n8085\,
            carryout => \c0.n8086\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_6_lut_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33758\,
            in2 => \_gnd_net_\,
            in3 => \N__32415\,
            lcout => \c0.data_out_6_7_N_965_4\,
            ltout => OPEN,
            carryin => \c0.n8086\,
            carryout => \c0.n8087\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_7_lut_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33494\,
            in2 => \_gnd_net_\,
            in3 => \N__32412\,
            lcout => \data_out_6_7_N_965_5\,
            ltout => OPEN,
            carryin => \c0.n8087\,
            carryout => \c0.n8088\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_8_lut_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33443\,
            in2 => \_gnd_net_\,
            in3 => \N__32409\,
            lcout => \c0.data_out_6_7_N_965_6\,
            ltout => OPEN,
            carryin => \c0.n8088\,
            carryout => \c0.n8089\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_2248_9_lut_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33431\,
            in2 => \_gnd_net_\,
            in3 => \N__32406\,
            lcout => \c0.data_out_6_7_N_965_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_740_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__33780\,
            in1 => \N__33675\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n11\,
            ltout => \c0.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_691_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__33821\,
            in1 => \N__33727\,
            in2 => \N__32619\,
            in3 => \N__33910\,
            lcout => \tx_data_0_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_692_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__33911\,
            in1 => \N__33375\,
            in2 => \N__33842\,
            in3 => \N__33861\,
            lcout => OPEN,
            ltout => \tx_data_3_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34207\,
            in1 => \_gnd_net_\,
            in2 => \N__32616\,
            in3 => \N__33632\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33779\,
            in1 => \N__33674\,
            in2 => \_gnd_net_\,
            in3 => \N__33820\,
            lcout => \c0.n45_adj_1656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32613\,
            in1 => \N__34218\,
            in2 => \_gnd_net_\,
            in3 => \N__34079\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7754_4_lut_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__33918\,
            in1 => \N__33724\,
            in2 => \N__33379\,
            in3 => \N__33837\,
            lcout => \tx_data_7_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_564_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32607\,
            in1 => \N__32556\,
            in2 => \_gnd_net_\,
            in3 => \N__32507\,
            lcout => \c0.n8986\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_696_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__33917\,
            in1 => \N__32430\,
            in2 => \_gnd_net_\,
            in3 => \N__33725\,
            lcout => \tx_data_6_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_4_lut_4_lut_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001010"
        )
    port map (
            in0 => \N__33919\,
            in1 => \N__33726\,
            in2 => \N__33380\,
            in3 => \N__33838\,
            lcout => OPEN,
            ltout => \tx_data_5_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34219\,
            in2 => \N__33384\,
            in3 => \N__33584\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__33843\,
            in1 => \N__33920\,
            in2 => \N__33735\,
            in3 => \N__33381\,
            lcout => OPEN,
            ltout => \tx_data_2_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__33330\,
            in1 => \_gnd_net_\,
            in2 => \N__33351\,
            in3 => \N__34220\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33348\,
            in1 => \N__34221\,
            in2 => \_gnd_net_\,
            in3 => \N__33339\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000010000"
        )
    port map (
            in0 => \N__34003\,
            in1 => \N__35631\,
            in2 => \N__34568\,
            in3 => \N__34439\,
            lcout => OPEN,
            ltout => \n8705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__35632\,
            in1 => \_gnd_net_\,
            in2 => \N__33342\,
            in3 => \N__34044\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_7994_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__33338\,
            in1 => \N__33329\,
            in2 => \N__33987\,
            in3 => \N__35630\,
            lcout => n9452,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__34034\,
            in1 => \N__34004\,
            in2 => \_gnd_net_\,
            in3 => \N__34043\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n9680_bdd_4_lut_LC_13_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__33321\,
            in1 => \N__33273\,
            in2 => \N__33261\,
            in3 => \N__33096\,
            lcout => \c0.n9683\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_3_lut_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__34983\,
            in1 => \N__35850\,
            in2 => \_gnd_net_\,
            in3 => \N__34917\,
            lcout => OPEN,
            ltout => \c0.n17_adj_1663_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_671_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34125\,
            in1 => \N__34230\,
            in2 => \N__33453\,
            in3 => \N__33927\,
            lcout => \c0.n123\,
            ltout => \c0.n123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i4_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__35785\,
            in1 => \N__33770\,
            in2 => \N__33450\,
            in3 => \N__33543\,
            lcout => \c0.byte_transmit_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i2_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__33473\,
            in1 => \N__33719\,
            in2 => \N__35813\,
            in3 => \N__33408\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i6_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__34348\,
            in1 => \N__35786\,
            in2 => \N__33447\,
            in3 => \N__33555\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i7_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__33432\,
            in1 => \N__34349\,
            in2 => \N__35812\,
            in3 => \N__33531\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.UART_TRANSMITTER_state__i1_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__34350\,
            in1 => \N__35784\,
            in2 => \_gnd_net_\,
            in3 => \N__34283\,
            lcout => \UART_TRANSMITTER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__33419\,
            in1 => \N__33482\,
            in2 => \N__33396\,
            in3 => \N__33407\,
            lcout => \c0.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i0_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__33469\,
            in1 => \N__33395\,
            in2 => \N__35815\,
            in3 => \N__33835\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_672_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33506\,
            in2 => \_gnd_net_\,
            in3 => \N__33554\,
            lcout => OPEN,
            ltout => \c0.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_673_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33542\,
            in1 => \N__33530\,
            in2 => \N__33519\,
            in3 => \N__33516\,
            lcout => \c0.n7814\,
            ltout => \c0.n7814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_674_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__34347\,
            in1 => \_gnd_net_\,
            in2 => \N__33510\,
            in3 => \_gnd_net_\,
            lcout => n7204,
            ltout => \n7204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i5_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__33507\,
            in1 => \N__35817\,
            in2 => \N__33498\,
            in3 => \N__33495\,
            lcout => byte_transmit_counter_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_1995_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34547\,
            in1 => \N__34284\,
            in2 => \N__35827\,
            in3 => \N__34158\,
            lcout => \c0.tx_transmit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter__i1_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__33483\,
            in1 => \N__35816\,
            in2 => \N__33474\,
            in3 => \N__33913\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7750_3_lut_4_lut_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33677\,
            in1 => \N__33723\,
            in2 => \N__33921\,
            in3 => \N__33777\,
            lcout => \tx_data_1_N_keep\,
            ltout => \tx_data_1_N_keep_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34195\,
            in2 => \N__33456\,
            in3 => \N__33599\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35421\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_663_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__33676\,
            in1 => \N__33823\,
            in2 => \_gnd_net_\,
            in3 => \N__33776\,
            lcout => OPEN,
            ltout => \c0.n7779_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_693_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__33912\,
            in1 => \N__33639\,
            in2 => \N__33864\,
            in3 => \N__33860\,
            lcout => \tx_data_4_N_keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_737_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34167\,
            in2 => \_gnd_net_\,
            in3 => \N__34153\,
            lcout => \c0.data_out_6__7__N_973\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7693_2_lut_3_lut_4_lut_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33822\,
            in1 => \N__33778\,
            in2 => \N__33731\,
            in3 => \N__33678\,
            lcout => \c0.n9291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33984\,
            in1 => \N__33633\,
            in2 => \N__33612\,
            in3 => \N__35645\,
            lcout => n9710,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33618\,
            in1 => \N__34196\,
            in2 => \_gnd_net_\,
            in3 => \N__33611\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35421\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n9710_bdd_4_lut_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__33973\,
            in1 => \N__33600\,
            in2 => \N__33585\,
            in3 => \N__33570\,
            lcout => OPEN,
            ltout => \n9713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i591325_i1_3_lut_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34033\,
            in1 => \_gnd_net_\,
            in2 => \N__33564\,
            in3 => \N__34065\,
            lcout => OPEN,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34501\,
            in2 => \N__33561\,
            in3 => \N__34427\,
            lcout => OPEN,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34097\,
            in2 => \N__33558\,
            in3 => \N__35538\,
            lcout => tx_o_adj_1726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n9452_bdd_4_lut_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__34086\,
            in1 => \N__34052\,
            in2 => \N__34080\,
            in3 => \N__33972\,
            lcout => n9455,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34053\,
            in1 => \N__34200\,
            in2 => \_gnd_net_\,
            in3 => \N__34059\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7402_4_lut_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__35536\,
            in1 => \N__35745\,
            in2 => \N__34500\,
            in3 => \N__34423\,
            lcout => n9073,
            ltout => \n9073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000010"
        )
    port map (
            in0 => \N__34035\,
            in1 => \N__34008\,
            in2 => \N__33990\,
            in3 => \N__33980\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35537\,
            in1 => \N__34658\,
            in2 => \_gnd_net_\,
            in3 => \N__34638\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Done_44_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111101100"
        )
    port map (
            in0 => \N__34512\,
            in1 => \N__34359\,
            in2 => \N__33936\,
            in3 => \N__35553\,
            lcout => n3892,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_669_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34719\,
            in1 => \N__34892\,
            in2 => \N__34854\,
            in3 => \N__34679\,
            lcout => \c0.n18_adj_1662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5731_2_lut_3_lut_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__34680\,
            in1 => \N__34339\,
            in2 => \_gnd_net_\,
            in3 => \N__34279\,
            lcout => \c0.n20_adj_1652\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5736_2_lut_3_lut_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__34282\,
            in1 => \_gnd_net_\,
            in2 => \N__34353\,
            in3 => \N__34893\,
            lcout => \c0.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5730_2_lut_3_lut_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__34698\,
            in1 => \N__34338\,
            in2 => \_gnd_net_\,
            in3 => \N__34278\,
            lcout => \c0.n21_adj_1653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5733_2_lut_3_lut_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__34281\,
            in1 => \_gnd_net_\,
            in2 => \N__34352\,
            in3 => \N__34958\,
            lcout => \c0.n18_adj_1650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_670_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34697\,
            in1 => \N__34937\,
            in2 => \N__34959\,
            in3 => \N__34874\,
            lcout => \c0.n19_adj_1664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5732_2_lut_3_lut_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__34982\,
            in1 => \N__34340\,
            in2 => \_gnd_net_\,
            in3 => \N__34280\,
            lcout => \c0.n19_adj_1651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5667_2_lut_3_lut_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__34272\,
            in1 => \N__34718\,
            in2 => \_gnd_net_\,
            in3 => \N__34332\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_675_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__34543\,
            in1 => \N__34271\,
            in2 => \_gnd_net_\,
            in3 => \N__34157\,
            lcout => \c0.n900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5734_2_lut_3_lut_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__34273\,
            in1 => \N__34938\,
            in2 => \_gnd_net_\,
            in3 => \N__34333\,
            lcout => \c0.n17_adj_1649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5738_2_lut_3_lut_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34336\,
            in1 => \N__34853\,
            in2 => \_gnd_net_\,
            in3 => \N__34276\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5739_2_lut_3_lut_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__34277\,
            in1 => \N__35846\,
            in2 => \_gnd_net_\,
            in3 => \N__34337\,
            lcout => \c0.n12_adj_1634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5737_2_lut_3_lut_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34335\,
            in1 => \N__34875\,
            in2 => \_gnd_net_\,
            in3 => \N__34275\,
            lcout => \c0.n14_adj_1639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5735_2_lut_3_lut_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34334\,
            in1 => \N__34916\,
            in2 => \_gnd_net_\,
            in3 => \N__34274\,
            lcout => \c0.n16_adj_1641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_668_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34540\,
            in2 => \_gnd_net_\,
            in3 => \N__34154\,
            lcout => \c0.n117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_2_lut_3_lut_4_lut_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__35534\,
            in1 => \N__34419\,
            in2 => \N__34502\,
            in3 => \N__34541\,
            lcout => n3747,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_prev_1994_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx_active_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7727_3_lut_4_lut_4_lut_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001110000000"
        )
    port map (
            in0 => \N__35735\,
            in1 => \N__34420\,
            in2 => \N__34503\,
            in3 => \N__34542\,
            lcout => OPEN,
            ltout => \n8749_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010111010"
        )
    port map (
            in0 => \N__34155\,
            in1 => \N__35535\,
            in2 => \N__34161\,
            in3 => \N__34428\,
            lcout => tx_active,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7389_2_lut_3_lut_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__35710\,
            in1 => \N__34410\,
            in2 => \_gnd_net_\,
            in3 => \N__35513\,
            lcout => \c0.tx.n9059\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_3_lut_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__35512\,
            in1 => \_gnd_net_\,
            in2 => \N__34429\,
            in3 => \N__35709\,
            lcout => OPEN,
            ltout => \c0.tx.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_509_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__35683\,
            in1 => \N__34479\,
            in2 => \N__34128\,
            in3 => \N__34578\,
            lcout => \c0.tx.n9027\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__35516\,
            in1 => \N__35736\,
            in2 => \N__34499\,
            in3 => \N__34426\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34425\,
            in1 => \N__34484\,
            in2 => \N__35744\,
            in3 => \N__35515\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i6328_4_lut_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__34424\,
            in2 => \N__34572\,
            in3 => \N__34548\,
            lcout => OPEN,
            ltout => \n3151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110100"
        )
    port map (
            in0 => \N__35737\,
            in1 => \N__34483\,
            in2 => \N__34515\,
            in3 => \N__35514\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_747_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34421\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34486\,
            lcout => n11_adj_1752,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__34627\,
            in1 => \N__35572\,
            in2 => \N__34659\,
            in3 => \N__34603\,
            lcout => OPEN,
            ltout => \c0.tx.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_adj_508_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__35596\,
            in1 => \N__34825\,
            in2 => \N__34506\,
            in3 => \N__35452\,
            lcout => \c0.tx.n23\,
            ltout => \c0.tx.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7651_2_lut_3_lut_4_lut_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__34485\,
            in1 => \N__35689\,
            in2 => \N__34443\,
            in3 => \N__34422\,
            lcout => n9259,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34604\,
            in1 => \_gnd_net_\,
            in2 => \N__35556\,
            in3 => \N__34590\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_15_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34826\,
            in1 => \N__35550\,
            in2 => \_gnd_net_\,
            in3 => \N__34812\,
            lcout => \r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_510_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34668\,
            lcout => \c0.tx.n7916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34628\,
            in1 => \N__35546\,
            in2 => \_gnd_net_\,
            in3 => \N__34614\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34792\,
            in1 => \N__34751\,
            in2 => \_gnd_net_\,
            in3 => \N__34662\,
            lcout => n9249,
            ltout => OPEN,
            carryin => \bfn_15_30_0_\,
            carryout => \c0.tx.n8090\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34796\,
            in1 => \N__34657\,
            in2 => \_gnd_net_\,
            in3 => \N__34632\,
            lcout => \c0.tx.n9290\,
            ltout => OPEN,
            carryin => \c0.tx.n8090\,
            carryout => \c0.tx.n8091\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34793\,
            in1 => \N__34629\,
            in2 => \_gnd_net_\,
            in3 => \N__34608\,
            lcout => \c0.tx.n9313\,
            ltout => OPEN,
            carryin => \c0.tx.n8091\,
            carryout => \c0.tx.n8092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_15_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34797\,
            in1 => \N__34605\,
            in2 => \_gnd_net_\,
            in3 => \N__34584\,
            lcout => \c0.tx.n9281\,
            ltout => OPEN,
            carryin => \c0.tx.n8092\,
            carryout => \c0.tx.n8093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34794\,
            in1 => \N__35597\,
            in2 => \_gnd_net_\,
            in3 => \N__34581\,
            lcout => n9305,
            ltout => OPEN,
            carryin => \c0.tx.n8093\,
            carryout => \c0.tx.n8094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34798\,
            in1 => \N__35573\,
            in2 => \_gnd_net_\,
            in3 => \N__34830\,
            lcout => \c0.tx.n9314\,
            ltout => OPEN,
            carryin => \c0.tx.n8094\,
            carryout => \c0.tx.n8095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34795\,
            in1 => \N__34827\,
            in2 => \_gnd_net_\,
            in3 => \N__34806\,
            lcout => n9304,
            ltout => OPEN,
            carryin => \c0.tx.n8095\,
            carryout => \c0.tx.n8096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_15_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34799\,
            in1 => \N__35453\,
            in2 => \_gnd_net_\,
            in3 => \N__34803\,
            lcout => n9303,
            ltout => OPEN,
            carryin => \c0.tx.n8096\,
            carryout => \c0.tx.n8097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__34800\,
            in1 => \N__35681\,
            in2 => \_gnd_net_\,
            in3 => \N__34761\,
            lcout => n9266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34758\,
            in1 => \N__34752\,
            in2 => \_gnd_net_\,
            in3 => \N__35551\,
            lcout => \r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_15_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35682\,
            in1 => \N__35552\,
            in2 => \_gnd_net_\,
            in3 => \N__34740\,
            lcout => \r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i0_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34734\,
            in2 => \N__34728\,
            in3 => \_gnd_net_\,
            lcout => \c0.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => \c0.n8120\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i1_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34704\,
            in2 => \_gnd_net_\,
            in3 => \N__34689\,
            lcout => \c0.delay_counter_1\,
            ltout => OPEN,
            carryin => \c0.n8120\,
            carryout => \c0.n8121\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i2_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34686\,
            in2 => \_gnd_net_\,
            in3 => \N__34671\,
            lcout => \c0.delay_counter_2\,
            ltout => OPEN,
            carryin => \c0.n8121\,
            carryout => \c0.n8122\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i3_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34989\,
            in2 => \_gnd_net_\,
            in3 => \N__34968\,
            lcout => \c0.delay_counter_3\,
            ltout => OPEN,
            carryin => \c0.n8122\,
            carryout => \c0.n8123\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i4_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34965\,
            in2 => \_gnd_net_\,
            in3 => \N__34947\,
            lcout => \c0.delay_counter_4\,
            ltout => OPEN,
            carryin => \c0.n8123\,
            carryout => \c0.n8124\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i5_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34944\,
            in2 => \_gnd_net_\,
            in3 => \N__34926\,
            lcout => \c0.delay_counter_5\,
            ltout => OPEN,
            carryin => \c0.n8124\,
            carryout => \c0.n8125\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i6_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34923\,
            in2 => \_gnd_net_\,
            in3 => \N__34902\,
            lcout => \c0.delay_counter_6\,
            ltout => OPEN,
            carryin => \c0.n8125\,
            carryout => \c0.n8126\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i7_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34899\,
            in2 => \_gnd_net_\,
            in3 => \N__34884\,
            lcout => \c0.delay_counter_7\,
            ltout => OPEN,
            carryin => \c0.n8126\,
            carryout => \c0.n8127\,
            clk => \N__35422\,
            ce => \N__35832\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i8_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34881\,
            in2 => \_gnd_net_\,
            in3 => \N__34863\,
            lcout => \c0.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_16_26_0_\,
            carryout => \c0.n8128\,
            clk => \N__35428\,
            ce => \N__35831\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i9_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34860\,
            in2 => \_gnd_net_\,
            in3 => \N__34839\,
            lcout => \c0.delay_counter_9\,
            ltout => OPEN,
            carryin => \c0.n8128\,
            carryout => \c0.n8129\,
            clk => \N__35428\,
            ce => \N__35831\,
            sr => \_gnd_net_\
        );

    \c0.delay_counter_424__i10_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34836\,
            in2 => \_gnd_net_\,
            in3 => \N__35853\,
            lcout => \c0.delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35428\,
            ce => \N__35831\,
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35690\,
            in2 => \_gnd_net_\,
            in3 => \N__35711\,
            lcout => \r_SM_Main_2_N_1480_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i7696_2_lut_3_lut_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__35712\,
            in1 => \_gnd_net_\,
            in2 => \N__35694\,
            in3 => \N__35649\,
            lcout => \c0.tx.n9310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35539\,
            in1 => \N__35598\,
            in2 => \_gnd_net_\,
            in3 => \N__35604\,
            lcout => \r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_16_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35554\,
            in1 => \N__35574\,
            in2 => \_gnd_net_\,
            in3 => \N__35580\,
            lcout => \c0.tx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35555\,
            in1 => \N__35454\,
            in2 => \_gnd_net_\,
            in3 => \N__35460\,
            lcout => \r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35436\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
